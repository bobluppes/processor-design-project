library ieee;
use ieee.std_logic_1164.all;

package main_pack_zynq is

    constant cpu_width : integer := 32;
    constant ram_size : integer := 78971;
    subtype word_type is std_logic_vector(cpu_width-1 downto 0);
    type ram_type is array(0 to ram_size-1) of word_type;
    function load_hex return ram_type;
end package;

package body main_pack_zynq is

    function load_hex return ram_type is
        variable ram_buffer : ram_type := (others=>(others=>'0'));
    begin
        ram_buffer(0) := X"3C1C100D";
        ram_buffer(1) := X"279C5050";
        ram_buffer(2) := X"3C05100D";
        ram_buffer(3) := X"24A5D1EC";
        ram_buffer(4) := X"3C04100D";
        ram_buffer(5) := X"2484DEC4";
        ram_buffer(6) := X"3C1D11FF";
        ram_buffer(7) := X"37BDFF00";
        ram_buffer(8) := X"ACA00000";
        ram_buffer(9) := X"00A4182A";
        ram_buffer(10) := X"1460FFFD";
        ram_buffer(11) := X"24A50004";
        ram_buffer(12) := X"0C02001C";
        ram_buffer(13) := X"00000000";
        ram_buffer(14) := X"27A50020";
        ram_buffer(15) := X"27A60028";
        ram_buffer(16) := X"ACA00000";
        ram_buffer(17) := X"ACC00000";
        ram_buffer(18) := X"0C0200CE";
        ram_buffer(19) := X"00002021";
        ram_buffer(20) := X"08020014";
        ram_buffer(21) := X"00000000";
        ram_buffer(22) := X"00000100";
        ram_buffer(23) := X"01000003";
        ram_buffer(24) := X"00000000";
        ram_buffer(25) := X"00000000";
        ram_buffer(26) := X"00000000";
        ram_buffer(27) := X"00000000";
        ram_buffer(28) := X"27BDFFE0";
        ram_buffer(29) := X"AFBF0014";
        ram_buffer(30) := X"04110001";
        ram_buffer(31) := X"00000000";
        ram_buffer(32) := X"0C02017C";
        ram_buffer(33) := X"00000000";
        ram_buffer(34) := X"04110001";
        ram_buffer(35) := X"00000000";
        ram_buffer(36) := X"0C031D53";
        ram_buffer(37) := X"00000000";
        ram_buffer(38) := X"8FBF0014";
        ram_buffer(39) := X"27BD0020";
        ram_buffer(40) := X"03E00008";
        ram_buffer(41) := X"00000000";
        ram_buffer(42) := X"8F828098";
        ram_buffer(43) := X"8F8681A4";
        ram_buffer(44) := X"8C44000C";
        ram_buffer(45) := X"3C05100C";
        ram_buffer(46) := X"27BDFFE8";
        ram_buffer(47) := X"24A575D8";
        ram_buffer(48) := X"AFBF0014";
        ram_buffer(49) := X"0C027196";
        ram_buffer(50) := X"AFB00010";
        ram_buffer(51) := X"8F828098";
        ram_buffer(52) := X"3C04100C";
        ram_buffer(53) := X"8C47000C";
        ram_buffer(54) := X"2406000C";
        ram_buffer(55) := X"24050001";
        ram_buffer(56) := X"0C0278D7";
        ram_buffer(57) := X"248475F0";
        ram_buffer(58) := X"8F828098";
        ram_buffer(59) := X"3C04100C";
        ram_buffer(60) := X"8C47000C";
        ram_buffer(61) := X"24060025";
        ram_buffer(62) := X"24050001";
        ram_buffer(63) := X"0C0278D7";
        ram_buffer(64) := X"24847600";
        ram_buffer(65) := X"8F828098";
        ram_buffer(66) := X"3C04100C";
        ram_buffer(67) := X"8C47000C";
        ram_buffer(68) := X"24060044";
        ram_buffer(69) := X"24050001";
        ram_buffer(70) := X"0C0278D7";
        ram_buffer(71) := X"24847628";
        ram_buffer(72) := X"8F828098";
        ram_buffer(73) := X"3C04100C";
        ram_buffer(74) := X"8C47000C";
        ram_buffer(75) := X"2406002D";
        ram_buffer(76) := X"24050001";
        ram_buffer(77) := X"0C0278D7";
        ram_buffer(78) := X"24847670";
        ram_buffer(79) := X"8F828098";
        ram_buffer(80) := X"3C04100C";
        ram_buffer(81) := X"8C47000C";
        ram_buffer(82) := X"2406004D";
        ram_buffer(83) := X"24050001";
        ram_buffer(84) := X"0C0278D7";
        ram_buffer(85) := X"248476A0";
        ram_buffer(86) := X"8F828098";
        ram_buffer(87) := X"3C04100C";
        ram_buffer(88) := X"8C47000C";
        ram_buffer(89) := X"2406002E";
        ram_buffer(90) := X"24050001";
        ram_buffer(91) := X"0C0278D7";
        ram_buffer(92) := X"248476F0";
        ram_buffer(93) := X"8F828098";
        ram_buffer(94) := X"3C04100C";
        ram_buffer(95) := X"8C47000C";
        ram_buffer(96) := X"24060041";
        ram_buffer(97) := X"24050001";
        ram_buffer(98) := X"0C0278D7";
        ram_buffer(99) := X"24847720";
        ram_buffer(100) := X"8F828098";
        ram_buffer(101) := X"3C04100C";
        ram_buffer(102) := X"8C47000C";
        ram_buffer(103) := X"2406001D";
        ram_buffer(104) := X"24050001";
        ram_buffer(105) := X"0C0278D7";
        ram_buffer(106) := X"24847764";
        ram_buffer(107) := X"8F828098";
        ram_buffer(108) := X"3C06100C";
        ram_buffer(109) := X"8C44000C";
        ram_buffer(110) := X"3C05100C";
        ram_buffer(111) := X"24C67784";
        ram_buffer(112) := X"0C027196";
        ram_buffer(113) := X"24A57790";
        ram_buffer(114) := X"8F828098";
        ram_buffer(115) := X"3C10100C";
        ram_buffer(116) := X"8C44000C";
        ram_buffer(117) := X"3C05100C";
        ram_buffer(118) := X"2606766C";
        ram_buffer(119) := X"0C027196";
        ram_buffer(120) := X"24A577BC";
        ram_buffer(121) := X"8F828098";
        ram_buffer(122) := X"3C05100C";
        ram_buffer(123) := X"8C44000C";
        ram_buffer(124) := X"2606766C";
        ram_buffer(125) := X"0C027196";
        ram_buffer(126) := X"24A577F8";
        ram_buffer(127) := X"8F828098";
        ram_buffer(128) := X"3C04100C";
        ram_buffer(129) := X"8C47000C";
        ram_buffer(130) := X"24060043";
        ram_buffer(131) := X"24050001";
        ram_buffer(132) := X"0C0278D7";
        ram_buffer(133) := X"2484782C";
        ram_buffer(134) := X"8F828098";
        ram_buffer(135) := X"3C04100C";
        ram_buffer(136) := X"8C47000C";
        ram_buffer(137) := X"2406003E";
        ram_buffer(138) := X"24050001";
        ram_buffer(139) := X"0C0278D7";
        ram_buffer(140) := X"24847870";
        ram_buffer(141) := X"8F828098";
        ram_buffer(142) := X"3C04100C";
        ram_buffer(143) := X"8C47000C";
        ram_buffer(144) := X"24060033";
        ram_buffer(145) := X"24050001";
        ram_buffer(146) := X"0C0278D7";
        ram_buffer(147) := X"248478B0";
        ram_buffer(148) := X"8F828098";
        ram_buffer(149) := X"3C04100C";
        ram_buffer(150) := X"8C47000C";
        ram_buffer(151) := X"2406002E";
        ram_buffer(152) := X"24050001";
        ram_buffer(153) := X"0C0278D7";
        ram_buffer(154) := X"248478E4";
        ram_buffer(155) := X"8F828098";
        ram_buffer(156) := X"3C04100C";
        ram_buffer(157) := X"8C47000C";
        ram_buffer(158) := X"2406002B";
        ram_buffer(159) := X"24050001";
        ram_buffer(160) := X"0C0278D7";
        ram_buffer(161) := X"24847914";
        ram_buffer(162) := X"8F828098";
        ram_buffer(163) := X"3C04100C";
        ram_buffer(164) := X"8C47000C";
        ram_buffer(165) := X"24060016";
        ram_buffer(166) := X"24050001";
        ram_buffer(167) := X"0C0278D7";
        ram_buffer(168) := X"24847940";
        ram_buffer(169) := X"8F828098";
        ram_buffer(170) := X"3C04100C";
        ram_buffer(171) := X"8C47000C";
        ram_buffer(172) := X"24060027";
        ram_buffer(173) := X"24050001";
        ram_buffer(174) := X"0C0278D7";
        ram_buffer(175) := X"24847958";
        ram_buffer(176) := X"8F828098";
        ram_buffer(177) := X"3C04100C";
        ram_buffer(178) := X"8C47000C";
        ram_buffer(179) := X"24060037";
        ram_buffer(180) := X"24050001";
        ram_buffer(181) := X"0C0278D7";
        ram_buffer(182) := X"24847980";
        ram_buffer(183) := X"8F828098";
        ram_buffer(184) := X"3C04100C";
        ram_buffer(185) := X"8C47000C";
        ram_buffer(186) := X"24060037";
        ram_buffer(187) := X"24050001";
        ram_buffer(188) := X"0C0278D7";
        ram_buffer(189) := X"248479B8";
        ram_buffer(190) := X"8F828098";
        ram_buffer(191) := X"3C04100C";
        ram_buffer(192) := X"8C47000C";
        ram_buffer(193) := X"24060034";
        ram_buffer(194) := X"24050001";
        ram_buffer(195) := X"0C0278D7";
        ram_buffer(196) := X"248479F0";
        ram_buffer(197) := X"8F828098";
        ram_buffer(198) := X"3C04100C";
        ram_buffer(199) := X"8C47000C";
        ram_buffer(200) := X"24847A28";
        ram_buffer(201) := X"24060038";
        ram_buffer(202) := X"0C0278D7";
        ram_buffer(203) := X"24050001";
        ram_buffer(204) := X"0C026D37";
        ram_buffer(205) := X"24040001";
        ram_buffer(206) := X"27BDFD98";
        ram_buffer(207) := X"3C05100C";
        ram_buffer(208) := X"AFB3025C";
        ram_buffer(209) := X"27B3023C";
        ram_buffer(210) := X"02602021";
        ram_buffer(211) := X"2406000D";
        ram_buffer(212) := X"24A57CBC";
        ram_buffer(213) := X"AFBF0264";
        ram_buffer(214) := X"AFB40260";
        ram_buffer(215) := X"AFB20258";
        ram_buffer(216) := X"AFB10254";
        ram_buffer(217) := X"0C027F93";
        ram_buffer(218) := X"AFB00250";
        ram_buffer(219) := X"3C05100C";
        ram_buffer(220) := X"24060013";
        ram_buffer(221) := X"24A57CCC";
        ram_buffer(222) := X"0C027F93";
        ram_buffer(223) := X"27A40228";
        ram_buffer(224) := X"3C02100C";
        ram_buffer(225) := X"24427BCC";
        ram_buffer(226) := X"AFA20210";
        ram_buffer(227) := X"3C02100C";
        ram_buffer(228) := X"24427C0C";
        ram_buffer(229) := X"AFA20214";
        ram_buffer(230) := X"3C02100C";
        ram_buffer(231) := X"24427C18";
        ram_buffer(232) := X"AFA20218";
        ram_buffer(233) := X"3C02100C";
        ram_buffer(234) := X"24427C1C";
        ram_buffer(235) := X"AFA2021C";
        ram_buffer(236) := X"3C02100C";
        ram_buffer(237) := X"2442766C";
        ram_buffer(238) := X"AFA20220";
        ram_buffer(239) := X"3C04100C";
        ram_buffer(240) := X"3C02100C";
        ram_buffer(241) := X"24847C38";
        ram_buffer(242) := X"24427C28";
        ram_buffer(243) := X"0C028186";
        ram_buffer(244) := X"AFA20224";
        ram_buffer(245) := X"0C03070B";
        ram_buffer(246) := X"AFB30220";
        ram_buffer(247) := X"27A50210";
        ram_buffer(248) := X"24040006";
        ram_buffer(249) := X"00608821";
        ram_buffer(250) := X"0C020366";
        ram_buffer(251) := X"0040A021";
        ram_buffer(252) := X"0C03070B";
        ram_buffer(253) := X"00000000";
        ram_buffer(254) := X"27A60010";
        ram_buffer(255) := X"02602821";
        ram_buffer(256) := X"27A40228";
        ram_buffer(257) := X"00608021";
        ram_buffer(258) := X"00409021";
        ram_buffer(259) := X"0C0303D0";
        ram_buffer(260) := X"3C13100C";
        ram_buffer(261) := X"0C028186";
        ram_buffer(262) := X"27A40010";
        ram_buffer(263) := X"0C028186";
        ram_buffer(264) := X"26647C54";
        ram_buffer(265) := X"02112823";
        ram_buffer(266) := X"0205802B";
        ram_buffer(267) := X"02542023";
        ram_buffer(268) := X"0C031C00";
        ram_buffer(269) := X"00902023";
        ram_buffer(270) := X"8F87801C";
        ram_buffer(271) := X"8F868018";
        ram_buffer(272) := X"00602821";
        ram_buffer(273) := X"0C03144F";
        ram_buffer(274) := X"00402021";
        ram_buffer(275) := X"3C04100C";
        ram_buffer(276) := X"00603821";
        ram_buffer(277) := X"00403021";
        ram_buffer(278) := X"0C028116";
        ram_buffer(279) := X"24847C90";
        ram_buffer(280) := X"0C028186";
        ram_buffer(281) := X"26647C54";
        ram_buffer(282) := X"3C04100C";
        ram_buffer(283) := X"240500FE";
        ram_buffer(284) := X"0C028116";
        ram_buffer(285) := X"24847CB8";
        ram_buffer(286) := X"8FBF0264";
        ram_buffer(287) := X"8FB40260";
        ram_buffer(288) := X"8FB3025C";
        ram_buffer(289) := X"8FB20258";
        ram_buffer(290) := X"8FB10254";
        ram_buffer(291) := X"8FB00250";
        ram_buffer(292) := X"00001021";
        ram_buffer(293) := X"03E00008";
        ram_buffer(294) := X"27BD0268";
        ram_buffer(295) := X"3C04100D";
        ram_buffer(296) := X"3C02100D";
        ram_buffer(297) := X"2484D060";
        ram_buffer(298) := X"2442D063";
        ram_buffer(299) := X"00441023";
        ram_buffer(300) := X"2C420007";
        ram_buffer(301) := X"14400006";
        ram_buffer(302) := X"3C190000";
        ram_buffer(303) := X"27390000";
        ram_buffer(304) := X"13200003";
        ram_buffer(305) := X"00000000";
        ram_buffer(306) := X"03200008";
        ram_buffer(307) := X"00000000";
        ram_buffer(308) := X"03E00008";
        ram_buffer(309) := X"00000000";
        ram_buffer(310) := X"3C04100D";
        ram_buffer(311) := X"3C02100D";
        ram_buffer(312) := X"2484D060";
        ram_buffer(313) := X"2442D060";
        ram_buffer(314) := X"00441023";
        ram_buffer(315) := X"00021083";
        ram_buffer(316) := X"00022FC2";
        ram_buffer(317) := X"00A22821";
        ram_buffer(318) := X"00052843";
        ram_buffer(319) := X"10A00006";
        ram_buffer(320) := X"3C190000";
        ram_buffer(321) := X"27390000";
        ram_buffer(322) := X"13200003";
        ram_buffer(323) := X"00000000";
        ram_buffer(324) := X"03200008";
        ram_buffer(325) := X"00000000";
        ram_buffer(326) := X"03E00008";
        ram_buffer(327) := X"00000000";
        ram_buffer(328) := X"27BDFFD8";
        ram_buffer(329) := X"AFB30020";
        ram_buffer(330) := X"3C13100D";
        ram_buffer(331) := X"9262D240";
        ram_buffer(332) := X"AFBF0024";
        ram_buffer(333) := X"AFB2001C";
        ram_buffer(334) := X"AFB10018";
        ram_buffer(335) := X"14400025";
        ram_buffer(336) := X"AFB00014";
        ram_buffer(337) := X"3C11100D";
        ram_buffer(338) := X"3C02100D";
        ram_buffer(339) := X"2442C7AC";
        ram_buffer(340) := X"2631C7A8";
        ram_buffer(341) := X"00518823";
        ram_buffer(342) := X"3C10100D";
        ram_buffer(343) := X"8E02D244";
        ram_buffer(344) := X"00118883";
        ram_buffer(345) := X"2631FFFF";
        ram_buffer(346) := X"3C04100D";
        ram_buffer(347) := X"0051182B";
        ram_buffer(348) := X"2492C7A8";
        ram_buffer(349) := X"1060000C";
        ram_buffer(350) := X"24420001";
        ram_buffer(351) := X"00021880";
        ram_buffer(352) := X"02431821";
        ram_buffer(353) := X"8C630000";
        ram_buffer(354) := X"00000000";
        ram_buffer(355) := X"0060F809";
        ram_buffer(356) := X"AE02D244";
        ram_buffer(357) := X"8E02D244";
        ram_buffer(358) := X"00000000";
        ram_buffer(359) := X"0051182B";
        ram_buffer(360) := X"1460FFF6";
        ram_buffer(361) := X"24420001";
        ram_buffer(362) := X"0C020127";
        ram_buffer(363) := X"00000000";
        ram_buffer(364) := X"3C020000";
        ram_buffer(365) := X"24420000";
        ram_buffer(366) := X"10400005";
        ram_buffer(367) := X"24020001";
        ram_buffer(368) := X"3C04100D";
        ram_buffer(369) := X"0C000000";
        ram_buffer(370) := X"2484B760";
        ram_buffer(371) := X"24020001";
        ram_buffer(372) := X"A262D240";
        ram_buffer(373) := X"8FBF0024";
        ram_buffer(374) := X"8FB30020";
        ram_buffer(375) := X"8FB2001C";
        ram_buffer(376) := X"8FB10018";
        ram_buffer(377) := X"8FB00014";
        ram_buffer(378) := X"03E00008";
        ram_buffer(379) := X"27BD0028";
        ram_buffer(380) := X"3C020000";
        ram_buffer(381) := X"27BDFFE8";
        ram_buffer(382) := X"24420000";
        ram_buffer(383) := X"10400006";
        ram_buffer(384) := X"AFBF0014";
        ram_buffer(385) := X"3C05100D";
        ram_buffer(386) := X"3C04100D";
        ram_buffer(387) := X"24A5D248";
        ram_buffer(388) := X"0C000000";
        ram_buffer(389) := X"2484B760";
        ram_buffer(390) := X"3C02100D";
        ram_buffer(391) := X"2444C7B0";
        ram_buffer(392) := X"8C820000";
        ram_buffer(393) := X"00000000";
        ram_buffer(394) := X"14400004";
        ram_buffer(395) := X"3C020000";
        ram_buffer(396) := X"8FBF0014";
        ram_buffer(397) := X"08020136";
        ram_buffer(398) := X"27BD0018";
        ram_buffer(399) := X"24420000";
        ram_buffer(400) := X"1040FFFB";
        ram_buffer(401) := X"00000000";
        ram_buffer(402) := X"0040F809";
        ram_buffer(403) := X"00000000";
        ram_buffer(404) := X"1000FFF7";
        ram_buffer(405) := X"00000000";
        ram_buffer(406) := X"27BDFF80";
        ram_buffer(407) := X"8C830000";
        ram_buffer(408) := X"28A20002";
        ram_buffer(409) := X"AFB5006C";
        ram_buffer(410) := X"00A0A821";
        ram_buffer(411) := X"2405004B";
        ram_buffer(412) := X"AFB70074";
        ram_buffer(413) := X"AFBF007C";
        ram_buffer(414) := X"AFBE0078";
        ram_buffer(415) := X"AFB60070";
        ram_buffer(416) := X"AFB40068";
        ram_buffer(417) := X"AFB30064";
        ram_buffer(418) := X"AFB20060";
        ram_buffer(419) := X"AFB1005C";
        ram_buffer(420) := X"AFB00058";
        ram_buffer(421) := X"00E0B821";
        ram_buffer(422) := X"AFA5001C";
        ram_buffer(423) := X"AF8081A8";
        ram_buffer(424) := X"AF8081A0";
        ram_buffer(425) := X"144000A1";
        ram_buffer(426) := X"AC600068";
        ram_buffer(427) := X"24020064";
        ram_buffer(428) := X"3C11100C";
        ram_buffer(429) := X"AFA20040";
        ram_buffer(430) := X"26227A64";
        ram_buffer(431) := X"AFA20038";
        ram_buffer(432) := X"3C02100C";
        ram_buffer(433) := X"24427A9C";
        ram_buffer(434) := X"AFA2003C";
        ram_buffer(435) := X"3C02100C";
        ram_buffer(436) := X"AFA20044";
        ram_buffer(437) := X"3C02100C";
        ram_buffer(438) := X"24427AC0";
        ram_buffer(439) := X"AFA20048";
        ram_buffer(440) := X"3C02100C";
        ram_buffer(441) := X"0080A021";
        ram_buffer(442) := X"00C0B021";
        ram_buffer(443) := X"00009821";
        ram_buffer(444) := X"AFA00028";
        ram_buffer(445) := X"AFA0002C";
        ram_buffer(446) := X"AFA00030";
        ram_buffer(447) := X"AFA00034";
        ram_buffer(448) := X"00009021";
        ram_buffer(449) := X"241E0001";
        ram_buffer(450) := X"AFA2004C";
        ram_buffer(451) := X"001E3880";
        ram_buffer(452) := X"02C78821";
        ram_buffer(453) := X"8E300000";
        ram_buffer(454) := X"2402002D";
        ram_buffer(455) := X"82040000";
        ram_buffer(456) := X"00000000";
        ram_buffer(457) := X"10820010";
        ram_buffer(458) := X"24060001";
        ram_buffer(459) := X"16E00023";
        ram_buffer(460) := X"00000000";
        ram_buffer(461) := X"8FBF007C";
        ram_buffer(462) := X"03C01021";
        ram_buffer(463) := X"8FB70074";
        ram_buffer(464) := X"8FBE0078";
        ram_buffer(465) := X"8FB60070";
        ram_buffer(466) := X"8FB5006C";
        ram_buffer(467) := X"8FB40068";
        ram_buffer(468) := X"8FB30064";
        ram_buffer(469) := X"8FB20060";
        ram_buffer(470) := X"8FB1005C";
        ram_buffer(471) := X"8FB00058";
        ram_buffer(472) := X"03E00008";
        ram_buffer(473) := X"27BD0080";
        ram_buffer(474) := X"26100001";
        ram_buffer(475) := X"8FA50038";
        ram_buffer(476) := X"02002021";
        ram_buffer(477) := X"0C021920";
        ram_buffer(478) := X"AFA70050";
        ram_buffer(479) := X"8FA70050";
        ram_buffer(480) := X"144000C0";
        ram_buffer(481) := X"24060001";
        ram_buffer(482) := X"8FA5003C";
        ram_buffer(483) := X"02002021";
        ram_buffer(484) := X"0C021920";
        ram_buffer(485) := X"AFA70050";
        ram_buffer(486) := X"10400036";
        ram_buffer(487) := X"24060002";
        ram_buffer(488) := X"24120001";
        ram_buffer(489) := X"27DE0001";
        ram_buffer(490) := X"03D5102A";
        ram_buffer(491) := X"1440FFD8";
        ram_buffer(492) := X"001E3880";
        ram_buffer(493) := X"12E0FFDF";
        ram_buffer(494) := X"00000000";
        ram_buffer(495) := X"8FA5001C";
        ram_buffer(496) := X"02403021";
        ram_buffer(497) := X"0C021CBA";
        ram_buffer(498) := X"02802021";
        ram_buffer(499) := X"8FA20034";
        ram_buffer(500) := X"00000000";
        ram_buffer(501) := X"10400007";
        ram_buffer(502) := X"02403821";
        ram_buffer(503) := X"8FA60040";
        ram_buffer(504) := X"00402821";
        ram_buffer(505) := X"0C02170E";
        ram_buffer(506) := X"02802021";
        ram_buffer(507) := X"1040001B";
        ram_buffer(508) := X"00000000";
        ram_buffer(509) := X"8FA20030";
        ram_buffer(510) := X"00000000";
        ram_buffer(511) := X"10400005";
        ram_buffer(512) := X"00402821";
        ram_buffer(513) := X"0C021860";
        ram_buffer(514) := X"02802021";
        ram_buffer(515) := X"10400013";
        ram_buffer(516) := X"00000000";
        ram_buffer(517) := X"8FA2002C";
        ram_buffer(518) := X"00000000";
        ram_buffer(519) := X"10400005";
        ram_buffer(520) := X"00402821";
        ram_buffer(521) := X"0C0218B3";
        ram_buffer(522) := X"02802021";
        ram_buffer(523) := X"1040000B";
        ram_buffer(524) := X"00000000";
        ram_buffer(525) := X"8FA20028";
        ram_buffer(526) := X"00000000";
        ram_buffer(527) := X"14400009";
        ram_buffer(528) := X"00000000";
        ram_buffer(529) := X"1260FFBB";
        ram_buffer(530) := X"02602821";
        ram_buffer(531) := X"0C02177C";
        ram_buffer(532) := X"02802021";
        ram_buffer(533) := X"1440FFB7";
        ram_buffer(534) := X"00000000";
        ram_buffer(535) := X"0C02002A";
        ram_buffer(536) := X"00000000";
        ram_buffer(537) := X"0C0220DD";
        ram_buffer(538) := X"02802021";
        ram_buffer(539) := X"1000FFF5";
        ram_buffer(540) := X"00000000";
        ram_buffer(541) := X"8FA20044";
        ram_buffer(542) := X"00000000";
        ram_buffer(543) := X"24457AA8";
        ram_buffer(544) := X"0C021920";
        ram_buffer(545) := X"02002021";
        ram_buffer(546) := X"10400018";
        ram_buffer(547) := X"24060001";
        ram_buffer(548) := X"27DE0001";
        ram_buffer(549) := X"03D5102A";
        ram_buffer(550) := X"8FA70050";
        ram_buffer(551) := X"1040FFEF";
        ram_buffer(552) := X"3C05100C";
        ram_buffer(553) := X"24F00004";
        ram_buffer(554) := X"02D08021";
        ram_buffer(555) := X"8E040000";
        ram_buffer(556) := X"24060001";
        ram_buffer(557) := X"0C021920";
        ram_buffer(558) := X"24A57AAC";
        ram_buffer(559) := X"10400003";
        ram_buffer(560) := X"24060002";
        ram_buffer(561) := X"1000FFB7";
        ram_buffer(562) := X"AE8000BC";
        ram_buffer(563) := X"3C05100C";
        ram_buffer(564) := X"8E040000";
        ram_buffer(565) := X"0C021920";
        ram_buffer(566) := X"24A57AB0";
        ram_buffer(567) := X"1040003F";
        ram_buffer(568) := X"24020001";
        ram_buffer(569) := X"1000FFAF";
        ram_buffer(570) := X"AE8200BC";
        ram_buffer(571) := X"8FA50048";
        ram_buffer(572) := X"0C021920";
        ram_buffer(573) := X"02002021";
        ram_buffer(574) := X"10400014";
        ram_buffer(575) := X"24060001";
        ram_buffer(576) := X"8F82819C";
        ram_buffer(577) := X"00000000";
        ram_buffer(578) := X"10400028";
        ram_buffer(579) := X"3C07100C";
        ram_buffer(580) := X"8E840000";
        ram_buffer(581) := X"00000000";
        ram_buffer(582) := X"8C820068";
        ram_buffer(583) := X"00000000";
        ram_buffer(584) := X"24420001";
        ram_buffer(585) := X"1000FF9F";
        ram_buffer(586) := X"AC820068";
        ram_buffer(587) := X"14E00003";
        ram_buffer(588) := X"00003021";
        ram_buffer(589) := X"1000FF7F";
        ram_buffer(590) := X"241E0001";
        ram_buffer(591) := X"0C021CBA";
        ram_buffer(592) := X"2405004B";
        ram_buffer(593) := X"1000FF7B";
        ram_buffer(594) := X"241E0001";
        ram_buffer(595) := X"8FA2004C";
        ram_buffer(596) := X"00000000";
        ram_buffer(597) := X"24457AC8";
        ram_buffer(598) := X"0C021920";
        ram_buffer(599) := X"02002021";
        ram_buffer(600) := X"1440FFE7";
        ram_buffer(601) := X"3C05100C";
        ram_buffer(602) := X"24060002";
        ram_buffer(603) := X"24A57B34";
        ram_buffer(604) := X"0C021920";
        ram_buffer(605) := X"02002021";
        ram_buffer(606) := X"14400008";
        ram_buffer(607) := X"24050001";
        ram_buffer(608) := X"3C05100C";
        ram_buffer(609) := X"24060002";
        ram_buffer(610) := X"24A57B40";
        ram_buffer(611) := X"0C021920";
        ram_buffer(612) := X"02002021";
        ram_buffer(613) := X"1040001A";
        ram_buffer(614) := X"24050001";
        ram_buffer(615) := X"0C021E7D";
        ram_buffer(616) := X"02802021";
        ram_buffer(617) := X"1000FF80";
        ram_buffer(618) := X"27DE0001";
        ram_buffer(619) := X"8F828098";
        ram_buffer(620) := X"00000000";
        ram_buffer(621) := X"8C44000C";
        ram_buffer(622) := X"3C06100C";
        ram_buffer(623) := X"3C05100C";
        ram_buffer(624) := X"24E77AD0";
        ram_buffer(625) := X"24C67AF4";
        ram_buffer(626) := X"0C027196";
        ram_buffer(627) := X"24A57B04";
        ram_buffer(628) := X"24020001";
        ram_buffer(629) := X"1000FFCE";
        ram_buffer(630) := X"AF82819C";
        ram_buffer(631) := X"3C05100C";
        ram_buffer(632) := X"8E040000";
        ram_buffer(633) := X"24060002";
        ram_buffer(634) := X"0C021920";
        ram_buffer(635) := X"24A57AB8";
        ram_buffer(636) := X"1040FF9A";
        ram_buffer(637) := X"24020002";
        ram_buffer(638) := X"1000FF6A";
        ram_buffer(639) := X"AE8200BC";
        ram_buffer(640) := X"3C05100C";
        ram_buffer(641) := X"24060003";
        ram_buffer(642) := X"24A57B4C";
        ram_buffer(643) := X"0C021920";
        ram_buffer(644) := X"02002021";
        ram_buffer(645) := X"10400029";
        ram_buffer(646) := X"24040078";
        ram_buffer(647) := X"27DE0001";
        ram_buffer(648) := X"03D5102A";
        ram_buffer(649) := X"1040FF8D";
        ram_buffer(650) := X"A3A40021";
        ram_buffer(651) := X"3C05100C";
        ram_buffer(652) := X"8E240004";
        ram_buffer(653) := X"27A70021";
        ram_buffer(654) := X"27A60018";
        ram_buffer(655) := X"0C028409";
        ram_buffer(656) := X"24A57B58";
        ram_buffer(657) := X"1840FF85";
        ram_buffer(658) := X"00000000";
        ram_buffer(659) := X"93A20021";
        ram_buffer(660) := X"2404004D";
        ram_buffer(661) := X"304200DF";
        ram_buffer(662) := X"00021600";
        ram_buffer(663) := X"00021603";
        ram_buffer(664) := X"10440010";
        ram_buffer(665) := X"240403E8";
        ram_buffer(666) := X"8FA20018";
        ram_buffer(667) := X"240403E8";
        ram_buffer(668) := X"00440018";
        ram_buffer(669) := X"8E840004";
        ram_buffer(670) := X"00001012";
        ram_buffer(671) := X"1000FF49";
        ram_buffer(672) := X"AC82002C";
        ram_buffer(673) := X"8F828098";
        ram_buffer(674) := X"8F8681A4";
        ram_buffer(675) := X"8C44000C";
        ram_buffer(676) := X"3C05100C";
        ram_buffer(677) := X"0C027196";
        ram_buffer(678) := X"24A57A70";
        ram_buffer(679) := X"0C026D37";
        ram_buffer(680) := X"24040001";
        ram_buffer(681) := X"8FA20018";
        ram_buffer(682) := X"00000000";
        ram_buffer(683) := X"00440018";
        ram_buffer(684) := X"00001012";
        ram_buffer(685) := X"1000FFED";
        ram_buffer(686) := X"AFA20018";
        ram_buffer(687) := X"3C05100C";
        ram_buffer(688) := X"24060001";
        ram_buffer(689) := X"24A57B60";
        ram_buffer(690) := X"0C021920";
        ram_buffer(691) := X"02002021";
        ram_buffer(692) := X"10400004";
        ram_buffer(693) := X"3C05100C";
        ram_buffer(694) := X"24020001";
        ram_buffer(695) := X"1000FF31";
        ram_buffer(696) := X"AE8200B0";
        ram_buffer(697) := X"24060001";
        ram_buffer(698) := X"24A57B6C";
        ram_buffer(699) := X"0C021920";
        ram_buffer(700) := X"02002021";
        ram_buffer(701) := X"1440FFF9";
        ram_buffer(702) := X"24020001";
        ram_buffer(703) := X"3C05100C";
        ram_buffer(704) := X"24060004";
        ram_buffer(705) := X"24A57B78";
        ram_buffer(706) := X"0C021920";
        ram_buffer(707) := X"02002021";
        ram_buffer(708) := X"10400008";
        ram_buffer(709) := X"3C05100C";
        ram_buffer(710) := X"27DE0001";
        ram_buffer(711) := X"03D5102A";
        ram_buffer(712) := X"1040FF4E";
        ram_buffer(713) := X"00000000";
        ram_buffer(714) := X"8E220004";
        ram_buffer(715) := X"1000FF1D";
        ram_buffer(716) := X"AF8281A0";
        ram_buffer(717) := X"24060001";
        ram_buffer(718) := X"24A57B80";
        ram_buffer(719) := X"0C021920";
        ram_buffer(720) := X"02002021";
        ram_buffer(721) := X"10400003";
        ram_buffer(722) := X"24020001";
        ram_buffer(723) := X"1000FF15";
        ram_buffer(724) := X"AFA20028";
        ram_buffer(725) := X"3C05100C";
        ram_buffer(726) := X"24060001";
        ram_buffer(727) := X"24A57B8C";
        ram_buffer(728) := X"0C021920";
        ram_buffer(729) := X"02002021";
        ram_buffer(730) := X"10400011";
        ram_buffer(731) := X"3C05100C";
        ram_buffer(732) := X"27DE0001";
        ram_buffer(733) := X"03D5102A";
        ram_buffer(734) := X"1040FF38";
        ram_buffer(735) := X"3C05100D";
        ram_buffer(736) := X"8E240004";
        ram_buffer(737) := X"27A6001C";
        ram_buffer(738) := X"0C028409";
        ram_buffer(739) := X"24A59658";
        ram_buffer(740) := X"24040001";
        ram_buffer(741) := X"1444FF31";
        ram_buffer(742) := X"00000000";
        ram_buffer(743) := X"8FA4001C";
        ram_buffer(744) := X"0C021CA3";
        ram_buffer(745) := X"27DE0001";
        ram_buffer(746) := X"1000FEFF";
        ram_buffer(747) := X"AFA20040";
        ram_buffer(748) := X"24060002";
        ram_buffer(749) := X"24A57B94";
        ram_buffer(750) := X"0C021920";
        ram_buffer(751) := X"02002021";
        ram_buffer(752) := X"10400008";
        ram_buffer(753) := X"3C05100C";
        ram_buffer(754) := X"27DE0001";
        ram_buffer(755) := X"03D5102A";
        ram_buffer(756) := X"1040FF22";
        ram_buffer(757) := X"00000000";
        ram_buffer(758) := X"8E220004";
        ram_buffer(759) := X"1000FEF1";
        ram_buffer(760) := X"AFA20030";
        ram_buffer(761) := X"24060002";
        ram_buffer(762) := X"24A57B9C";
        ram_buffer(763) := X"0C021920";
        ram_buffer(764) := X"02002021";
        ram_buffer(765) := X"10400008";
        ram_buffer(766) := X"3C05100C";
        ram_buffer(767) := X"27DE0001";
        ram_buffer(768) := X"03D5102A";
        ram_buffer(769) := X"1040FF15";
        ram_buffer(770) := X"00000000";
        ram_buffer(771) := X"8E220004";
        ram_buffer(772) := X"1000FEE4";
        ram_buffer(773) := X"AFA20034";
        ram_buffer(774) := X"24060001";
        ram_buffer(775) := X"24A57BA4";
        ram_buffer(776) := X"02002021";
        ram_buffer(777) := X"0C021920";
        ram_buffer(778) := X"AFA20050";
        ram_buffer(779) := X"1040001D";
        ram_buffer(780) := X"24040078";
        ram_buffer(781) := X"27DE0001";
        ram_buffer(782) := X"03D5102A";
        ram_buffer(783) := X"1040FF07";
        ram_buffer(784) := X"A3A40020";
        ram_buffer(785) := X"3C05100C";
        ram_buffer(786) := X"8E240004";
        ram_buffer(787) := X"27A70020";
        ram_buffer(788) := X"27A60014";
        ram_buffer(789) := X"0C028409";
        ram_buffer(790) := X"24A57B58";
        ram_buffer(791) := X"1840FEFF";
        ram_buffer(792) := X"3C020001";
        ram_buffer(793) := X"8FA40014";
        ram_buffer(794) := X"00000000";
        ram_buffer(795) := X"0082102B";
        ram_buffer(796) := X"1040FEFA";
        ram_buffer(797) := X"24050042";
        ram_buffer(798) := X"93A20020";
        ram_buffer(799) := X"00000000";
        ram_buffer(800) := X"304200DF";
        ram_buffer(801) := X"00021600";
        ram_buffer(802) := X"00021603";
        ram_buffer(803) := X"8FAD0050";
        ram_buffer(804) := X"10450012";
        ram_buffer(805) := X"00000000";
        ram_buffer(806) := X"00806821";
        ram_buffer(807) := X"1000FEC1";
        ram_buffer(808) := X"AE8D00C4";
        ram_buffer(809) := X"3C05100C";
        ram_buffer(810) := X"24060002";
        ram_buffer(811) := X"24A57BAC";
        ram_buffer(812) := X"0C021920";
        ram_buffer(813) := X"02002021";
        ram_buffer(814) := X"1040000A";
        ram_buffer(815) := X"3C05100C";
        ram_buffer(816) := X"27DE0001";
        ram_buffer(817) := X"03D5102A";
        ram_buffer(818) := X"1040FEE4";
        ram_buffer(819) := X"00000000";
        ram_buffer(820) := X"8E220004";
        ram_buffer(821) := X"1000FEB3";
        ram_buffer(822) := X"AFA2002C";
        ram_buffer(823) := X"1000FFEF";
        ram_buffer(824) := X"AE8400C0";
        ram_buffer(825) := X"24060002";
        ram_buffer(826) := X"24A57BB4";
        ram_buffer(827) := X"0C021920";
        ram_buffer(828) := X"02002021";
        ram_buffer(829) := X"10400008";
        ram_buffer(830) := X"3C05100C";
        ram_buffer(831) := X"27DE0001";
        ram_buffer(832) := X"03D5102A";
        ram_buffer(833) := X"1040FED5";
        ram_buffer(834) := X"00000000";
        ram_buffer(835) := X"8E330004";
        ram_buffer(836) := X"1000FEA5";
        ram_buffer(837) := X"27DE0001";
        ram_buffer(838) := X"24060002";
        ram_buffer(839) := X"24A57BBC";
        ram_buffer(840) := X"0C021920";
        ram_buffer(841) := X"02002021";
        ram_buffer(842) := X"10400013";
        ram_buffer(843) := X"3C05100C";
        ram_buffer(844) := X"27DE0001";
        ram_buffer(845) := X"03D5102A";
        ram_buffer(846) := X"1040FEC8";
        ram_buffer(847) := X"3C05100D";
        ram_buffer(848) := X"8E240004";
        ram_buffer(849) := X"27A60010";
        ram_buffer(850) := X"0C028409";
        ram_buffer(851) := X"24A59658";
        ram_buffer(852) := X"24040001";
        ram_buffer(853) := X"1444FEC1";
        ram_buffer(854) := X"00000000";
        ram_buffer(855) := X"8FA20010";
        ram_buffer(856) := X"00000000";
        ram_buffer(857) := X"2C440065";
        ram_buffer(858) := X"1080FEBC";
        ram_buffer(859) := X"00000000";
        ram_buffer(860) := X"1000FE8C";
        ram_buffer(861) := X"AE8200B8";
        ram_buffer(862) := X"24060001";
        ram_buffer(863) := X"24A57BC4";
        ram_buffer(864) := X"0C021920";
        ram_buffer(865) := X"02002021";
        ram_buffer(866) := X"1040FEB4";
        ram_buffer(867) := X"24020001";
        ram_buffer(868) := X"1000FE84";
        ram_buffer(869) := X"AF8281A8";
        ram_buffer(870) := X"8CA20000";
        ram_buffer(871) := X"27BDFDE8";
        ram_buffer(872) := X"AF8281A4";
        ram_buffer(873) := X"AFB40210";
        ram_buffer(874) := X"AFB20208";
        ram_buffer(875) := X"AFBF0214";
        ram_buffer(876) := X"AFB3020C";
        ram_buffer(877) := X"AFB10204";
        ram_buffer(878) := X"AFB00200";
        ram_buffer(879) := X"00A0A021";
        ram_buffer(880) := X"10400053";
        ram_buffer(881) := X"00809021";
        ram_buffer(882) := X"80420000";
        ram_buffer(883) := X"00000000";
        ram_buffer(884) := X"10400050";
        ram_buffer(885) := X"3C02100C";
        ram_buffer(886) := X"0C02657F";
        ram_buffer(887) := X"27A40178";
        ram_buffer(888) := X"24060168";
        ram_buffer(889) := X"2405003D";
        ram_buffer(890) := X"27A40010";
        ram_buffer(891) := X"0C02194D";
        ram_buffer(892) := X"AFA20010";
        ram_buffer(893) := X"3C02100D";
        ram_buffer(894) := X"24428238";
        ram_buffer(895) := X"AFA201F0";
        ram_buffer(896) := X"240203E8";
        ram_buffer(897) := X"AFA201F4";
        ram_buffer(898) := X"24020413";
        ram_buffer(899) := X"27A40010";
        ram_buffer(900) := X"AFA201F8";
        ram_buffer(901) := X"24020002";
        ram_buffer(902) := X"0C021F65";
        ram_buffer(903) := X"AFA20034";
        ram_buffer(904) := X"00003821";
        ram_buffer(905) := X"02803021";
        ram_buffer(906) := X"02402821";
        ram_buffer(907) := X"0C020196";
        ram_buffer(908) := X"27A40010";
        ram_buffer(909) := X"2643FFFF";
        ram_buffer(910) := X"0043182A";
        ram_buffer(911) := X"146000C9";
        ram_buffer(912) := X"0052182A";
        ram_buffer(913) := X"10600036";
        ram_buffer(914) := X"00021080";
        ram_buffer(915) := X"02828021";
        ram_buffer(916) := X"8E040000";
        ram_buffer(917) := X"3C05100C";
        ram_buffer(918) := X"0C02716A";
        ram_buffer(919) := X"24A57BF0";
        ram_buffer(920) := X"104000B2";
        ram_buffer(921) := X"00408821";
        ram_buffer(922) := X"8F8481A0";
        ram_buffer(923) := X"00000000";
        ram_buffer(924) := X"10800031";
        ram_buffer(925) := X"00000000";
        ram_buffer(926) := X"3C05100C";
        ram_buffer(927) := X"0C02716A";
        ram_buffer(928) := X"24A57C08";
        ram_buffer(929) := X"104000B2";
        ram_buffer(930) := X"00409821";
        ram_buffer(931) := X"8F8281A8";
        ram_buffer(932) := X"00000000";
        ram_buffer(933) := X"1440002F";
        ram_buffer(934) := X"00000000";
        ram_buffer(935) := X"8E220004";
        ram_buffer(936) := X"00000000";
        ram_buffer(937) := X"2442FFFF";
        ram_buffer(938) := X"04400086";
        ram_buffer(939) := X"AE220004";
        ram_buffer(940) := X"8E220000";
        ram_buffer(941) := X"00000000";
        ram_buffer(942) := X"24430001";
        ram_buffer(943) := X"AE230000";
        ram_buffer(944) := X"90500000";
        ram_buffer(945) := X"02202821";
        ram_buffer(946) := X"0C029D83";
        ram_buffer(947) := X"02002021";
        ram_buffer(948) := X"2403FFFF";
        ram_buffer(949) := X"1043008D";
        ram_buffer(950) := X"00000000";
        ram_buffer(951) := X"24020042";
        ram_buffer(952) := X"12020074";
        ram_buffer(953) := X"2A020043";
        ram_buffer(954) := X"14400064";
        ram_buffer(955) := X"24020047";
        ram_buffer(956) := X"1202006C";
        ram_buffer(957) := X"24020050";
        ram_buffer(958) := X"16020062";
        ram_buffer(959) := X"00000000";
        ram_buffer(960) := X"0C020754";
        ram_buffer(961) := X"27A40010";
        ram_buffer(962) := X"10000015";
        ram_buffer(963) := X"00408021";
        ram_buffer(964) := X"3C02100C";
        ram_buffer(965) := X"24427BCC";
        ram_buffer(966) := X"1000FFAF";
        ram_buffer(967) := X"AF8281A4";
        ram_buffer(968) := X"0C021943";
        ram_buffer(969) := X"00000000";
        ram_buffer(970) := X"8F8481A0";
        ram_buffer(971) := X"00000000";
        ram_buffer(972) := X"1480FFD1";
        ram_buffer(973) := X"00408821";
        ram_buffer(974) := X"0C021948";
        ram_buffer(975) := X"00000000";
        ram_buffer(976) := X"00409821";
        ram_buffer(977) := X"8F8281A8";
        ram_buffer(978) := X"00000000";
        ram_buffer(979) := X"1040FFD3";
        ram_buffer(980) := X"00000000";
        ram_buffer(981) := X"0C0211E5";
        ram_buffer(982) := X"27A40010";
        ram_buffer(983) := X"00408021";
        ram_buffer(984) := X"8E020000";
        ram_buffer(985) := X"02002821";
        ram_buffer(986) := X"27A40010";
        ram_buffer(987) := X"0040F809";
        ram_buffer(988) := X"AE11000C";
        ram_buffer(989) := X"0C021D7F";
        ram_buffer(990) := X"27A40010";
        ram_buffer(991) := X"24070001";
        ram_buffer(992) := X"02803021";
        ram_buffer(993) := X"02402821";
        ram_buffer(994) := X"0C020196";
        ram_buffer(995) := X"27A40010";
        ram_buffer(996) := X"02602821";
        ram_buffer(997) := X"0C022264";
        ram_buffer(998) := X"27A40010";
        ram_buffer(999) := X"24050001";
        ram_buffer(1000) := X"0C021A9F";
        ram_buffer(1001) := X"27A40010";
        ram_buffer(1002) := X"8FA3002C";
        ram_buffer(1003) := X"8FA200E8";
        ram_buffer(1004) := X"00000000";
        ram_buffer(1005) := X"0043102B";
        ram_buffer(1006) := X"1040000F";
        ram_buffer(1007) := X"00000000";
        ram_buffer(1008) := X"8E020004";
        ram_buffer(1009) := X"02002821";
        ram_buffer(1010) := X"0040F809";
        ram_buffer(1011) := X"27A40010";
        ram_buffer(1012) := X"8E050010";
        ram_buffer(1013) := X"00403021";
        ram_buffer(1014) := X"0C021AD5";
        ram_buffer(1015) := X"27A40010";
        ram_buffer(1016) := X"8FA3002C";
        ram_buffer(1017) := X"8FA200E8";
        ram_buffer(1018) := X"00000000";
        ram_buffer(1019) := X"0043102B";
        ram_buffer(1020) := X"1440FFF3";
        ram_buffer(1021) := X"00000000";
        ram_buffer(1022) := X"8E020008";
        ram_buffer(1023) := X"02002821";
        ram_buffer(1024) := X"0040F809";
        ram_buffer(1025) := X"27A40010";
        ram_buffer(1026) := X"0C0219D5";
        ram_buffer(1027) := X"27A40010";
        ram_buffer(1028) := X"0C021993";
        ram_buffer(1029) := X"27A40010";
        ram_buffer(1030) := X"8F828098";
        ram_buffer(1031) := X"00000000";
        ram_buffer(1032) := X"8C430004";
        ram_buffer(1033) := X"00000000";
        ram_buffer(1034) := X"12230005";
        ram_buffer(1035) := X"00000000";
        ram_buffer(1036) := X"0C026DBB";
        ram_buffer(1037) := X"02202021";
        ram_buffer(1038) := X"8F828098";
        ram_buffer(1039) := X"00000000";
        ram_buffer(1040) := X"8C420008";
        ram_buffer(1041) := X"00000000";
        ram_buffer(1042) := X"12620003";
        ram_buffer(1043) := X"00000000";
        ram_buffer(1044) := X"0C026DBB";
        ram_buffer(1045) := X"02602021";
        ram_buffer(1046) := X"8FBF0214";
        ram_buffer(1047) := X"8FB40210";
        ram_buffer(1048) := X"8FB3020C";
        ram_buffer(1049) := X"8FB20208";
        ram_buffer(1050) := X"8FB10204";
        ram_buffer(1051) := X"8FB00200";
        ram_buffer(1052) := X"00001021";
        ram_buffer(1053) := X"03E00008";
        ram_buffer(1054) := X"27BD0218";
        ram_buffer(1055) := X"1200FFB5";
        ram_buffer(1056) := X"00000000";
        ram_buffer(1057) := X"8FA20010";
        ram_buffer(1058) := X"24040411";
        ram_buffer(1059) := X"8C430000";
        ram_buffer(1060) := X"AC440014";
        ram_buffer(1061) := X"0060F809";
        ram_buffer(1062) := X"27A40010";
        ram_buffer(1063) := X"AC11000C";
        ram_buffer(1064) := X"0000000D";
        ram_buffer(1065) := X"0C020E0C";
        ram_buffer(1066) := X"27A40010";
        ram_buffer(1067) := X"1000FFAC";
        ram_buffer(1068) := X"00408021";
        ram_buffer(1069) := X"0C0215F7";
        ram_buffer(1070) := X"27A40010";
        ram_buffer(1071) := X"1000FFA8";
        ram_buffer(1072) := X"00408021";
        ram_buffer(1073) := X"8F848098";
        ram_buffer(1074) := X"0C028350";
        ram_buffer(1075) := X"02202821";
        ram_buffer(1076) := X"00408021";
        ram_buffer(1077) := X"2402FFFF";
        ram_buffer(1078) := X"1602FF7A";
        ram_buffer(1079) := X"24050029";
        ram_buffer(1080) := X"8FA20010";
        ram_buffer(1081) := X"00000000";
        ram_buffer(1082) := X"8C430000";
        ram_buffer(1083) := X"27A40010";
        ram_buffer(1084) := X"0060F809";
        ram_buffer(1085) := X"AC450014";
        ram_buffer(1086) := X"02202821";
        ram_buffer(1087) := X"0C029D83";
        ram_buffer(1088) := X"2404FFFF";
        ram_buffer(1089) := X"1450FFDF";
        ram_buffer(1090) := X"00000000";
        ram_buffer(1091) := X"8FA20010";
        ram_buffer(1092) := X"24040410";
        ram_buffer(1093) := X"8C430000";
        ram_buffer(1094) := X"AC440014";
        ram_buffer(1095) := X"0060F809";
        ram_buffer(1096) := X"27A40010";
        ram_buffer(1097) := X"1000FF6E";
        ram_buffer(1098) := X"24020042";
        ram_buffer(1099) := X"8F828098";
        ram_buffer(1100) := X"8E070000";
        ram_buffer(1101) := X"8C44000C";
        ram_buffer(1102) := X"8F8681A4";
        ram_buffer(1103) := X"3C05100C";
        ram_buffer(1104) := X"0C027196";
        ram_buffer(1105) := X"24A57BF4";
        ram_buffer(1106) := X"0C026D37";
        ram_buffer(1107) := X"24040001";
        ram_buffer(1108) := X"8F828098";
        ram_buffer(1109) := X"8F8781A0";
        ram_buffer(1110) := X"8C44000C";
        ram_buffer(1111) := X"1000FFF6";
        ram_buffer(1112) := X"00000000";
        ram_buffer(1113) := X"8F828098";
        ram_buffer(1114) := X"8F8681A4";
        ram_buffer(1115) := X"8C44000C";
        ram_buffer(1116) := X"3C05100C";
        ram_buffer(1117) := X"0C027196";
        ram_buffer(1118) := X"24A57BD4";
        ram_buffer(1119) := X"0C02002A";
        ram_buffer(1120) := X"00000000";
        ram_buffer(1121) := X"03E00008";
        ram_buffer(1122) := X"00000000";
        ram_buffer(1123) := X"27BDFFE0";
        ram_buffer(1124) := X"8CA7000C";
        ram_buffer(1125) := X"8CA60020";
        ram_buffer(1126) := X"AFB20018";
        ram_buffer(1127) := X"00809021";
        ram_buffer(1128) := X"8CA40018";
        ram_buffer(1129) := X"AFB10014";
        ram_buffer(1130) := X"00A08821";
        ram_buffer(1131) := X"AFB00010";
        ram_buffer(1132) := X"AFBF001C";
        ram_buffer(1133) := X"8E300024";
        ram_buffer(1134) := X"0C0272E9";
        ram_buffer(1135) := X"24050001";
        ram_buffer(1136) := X"8E230020";
        ram_buffer(1137) := X"00000000";
        ram_buffer(1138) := X"10430007";
        ram_buffer(1139) := X"00000000";
        ram_buffer(1140) := X"8E420000";
        ram_buffer(1141) := X"2404002A";
        ram_buffer(1142) := X"8C430000";
        ram_buffer(1143) := X"AC440014";
        ram_buffer(1144) := X"0060F809";
        ram_buffer(1145) := X"02402021";
        ram_buffer(1146) := X"8E220010";
        ram_buffer(1147) := X"8E450018";
        ram_buffer(1148) := X"8C430000";
        ram_buffer(1149) := X"8E220018";
        ram_buffer(1150) := X"10A00016";
        ram_buffer(1151) := X"00000000";
        ram_buffer(1152) := X"00052040";
        ram_buffer(1153) := X"00852821";
        ram_buffer(1154) := X"00452821";
        ram_buffer(1155) := X"90440000";
        ram_buffer(1156) := X"24630003";
        ram_buffer(1157) := X"02042021";
        ram_buffer(1158) := X"90840000";
        ram_buffer(1159) := X"24420003";
        ram_buffer(1160) := X"A064FFFD";
        ram_buffer(1161) := X"9044FFFE";
        ram_buffer(1162) := X"00000000";
        ram_buffer(1163) := X"02042021";
        ram_buffer(1164) := X"90840000";
        ram_buffer(1165) := X"00000000";
        ram_buffer(1166) := X"A064FFFE";
        ram_buffer(1167) := X"9044FFFF";
        ram_buffer(1168) := X"00000000";
        ram_buffer(1169) := X"02042021";
        ram_buffer(1170) := X"90840000";
        ram_buffer(1171) := X"1445FFEF";
        ram_buffer(1172) := X"A064FFFF";
        ram_buffer(1173) := X"8FBF001C";
        ram_buffer(1174) := X"8FB20018";
        ram_buffer(1175) := X"8FB10014";
        ram_buffer(1176) := X"8FB00010";
        ram_buffer(1177) := X"24020001";
        ram_buffer(1178) := X"03E00008";
        ram_buffer(1179) := X"27BD0020";
        ram_buffer(1180) := X"27BDFFE0";
        ram_buffer(1181) := X"8CA7000C";
        ram_buffer(1182) := X"8CA60020";
        ram_buffer(1183) := X"AFB20018";
        ram_buffer(1184) := X"00809021";
        ram_buffer(1185) := X"8CA40018";
        ram_buffer(1186) := X"AFB10014";
        ram_buffer(1187) := X"00A08821";
        ram_buffer(1188) := X"AFB00010";
        ram_buffer(1189) := X"AFBF001C";
        ram_buffer(1190) := X"8E300024";
        ram_buffer(1191) := X"0C0272E9";
        ram_buffer(1192) := X"24050001";
        ram_buffer(1193) := X"8E230020";
        ram_buffer(1194) := X"00000000";
        ram_buffer(1195) := X"10430007";
        ram_buffer(1196) := X"2404002A";
        ram_buffer(1197) := X"8E420000";
        ram_buffer(1198) := X"00000000";
        ram_buffer(1199) := X"8C430000";
        ram_buffer(1200) := X"AC440014";
        ram_buffer(1201) := X"0060F809";
        ram_buffer(1202) := X"02402021";
        ram_buffer(1203) := X"8E220010";
        ram_buffer(1204) := X"8E460018";
        ram_buffer(1205) := X"8C440000";
        ram_buffer(1206) := X"8E220018";
        ram_buffer(1207) := X"10C0001C";
        ram_buffer(1208) := X"00000000";
        ram_buffer(1209) := X"00061840";
        ram_buffer(1210) := X"00663021";
        ram_buffer(1211) := X"00863021";
        ram_buffer(1212) := X"90430001";
        ram_buffer(1213) := X"90450000";
        ram_buffer(1214) := X"00031A00";
        ram_buffer(1215) := X"00651825";
        ram_buffer(1216) := X"02031821";
        ram_buffer(1217) := X"90630000";
        ram_buffer(1218) := X"24420006";
        ram_buffer(1219) := X"A0830000";
        ram_buffer(1220) := X"9043FFFD";
        ram_buffer(1221) := X"9045FFFC";
        ram_buffer(1222) := X"00031A00";
        ram_buffer(1223) := X"00651825";
        ram_buffer(1224) := X"02031821";
        ram_buffer(1225) := X"90630000";
        ram_buffer(1226) := X"24840003";
        ram_buffer(1227) := X"A083FFFE";
        ram_buffer(1228) := X"9043FFFF";
        ram_buffer(1229) := X"9045FFFE";
        ram_buffer(1230) := X"00031A00";
        ram_buffer(1231) := X"00651825";
        ram_buffer(1232) := X"02031821";
        ram_buffer(1233) := X"90630000";
        ram_buffer(1234) := X"1486FFE9";
        ram_buffer(1235) := X"A083FFFF";
        ram_buffer(1236) := X"8FBF001C";
        ram_buffer(1237) := X"8FB20018";
        ram_buffer(1238) := X"8FB10014";
        ram_buffer(1239) := X"8FB00010";
        ram_buffer(1240) := X"24020001";
        ram_buffer(1241) := X"03E00008";
        ram_buffer(1242) := X"27BD0020";
        ram_buffer(1243) := X"27BDFFE0";
        ram_buffer(1244) := X"8CA7000C";
        ram_buffer(1245) := X"8CA60020";
        ram_buffer(1246) := X"AFB20018";
        ram_buffer(1247) := X"00809021";
        ram_buffer(1248) := X"8CA40018";
        ram_buffer(1249) := X"AFB10014";
        ram_buffer(1250) := X"00A08821";
        ram_buffer(1251) := X"AFB00010";
        ram_buffer(1252) := X"AFBF001C";
        ram_buffer(1253) := X"8E300024";
        ram_buffer(1254) := X"0C0272E9";
        ram_buffer(1255) := X"24050001";
        ram_buffer(1256) := X"8E230020";
        ram_buffer(1257) := X"00000000";
        ram_buffer(1258) := X"10430007";
        ram_buffer(1259) := X"2404002A";
        ram_buffer(1260) := X"8E420000";
        ram_buffer(1261) := X"00000000";
        ram_buffer(1262) := X"8C430000";
        ram_buffer(1263) := X"AC440014";
        ram_buffer(1264) := X"0060F809";
        ram_buffer(1265) := X"02402021";
        ram_buffer(1266) := X"8E220010";
        ram_buffer(1267) := X"8E430018";
        ram_buffer(1268) := X"8C420000";
        ram_buffer(1269) := X"8E240018";
        ram_buffer(1270) := X"10600008";
        ram_buffer(1271) := X"00432821";
        ram_buffer(1272) := X"24840001";
        ram_buffer(1273) := X"9083FFFF";
        ram_buffer(1274) := X"24420001";
        ram_buffer(1275) := X"02031821";
        ram_buffer(1276) := X"90630000";
        ram_buffer(1277) := X"1445FFFA";
        ram_buffer(1278) := X"A043FFFF";
        ram_buffer(1279) := X"8FBF001C";
        ram_buffer(1280) := X"8FB20018";
        ram_buffer(1281) := X"8FB10014";
        ram_buffer(1282) := X"8FB00010";
        ram_buffer(1283) := X"24020001";
        ram_buffer(1284) := X"03E00008";
        ram_buffer(1285) := X"27BD0020";
        ram_buffer(1286) := X"27BDFFE0";
        ram_buffer(1287) := X"8CA7000C";
        ram_buffer(1288) := X"8CA60020";
        ram_buffer(1289) := X"AFB20018";
        ram_buffer(1290) := X"00809021";
        ram_buffer(1291) := X"8CA40018";
        ram_buffer(1292) := X"AFB10014";
        ram_buffer(1293) := X"00A08821";
        ram_buffer(1294) := X"AFB00010";
        ram_buffer(1295) := X"AFBF001C";
        ram_buffer(1296) := X"8E300024";
        ram_buffer(1297) := X"0C0272E9";
        ram_buffer(1298) := X"24050001";
        ram_buffer(1299) := X"8E230020";
        ram_buffer(1300) := X"00000000";
        ram_buffer(1301) := X"10430007";
        ram_buffer(1302) := X"2404002A";
        ram_buffer(1303) := X"8E420000";
        ram_buffer(1304) := X"00000000";
        ram_buffer(1305) := X"8C430000";
        ram_buffer(1306) := X"AC440014";
        ram_buffer(1307) := X"0060F809";
        ram_buffer(1308) := X"02402021";
        ram_buffer(1309) := X"8E230010";
        ram_buffer(1310) := X"8E420018";
        ram_buffer(1311) := X"8C630000";
        ram_buffer(1312) := X"8E240018";
        ram_buffer(1313) := X"1040000B";
        ram_buffer(1314) := X"00623021";
        ram_buffer(1315) := X"90850000";
        ram_buffer(1316) := X"24840002";
        ram_buffer(1317) := X"9082FFFF";
        ram_buffer(1318) := X"24630001";
        ram_buffer(1319) := X"00021200";
        ram_buffer(1320) := X"00451025";
        ram_buffer(1321) := X"02021021";
        ram_buffer(1322) := X"90420000";
        ram_buffer(1323) := X"1466FFF7";
        ram_buffer(1324) := X"A062FFFF";
        ram_buffer(1325) := X"8FBF001C";
        ram_buffer(1326) := X"8FB20018";
        ram_buffer(1327) := X"8FB10014";
        ram_buffer(1328) := X"8FB00010";
        ram_buffer(1329) := X"24020001";
        ram_buffer(1330) := X"03E00008";
        ram_buffer(1331) := X"27BD0020";
        ram_buffer(1332) := X"27BDFFE0";
        ram_buffer(1333) := X"8CA7000C";
        ram_buffer(1334) := X"8CA60020";
        ram_buffer(1335) := X"AFB10018";
        ram_buffer(1336) := X"00808821";
        ram_buffer(1337) := X"8CA40018";
        ram_buffer(1338) := X"AFB00014";
        ram_buffer(1339) := X"00A08021";
        ram_buffer(1340) := X"AFBF001C";
        ram_buffer(1341) := X"0C0272E9";
        ram_buffer(1342) := X"24050001";
        ram_buffer(1343) := X"8E030020";
        ram_buffer(1344) := X"00000000";
        ram_buffer(1345) := X"10430007";
        ram_buffer(1346) := X"00000000";
        ram_buffer(1347) := X"8E220000";
        ram_buffer(1348) := X"2404002A";
        ram_buffer(1349) := X"8C430000";
        ram_buffer(1350) := X"AC440014";
        ram_buffer(1351) := X"0060F809";
        ram_buffer(1352) := X"02202021";
        ram_buffer(1353) := X"8FBF001C";
        ram_buffer(1354) := X"8FB10018";
        ram_buffer(1355) := X"8FB00014";
        ram_buffer(1356) := X"24020001";
        ram_buffer(1357) := X"03E00008";
        ram_buffer(1358) := X"27BD0020";
        ram_buffer(1359) := X"27BDFFD0";
        ram_buffer(1360) := X"AFB60028";
        ram_buffer(1361) := X"AFB50024";
        ram_buffer(1362) := X"AFB40020";
        ram_buffer(1363) := X"AFB3001C";
        ram_buffer(1364) := X"AFB20018";
        ram_buffer(1365) := X"AFB10014";
        ram_buffer(1366) := X"AFB00010";
        ram_buffer(1367) := X"AFBF002C";
        ram_buffer(1368) := X"0080A021";
        ram_buffer(1369) := X"00A08021";
        ram_buffer(1370) := X"24120020";
        ram_buffer(1371) := X"2415000D";
        ram_buffer(1372) := X"2416000A";
        ram_buffer(1373) := X"2413FFFF";
        ram_buffer(1374) := X"24110023";
        ram_buffer(1375) := X"8E020004";
        ram_buffer(1376) := X"00000000";
        ram_buffer(1377) := X"2442FFFF";
        ram_buffer(1378) := X"04400057";
        ram_buffer(1379) := X"AE020004";
        ram_buffer(1380) := X"8E030000";
        ram_buffer(1381) := X"00000000";
        ram_buffer(1382) := X"24640001";
        ram_buffer(1383) := X"AE040000";
        ram_buffer(1384) := X"90630000";
        ram_buffer(1385) := X"00000000";
        ram_buffer(1386) := X"10710043";
        ram_buffer(1387) := X"2442FFFF";
        ram_buffer(1388) := X"1072FFF2";
        ram_buffer(1389) := X"2462FFF7";
        ram_buffer(1390) := X"2C420002";
        ram_buffer(1391) := X"1440FFEF";
        ram_buffer(1392) := X"00000000";
        ram_buffer(1393) := X"1075FFED";
        ram_buffer(1394) := X"00000000";
        ram_buffer(1395) := X"2471FFD0";
        ram_buffer(1396) := X"2E22000A";
        ram_buffer(1397) := X"10400052";
        ram_buffer(1398) := X"02209021";
        ram_buffer(1399) := X"10000004";
        ram_buffer(1400) := X"24110023";
        ram_buffer(1401) := X"10800056";
        ram_buffer(1402) := X"00000000";
        ram_buffer(1403) := X"00629021";
        ram_buffer(1404) := X"8E020004";
        ram_buffer(1405) := X"00000000";
        ram_buffer(1406) := X"2442FFFF";
        ram_buffer(1407) := X"0440005B";
        ram_buffer(1408) := X"AE020004";
        ram_buffer(1409) := X"8E020000";
        ram_buffer(1410) := X"00000000";
        ram_buffer(1411) := X"24430001";
        ram_buffer(1412) := X"AE030000";
        ram_buffer(1413) := X"90420000";
        ram_buffer(1414) := X"00122040";
        ram_buffer(1415) := X"001218C0";
        ram_buffer(1416) := X"00831821";
        ram_buffer(1417) := X"2445FFD0";
        ram_buffer(1418) := X"2463FFD0";
        ram_buffer(1419) := X"1451FFED";
        ram_buffer(1420) := X"2CA4000A";
        ram_buffer(1421) := X"8E020004";
        ram_buffer(1422) := X"2411000A";
        ram_buffer(1423) := X"10000009";
        ram_buffer(1424) := X"2413FFFF";
        ram_buffer(1425) := X"8E030000";
        ram_buffer(1426) := X"00000000";
        ram_buffer(1427) := X"24640001";
        ram_buffer(1428) := X"AE040000";
        ram_buffer(1429) := X"90630000";
        ram_buffer(1430) := X"00000000";
        ram_buffer(1431) := X"10710038";
        ram_buffer(1432) := X"00000000";
        ram_buffer(1433) := X"2442FFFF";
        ram_buffer(1434) := X"0441FFF6";
        ram_buffer(1435) := X"AE020004";
        ram_buffer(1436) := X"8F848098";
        ram_buffer(1437) := X"0C028350";
        ram_buffer(1438) := X"02002821";
        ram_buffer(1439) := X"10510030";
        ram_buffer(1440) := X"00000000";
        ram_buffer(1441) := X"1053002E";
        ram_buffer(1442) := X"00000000";
        ram_buffer(1443) := X"8E020004";
        ram_buffer(1444) := X"1000FFF5";
        ram_buffer(1445) := X"2442FFFF";
        ram_buffer(1446) := X"8E030000";
        ram_buffer(1447) := X"00000000";
        ram_buffer(1448) := X"24640001";
        ram_buffer(1449) := X"AE040000";
        ram_buffer(1450) := X"90630000";
        ram_buffer(1451) := X"00000000";
        ram_buffer(1452) := X"1076FFB2";
        ram_buffer(1453) := X"2442FFFF";
        ram_buffer(1454) := X"0441FFF7";
        ram_buffer(1455) := X"AE020004";
        ram_buffer(1456) := X"8F848098";
        ram_buffer(1457) := X"0C028350";
        ram_buffer(1458) := X"02002821";
        ram_buffer(1459) := X"1056FFAB";
        ram_buffer(1460) := X"00000000";
        ram_buffer(1461) := X"1053000B";
        ram_buffer(1462) := X"00000000";
        ram_buffer(1463) := X"8E020004";
        ram_buffer(1464) := X"1000FFF5";
        ram_buffer(1465) := X"2442FFFF";
        ram_buffer(1466) := X"8F848098";
        ram_buffer(1467) := X"0C028350";
        ram_buffer(1468) := X"02002821";
        ram_buffer(1469) := X"1051FFF9";
        ram_buffer(1470) := X"00401821";
        ram_buffer(1471) := X"1453FFAC";
        ram_buffer(1472) := X"00000000";
        ram_buffer(1473) := X"8E820000";
        ram_buffer(1474) := X"2404002A";
        ram_buffer(1475) := X"8C430000";
        ram_buffer(1476) := X"AC440014";
        ram_buffer(1477) := X"0060F809";
        ram_buffer(1478) := X"02802021";
        ram_buffer(1479) := X"2411FFCF";
        ram_buffer(1480) := X"8E820000";
        ram_buffer(1481) := X"24040402";
        ram_buffer(1482) := X"8C430000";
        ram_buffer(1483) := X"AC440014";
        ram_buffer(1484) := X"0060F809";
        ram_buffer(1485) := X"02802021";
        ram_buffer(1486) := X"1000FFA8";
        ram_buffer(1487) := X"02209021";
        ram_buffer(1488) := X"8FBF002C";
        ram_buffer(1489) := X"02401021";
        ram_buffer(1490) := X"8FB60028";
        ram_buffer(1491) := X"8FB50024";
        ram_buffer(1492) := X"8FB40020";
        ram_buffer(1493) := X"8FB3001C";
        ram_buffer(1494) := X"8FB20018";
        ram_buffer(1495) := X"8FB10014";
        ram_buffer(1496) := X"8FB00010";
        ram_buffer(1497) := X"03E00008";
        ram_buffer(1498) := X"27BD0030";
        ram_buffer(1499) := X"8F848098";
        ram_buffer(1500) := X"0C028350";
        ram_buffer(1501) := X"02002821";
        ram_buffer(1502) := X"1000FFA8";
        ram_buffer(1503) := X"00122040";
        ram_buffer(1504) := X"27BDFFD0";
        ram_buffer(1505) := X"AFB10018";
        ram_buffer(1506) := X"00A08821";
        ram_buffer(1507) := X"8CA5000C";
        ram_buffer(1508) := X"AFB00014";
        ram_buffer(1509) := X"8CA20004";
        ram_buffer(1510) := X"AFBF002C";
        ram_buffer(1511) := X"2442FFFF";
        ram_buffer(1512) := X"AFB50028";
        ram_buffer(1513) := X"AFB40024";
        ram_buffer(1514) := X"AFB30020";
        ram_buffer(1515) := X"AFB2001C";
        ram_buffer(1516) := X"00808021";
        ram_buffer(1517) := X"0440010E";
        ram_buffer(1518) := X"ACA20004";
        ram_buffer(1519) := X"8CA20000";
        ram_buffer(1520) := X"00000000";
        ram_buffer(1521) := X"24430001";
        ram_buffer(1522) := X"ACA30000";
        ram_buffer(1523) := X"90420000";
        ram_buffer(1524) := X"00000000";
        ram_buffer(1525) := X"38420050";
        ram_buffer(1526) := X"0002102B";
        ram_buffer(1527) := X"144000D0";
        ram_buffer(1528) := X"24040403";
        ram_buffer(1529) := X"8E25000C";
        ram_buffer(1530) := X"00000000";
        ram_buffer(1531) := X"8CA20004";
        ram_buffer(1532) := X"00000000";
        ram_buffer(1533) := X"2442FFFF";
        ram_buffer(1534) := X"044000D6";
        ram_buffer(1535) := X"ACA20004";
        ram_buffer(1536) := X"8CA20000";
        ram_buffer(1537) := X"00000000";
        ram_buffer(1538) := X"24430001";
        ram_buffer(1539) := X"ACA30000";
        ram_buffer(1540) := X"90540000";
        ram_buffer(1541) := X"0C02054F";
        ram_buffer(1542) := X"02002021";
        ram_buffer(1543) := X"8E25000C";
        ram_buffer(1544) := X"02002021";
        ram_buffer(1545) := X"0C02054F";
        ram_buffer(1546) := X"00409821";
        ram_buffer(1547) := X"8E25000C";
        ram_buffer(1548) := X"02002021";
        ram_buffer(1549) := X"0C02054F";
        ram_buffer(1550) := X"0040A821";
        ram_buffer(1551) := X"12600003";
        ram_buffer(1552) := X"00409021";
        ram_buffer(1553) := X"16A0002E";
        ram_buffer(1554) := X"00000000";
        ram_buffer(1555) := X"8E020000";
        ram_buffer(1556) := X"24040403";
        ram_buffer(1557) := X"8C430000";
        ram_buffer(1558) := X"AC440014";
        ram_buffer(1559) := X"0060F809";
        ram_buffer(1560) := X"02002021";
        ram_buffer(1561) := X"24020008";
        ram_buffer(1562) := X"AE020030";
        ram_buffer(1563) := X"24020033";
        ram_buffer(1564) := X"AE130018";
        ram_buffer(1565) := X"12820029";
        ram_buffer(1566) := X"AE15001C";
        ram_buffer(1567) := X"2A820034";
        ram_buffer(1568) := X"14400092";
        ram_buffer(1569) := X"24020035";
        ram_buffer(1570) := X"1282004E";
        ram_buffer(1571) := X"24020036";
        ram_buffer(1572) := X"168200B6";
        ram_buffer(1573) := X"24030003";
        ram_buffer(1574) := X"8E020000";
        ram_buffer(1575) := X"AE030020";
        ram_buffer(1576) := X"24030002";
        ram_buffer(1577) := X"AE030024";
        ram_buffer(1578) := X"AC530018";
        ram_buffer(1579) := X"8E030000";
        ram_buffer(1580) := X"24040406";
        ram_buffer(1581) := X"AC440014";
        ram_buffer(1582) := X"AC75001C";
        ram_buffer(1583) := X"8E020000";
        ram_buffer(1584) := X"24050001";
        ram_buffer(1585) := X"8C420004";
        ram_buffer(1586) := X"00000000";
        ram_buffer(1587) := X"0040F809";
        ram_buffer(1588) := X"02002021";
        ram_buffer(1589) := X"2E420100";
        ram_buffer(1590) := X"104000C2";
        ram_buffer(1591) := X"3C021008";
        ram_buffer(1592) := X"240200FF";
        ram_buffer(1593) := X"124200C8";
        ram_buffer(1594) := X"3C021008";
        ram_buffer(1595) := X"2442118C";
        ram_buffer(1596) := X"AE220004";
        ram_buffer(1597) := X"24140001";
        ram_buffer(1598) := X"1000004B";
        ram_buffer(1599) := X"0000A821";
        ram_buffer(1600) := X"1040FFD2";
        ram_buffer(1601) := X"24020008";
        ram_buffer(1602) := X"AE020030";
        ram_buffer(1603) := X"24020033";
        ram_buffer(1604) := X"AE130018";
        ram_buffer(1605) := X"1682FFD9";
        ram_buffer(1606) := X"AE15001C";
        ram_buffer(1607) := X"8E020000";
        ram_buffer(1608) := X"24030003";
        ram_buffer(1609) := X"AE030020";
        ram_buffer(1610) := X"24030002";
        ram_buffer(1611) := X"AE030024";
        ram_buffer(1612) := X"AC530018";
        ram_buffer(1613) := X"8E030000";
        ram_buffer(1614) := X"24040407";
        ram_buffer(1615) := X"AC440014";
        ram_buffer(1616) := X"AC75001C";
        ram_buffer(1617) := X"8E020000";
        ram_buffer(1618) := X"24050001";
        ram_buffer(1619) := X"8C420004";
        ram_buffer(1620) := X"00000000";
        ram_buffer(1621) := X"0040F809";
        ram_buffer(1622) := X"02002021";
        ram_buffer(1623) := X"3C021008";
        ram_buffer(1624) := X"24421C20";
        ram_buffer(1625) := X"AE220004";
        ram_buffer(1626) := X"24140001";
        ram_buffer(1627) := X"8E060020";
        ram_buffer(1628) := X"8E020004";
        ram_buffer(1629) := X"02660018";
        ram_buffer(1630) := X"8C420008";
        ram_buffer(1631) := X"24070001";
        ram_buffer(1632) := X"24050001";
        ram_buffer(1633) := X"00003012";
        ram_buffer(1634) := X"0040F809";
        ram_buffer(1635) := X"02002021";
        ram_buffer(1636) := X"AE220010";
        ram_buffer(1637) := X"24020001";
        ram_buffer(1638) := X"16800034";
        ram_buffer(1639) := X"AE220014";
        ram_buffer(1640) := X"8FBF002C";
        ram_buffer(1641) := X"8FB50028";
        ram_buffer(1642) := X"8FB40024";
        ram_buffer(1643) := X"8FB30020";
        ram_buffer(1644) := X"8FB2001C";
        ram_buffer(1645) := X"8FB10018";
        ram_buffer(1646) := X"8FB00014";
        ram_buffer(1647) := X"03E00008";
        ram_buffer(1648) := X"27BD0030";
        ram_buffer(1649) := X"8E020000";
        ram_buffer(1650) := X"24030001";
        ram_buffer(1651) := X"AE030020";
        ram_buffer(1652) := X"AE030024";
        ram_buffer(1653) := X"AC530018";
        ram_buffer(1654) := X"8E030000";
        ram_buffer(1655) := X"24040404";
        ram_buffer(1656) := X"AC440014";
        ram_buffer(1657) := X"AC75001C";
        ram_buffer(1658) := X"8E020000";
        ram_buffer(1659) := X"24050001";
        ram_buffer(1660) := X"8C420004";
        ram_buffer(1661) := X"00000000";
        ram_buffer(1662) := X"0040F809";
        ram_buffer(1663) := X"02002021";
        ram_buffer(1664) := X"2E420100";
        ram_buffer(1665) := X"1040006F";
        ram_buffer(1666) := X"3C021008";
        ram_buffer(1667) := X"240200FF";
        ram_buffer(1668) := X"1242007D";
        ram_buffer(1669) := X"3C021008";
        ram_buffer(1670) := X"2442136C";
        ram_buffer(1671) := X"AE220004";
        ram_buffer(1672) := X"24140001";
        ram_buffer(1673) := X"0000A821";
        ram_buffer(1674) := X"8E060020";
        ram_buffer(1675) := X"8E020004";
        ram_buffer(1676) := X"02660018";
        ram_buffer(1677) := X"8C420000";
        ram_buffer(1678) := X"24050001";
        ram_buffer(1679) := X"02002021";
        ram_buffer(1680) := X"00003012";
        ram_buffer(1681) := X"0040F809";
        ram_buffer(1682) := X"AE260020";
        ram_buffer(1683) := X"12A0FFC7";
        ram_buffer(1684) := X"AE220018";
        ram_buffer(1685) := X"2623001C";
        ram_buffer(1686) := X"AE22001C";
        ram_buffer(1687) := X"24020001";
        ram_buffer(1688) := X"AE230010";
        ram_buffer(1689) := X"1280FFCE";
        ram_buffer(1690) := X"AE220014";
        ram_buffer(1691) := X"8E020004";
        ram_buffer(1692) := X"26530001";
        ram_buffer(1693) := X"8C420000";
        ram_buffer(1694) := X"02603021";
        ram_buffer(1695) := X"24050001";
        ram_buffer(1696) := X"0040F809";
        ram_buffer(1697) := X"02002021";
        ram_buffer(1698) := X"AE220024";
        ram_buffer(1699) := X"0640FFC4";
        ram_buffer(1700) := X"00121842";
        ram_buffer(1701) := X"10000002";
        ram_buffer(1702) := X"00002021";
        ram_buffer(1703) := X"8E220024";
        ram_buffer(1704) := X"16400002";
        ram_buffer(1705) := X"0072001B";
        ram_buffer(1706) := X"0007000D";
        ram_buffer(1707) := X"00441021";
        ram_buffer(1708) := X"24840001";
        ram_buffer(1709) := X"246300FF";
        ram_buffer(1710) := X"00002812";
        ram_buffer(1711) := X"1493FFF7";
        ram_buffer(1712) := X"A0450000";
        ram_buffer(1713) := X"1000FFB6";
        ram_buffer(1714) := X"00000000";
        ram_buffer(1715) := X"24020032";
        ram_buffer(1716) := X"16820026";
        ram_buffer(1717) := X"24030001";
        ram_buffer(1718) := X"8E020000";
        ram_buffer(1719) := X"AE030020";
        ram_buffer(1720) := X"AE030024";
        ram_buffer(1721) := X"AC530018";
        ram_buffer(1722) := X"8E030000";
        ram_buffer(1723) := X"24040405";
        ram_buffer(1724) := X"AC440014";
        ram_buffer(1725) := X"AC75001C";
        ram_buffer(1726) := X"8E020000";
        ram_buffer(1727) := X"24050001";
        ram_buffer(1728) := X"8C420004";
        ram_buffer(1729) := X"00000000";
        ram_buffer(1730) := X"0040F809";
        ram_buffer(1731) := X"02002021";
        ram_buffer(1732) := X"3C021008";
        ram_buffer(1733) := X"24421CD0";
        ram_buffer(1734) := X"1000FF93";
        ram_buffer(1735) := X"AE220004";
        ram_buffer(1736) := X"8E020000";
        ram_buffer(1737) := X"00000000";
        ram_buffer(1738) := X"8C430000";
        ram_buffer(1739) := X"AC440014";
        ram_buffer(1740) := X"0060F809";
        ram_buffer(1741) := X"02002021";
        ram_buffer(1742) := X"8E25000C";
        ram_buffer(1743) := X"00000000";
        ram_buffer(1744) := X"8CA20004";
        ram_buffer(1745) := X"00000000";
        ram_buffer(1746) := X"2442FFFF";
        ram_buffer(1747) := X"0441FF2C";
        ram_buffer(1748) := X"ACA20004";
        ram_buffer(1749) := X"8F848098";
        ram_buffer(1750) := X"0C028350";
        ram_buffer(1751) := X"00000000";
        ram_buffer(1752) := X"8E25000C";
        ram_buffer(1753) := X"1000FF2B";
        ram_buffer(1754) := X"0040A021";
        ram_buffer(1755) := X"8E020000";
        ram_buffer(1756) := X"24040403";
        ram_buffer(1757) := X"8C430000";
        ram_buffer(1758) := X"AC440014";
        ram_buffer(1759) := X"0060F809";
        ram_buffer(1760) := X"02002021";
        ram_buffer(1761) := X"8E060020";
        ram_buffer(1762) := X"2E420100";
        ram_buffer(1763) := X"02660018";
        ram_buffer(1764) := X"2C420001";
        ram_buffer(1765) := X"24420001";
        ram_buffer(1766) := X"00003012";
        ram_buffer(1767) := X"8E030004";
        ram_buffer(1768) := X"24050001";
        ram_buffer(1769) := X"00460018";
        ram_buffer(1770) := X"8C630000";
        ram_buffer(1771) := X"02002021";
        ram_buffer(1772) := X"00003012";
        ram_buffer(1773) := X"0060F809";
        ram_buffer(1774) := X"AE260020";
        ram_buffer(1775) := X"1000FF6A";
        ram_buffer(1776) := X"AE220018";
        ram_buffer(1777) := X"24421418";
        ram_buffer(1778) := X"AE220004";
        ram_buffer(1779) := X"8E060020";
        ram_buffer(1780) := X"00000000";
        ram_buffer(1781) := X"02660018";
        ram_buffer(1782) := X"00003012";
        ram_buffer(1783) := X"1000FFEF";
        ram_buffer(1784) := X"24020002";
        ram_buffer(1785) := X"24421270";
        ram_buffer(1786) := X"1000FFF8";
        ram_buffer(1787) := X"AE220004";
        ram_buffer(1788) := X"8F848098";
        ram_buffer(1789) := X"0C028350";
        ram_buffer(1790) := X"00000000";
        ram_buffer(1791) := X"38420050";
        ram_buffer(1792) := X"1000FEF6";
        ram_buffer(1793) := X"0002102B";
        ram_buffer(1794) := X"3C021008";
        ram_buffer(1795) := X"244214D0";
        ram_buffer(1796) := X"AE220004";
        ram_buffer(1797) := X"0000A021";
        ram_buffer(1798) := X"1000FF83";
        ram_buffer(1799) := X"24150001";
        ram_buffer(1800) := X"27BDFFD8";
        ram_buffer(1801) := X"8CA20010";
        ram_buffer(1802) := X"AFB10014";
        ram_buffer(1803) := X"8C910018";
        ram_buffer(1804) := X"AFB40020";
        ram_buffer(1805) := X"AFB3001C";
        ram_buffer(1806) := X"AFB00010";
        ram_buffer(1807) := X"AFBF0024";
        ram_buffer(1808) := X"AFB20018";
        ram_buffer(1809) := X"8CB4000C";
        ram_buffer(1810) := X"8CB30024";
        ram_buffer(1811) := X"8C500000";
        ram_buffer(1812) := X"12200016";
        ram_buffer(1813) := X"00809021";
        ram_buffer(1814) := X"02802821";
        ram_buffer(1815) := X"0C02054F";
        ram_buffer(1816) := X"02402021";
        ram_buffer(1817) := X"02621021";
        ram_buffer(1818) := X"90420000";
        ram_buffer(1819) := X"02802821";
        ram_buffer(1820) := X"A2020000";
        ram_buffer(1821) := X"0C02054F";
        ram_buffer(1822) := X"02402021";
        ram_buffer(1823) := X"02621021";
        ram_buffer(1824) := X"90420000";
        ram_buffer(1825) := X"02802821";
        ram_buffer(1826) := X"A2020001";
        ram_buffer(1827) := X"0C02054F";
        ram_buffer(1828) := X"02402021";
        ram_buffer(1829) := X"02621021";
        ram_buffer(1830) := X"90420000";
        ram_buffer(1831) := X"26100003";
        ram_buffer(1832) := X"2631FFFF";
        ram_buffer(1833) := X"1620FFEC";
        ram_buffer(1834) := X"A202FFFF";
        ram_buffer(1835) := X"8FBF0024";
        ram_buffer(1836) := X"8FB40020";
        ram_buffer(1837) := X"8FB3001C";
        ram_buffer(1838) := X"8FB20018";
        ram_buffer(1839) := X"8FB10014";
        ram_buffer(1840) := X"8FB00010";
        ram_buffer(1841) := X"24020001";
        ram_buffer(1842) := X"03E00008";
        ram_buffer(1843) := X"27BD0028";
        ram_buffer(1844) := X"27BDFFD8";
        ram_buffer(1845) := X"8CA20010";
        ram_buffer(1846) := X"AFB00010";
        ram_buffer(1847) := X"8C900018";
        ram_buffer(1848) := X"AFB40020";
        ram_buffer(1849) := X"AFB3001C";
        ram_buffer(1850) := X"AFB10014";
        ram_buffer(1851) := X"AFBF0024";
        ram_buffer(1852) := X"AFB20018";
        ram_buffer(1853) := X"8CB4000C";
        ram_buffer(1854) := X"8CB30024";
        ram_buffer(1855) := X"8C510000";
        ram_buffer(1856) := X"1200000A";
        ram_buffer(1857) := X"00809021";
        ram_buffer(1858) := X"02802821";
        ram_buffer(1859) := X"0C02054F";
        ram_buffer(1860) := X"02402021";
        ram_buffer(1861) := X"02621021";
        ram_buffer(1862) := X"90420000";
        ram_buffer(1863) := X"26310001";
        ram_buffer(1864) := X"2610FFFF";
        ram_buffer(1865) := X"1600FFF8";
        ram_buffer(1866) := X"A222FFFF";
        ram_buffer(1867) := X"8FBF0024";
        ram_buffer(1868) := X"8FB40020";
        ram_buffer(1869) := X"8FB3001C";
        ram_buffer(1870) := X"8FB20018";
        ram_buffer(1871) := X"8FB10014";
        ram_buffer(1872) := X"8FB00010";
        ram_buffer(1873) := X"24020001";
        ram_buffer(1874) := X"03E00008";
        ram_buffer(1875) := X"27BD0028";
        ram_buffer(1876) := X"8C820004";
        ram_buffer(1877) := X"27BDFFE8";
        ram_buffer(1878) := X"8C420000";
        ram_buffer(1879) := X"24060028";
        ram_buffer(1880) := X"AFBF0014";
        ram_buffer(1881) := X"0040F809";
        ram_buffer(1882) := X"24050001";
        ram_buffer(1883) := X"3C031008";
        ram_buffer(1884) := X"24631780";
        ram_buffer(1885) := X"AC430000";
        ram_buffer(1886) := X"8FBF0014";
        ram_buffer(1887) := X"3C031008";
        ram_buffer(1888) := X"24631184";
        ram_buffer(1889) := X"AC430008";
        ram_buffer(1890) := X"03E00008";
        ram_buffer(1891) := X"27BD0018";
        ram_buffer(1892) := X"8CA20170";
        ram_buffer(1893) := X"27BDFFD8";
        ram_buffer(1894) := X"30430007";
        ram_buffer(1895) := X"AFB20020";
        ram_buffer(1896) := X"00809021";
        ram_buffer(1897) := X"24040002";
        ram_buffer(1898) := X"AFB1001C";
        ram_buffer(1899) := X"AFB00018";
        ram_buffer(1900) := X"AFBF0024";
        ram_buffer(1901) := X"8CB0001C";
        ram_buffer(1902) := X"10640037";
        ram_buffer(1903) := X"00A08821";
        ram_buffer(1904) := X"28640003";
        ram_buffer(1905) := X"1480003C";
        ram_buffer(1906) := X"24040004";
        ram_buffer(1907) := X"14640030";
        ram_buffer(1908) := X"24040006";
        ram_buffer(1909) := X"8CA60174";
        ram_buffer(1910) := X"000210C2";
        ram_buffer(1911) := X"00463021";
        ram_buffer(1912) := X"8E420004";
        ram_buffer(1913) := X"8E25016C";
        ram_buffer(1914) := X"AFA00010";
        ram_buffer(1915) := X"8C42001C";
        ram_buffer(1916) := X"02402021";
        ram_buffer(1917) := X"0040F809";
        ram_buffer(1918) := X"24070001";
        ram_buffer(1919) := X"8C430000";
        ram_buffer(1920) := X"8E440018";
        ram_buffer(1921) := X"8E220010";
        ram_buffer(1922) := X"00000000";
        ram_buffer(1923) := X"8C420000";
        ram_buffer(1924) := X"10800015";
        ram_buffer(1925) := X"00643021";
        ram_buffer(1926) := X"24630001";
        ram_buffer(1927) := X"9065FFFF";
        ram_buffer(1928) := X"8E040000";
        ram_buffer(1929) := X"24420003";
        ram_buffer(1930) := X"00852021";
        ram_buffer(1931) := X"90840000";
        ram_buffer(1932) := X"00000000";
        ram_buffer(1933) := X"A044FFFD";
        ram_buffer(1934) := X"8E040004";
        ram_buffer(1935) := X"00000000";
        ram_buffer(1936) := X"00852021";
        ram_buffer(1937) := X"90840000";
        ram_buffer(1938) := X"00000000";
        ram_buffer(1939) := X"A044FFFE";
        ram_buffer(1940) := X"8E040008";
        ram_buffer(1941) := X"00000000";
        ram_buffer(1942) := X"00852021";
        ram_buffer(1943) := X"90840000";
        ram_buffer(1944) := X"1466FFED";
        ram_buffer(1945) := X"A044FFFF";
        ram_buffer(1946) := X"8E220170";
        ram_buffer(1947) := X"8FBF0024";
        ram_buffer(1948) := X"24420001";
        ram_buffer(1949) := X"AE220170";
        ram_buffer(1950) := X"8FB20020";
        ram_buffer(1951) := X"8FB1001C";
        ram_buffer(1952) := X"8FB00018";
        ram_buffer(1953) := X"24020001";
        ram_buffer(1954) := X"03E00008";
        ram_buffer(1955) := X"27BD0028";
        ram_buffer(1956) := X"14640005";
        ram_buffer(1957) := X"00000000";
        ram_buffer(1958) := X"8E260178";
        ram_buffer(1959) := X"00021082";
        ram_buffer(1960) := X"1000FFCF";
        ram_buffer(1961) := X"00463021";
        ram_buffer(1962) := X"8E26017C";
        ram_buffer(1963) := X"00021042";
        ram_buffer(1964) := X"1000FFCB";
        ram_buffer(1965) := X"00463021";
        ram_buffer(1966) := X"1460FFFB";
        ram_buffer(1967) := X"00000000";
        ram_buffer(1968) := X"1000FFC7";
        ram_buffer(1969) := X"000230C2";
        ram_buffer(1970) := X"03E00008";
        ram_buffer(1971) := X"00000000";
        ram_buffer(1972) := X"18A00080";
        ram_buffer(1973) := X"00000000";
        ram_buffer(1974) := X"27BDFFC8";
        ram_buffer(1975) := X"AFB6002C";
        ram_buffer(1976) := X"AFB50028";
        ram_buffer(1977) := X"AFB30020";
        ram_buffer(1978) := X"AFB2001C";
        ram_buffer(1979) := X"AFB10018";
        ram_buffer(1980) := X"AFB00014";
        ram_buffer(1981) := X"AFBF0034";
        ram_buffer(1982) := X"AFB70030";
        ram_buffer(1983) := X"AFB40024";
        ram_buffer(1984) := X"00008021";
        ram_buffer(1985) := X"00C0B021";
        ram_buffer(1986) := X"0080A821";
        ram_buffer(1987) := X"00A08821";
        ram_buffer(1988) := X"2413FFFF";
        ram_buffer(1989) := X"10000025";
        ram_buffer(1990) := X"2412002A";
        ram_buffer(1991) := X"8CA20000";
        ram_buffer(1992) := X"00000000";
        ram_buffer(1993) := X"24430001";
        ram_buffer(1994) := X"ACA30000";
        ram_buffer(1995) := X"90570000";
        ram_buffer(1996) := X"00000000";
        ram_buffer(1997) := X"A2970000";
        ram_buffer(1998) := X"8EA5000C";
        ram_buffer(1999) := X"8ED40004";
        ram_buffer(2000) := X"8CA20004";
        ram_buffer(2001) := X"0290A021";
        ram_buffer(2002) := X"2442FFFF";
        ram_buffer(2003) := X"04400033";
        ram_buffer(2004) := X"ACA20004";
        ram_buffer(2005) := X"8CA20000";
        ram_buffer(2006) := X"00000000";
        ram_buffer(2007) := X"24430001";
        ram_buffer(2008) := X"ACA30000";
        ram_buffer(2009) := X"90570000";
        ram_buffer(2010) := X"00000000";
        ram_buffer(2011) := X"A2970000";
        ram_buffer(2012) := X"8EA5000C";
        ram_buffer(2013) := X"8ED40008";
        ram_buffer(2014) := X"8CA20004";
        ram_buffer(2015) := X"0290A021";
        ram_buffer(2016) := X"2442FFFF";
        ram_buffer(2017) := X"0440003A";
        ram_buffer(2018) := X"ACA20004";
        ram_buffer(2019) := X"8CA20000";
        ram_buffer(2020) := X"00000000";
        ram_buffer(2021) := X"24430001";
        ram_buffer(2022) := X"ACA30000";
        ram_buffer(2023) := X"90570000";
        ram_buffer(2024) := X"26100001";
        ram_buffer(2025) := X"12300041";
        ram_buffer(2026) := X"A2970000";
        ram_buffer(2027) := X"8EA5000C";
        ram_buffer(2028) := X"8ED40000";
        ram_buffer(2029) := X"8CA20004";
        ram_buffer(2030) := X"0290A021";
        ram_buffer(2031) := X"2442FFFF";
        ram_buffer(2032) := X"0441FFD6";
        ram_buffer(2033) := X"ACA20004";
        ram_buffer(2034) := X"8F848098";
        ram_buffer(2035) := X"0C028350";
        ram_buffer(2036) := X"00000000";
        ram_buffer(2037) := X"1453FFD7";
        ram_buffer(2038) := X"0040B821";
        ram_buffer(2039) := X"8EA40018";
        ram_buffer(2040) := X"00000000";
        ram_buffer(2041) := X"8C820000";
        ram_buffer(2042) := X"00000000";
        ram_buffer(2043) := X"8C430000";
        ram_buffer(2044) := X"00000000";
        ram_buffer(2045) := X"0060F809";
        ram_buffer(2046) := X"AC520014";
        ram_buffer(2047) := X"A2970000";
        ram_buffer(2048) := X"8EA5000C";
        ram_buffer(2049) := X"8ED40004";
        ram_buffer(2050) := X"8CA20004";
        ram_buffer(2051) := X"0290A021";
        ram_buffer(2052) := X"2442FFFF";
        ram_buffer(2053) := X"0441FFCF";
        ram_buffer(2054) := X"ACA20004";
        ram_buffer(2055) := X"8F848098";
        ram_buffer(2056) := X"0C028350";
        ram_buffer(2057) := X"00000000";
        ram_buffer(2058) := X"1453FFD0";
        ram_buffer(2059) := X"0040B821";
        ram_buffer(2060) := X"8EA40018";
        ram_buffer(2061) := X"00000000";
        ram_buffer(2062) := X"8C820000";
        ram_buffer(2063) := X"00000000";
        ram_buffer(2064) := X"8C430000";
        ram_buffer(2065) := X"00000000";
        ram_buffer(2066) := X"0060F809";
        ram_buffer(2067) := X"AC520014";
        ram_buffer(2068) := X"A2970000";
        ram_buffer(2069) := X"8EA5000C";
        ram_buffer(2070) := X"8ED40008";
        ram_buffer(2071) := X"8CA20004";
        ram_buffer(2072) := X"0290A021";
        ram_buffer(2073) := X"2442FFFF";
        ram_buffer(2074) := X"0441FFC8";
        ram_buffer(2075) := X"ACA20004";
        ram_buffer(2076) := X"8F848098";
        ram_buffer(2077) := X"0C028350";
        ram_buffer(2078) := X"00000000";
        ram_buffer(2079) := X"1453FFC8";
        ram_buffer(2080) := X"0040B821";
        ram_buffer(2081) := X"8EA40018";
        ram_buffer(2082) := X"26100001";
        ram_buffer(2083) := X"8C820000";
        ram_buffer(2084) := X"00000000";
        ram_buffer(2085) := X"8C430000";
        ram_buffer(2086) := X"00000000";
        ram_buffer(2087) := X"0060F809";
        ram_buffer(2088) := X"AC520014";
        ram_buffer(2089) := X"1630FFC1";
        ram_buffer(2090) := X"A2970000";
        ram_buffer(2091) := X"8FBF0034";
        ram_buffer(2092) := X"8FB70030";
        ram_buffer(2093) := X"8FB6002C";
        ram_buffer(2094) := X"8FB50028";
        ram_buffer(2095) := X"8FB40024";
        ram_buffer(2096) := X"8FB30020";
        ram_buffer(2097) := X"8FB2001C";
        ram_buffer(2098) := X"8FB10018";
        ram_buffer(2099) := X"8FB00014";
        ram_buffer(2100) := X"27BD0038";
        ram_buffer(2101) := X"03E00008";
        ram_buffer(2102) := X"00000000";
        ram_buffer(2103) := X"8C82012C";
        ram_buffer(2104) := X"8C850140";
        ram_buffer(2105) := X"27BDFFD8";
        ram_buffer(2106) := X"8C830128";
        ram_buffer(2107) := X"AFB00010";
        ram_buffer(2108) := X"00808021";
        ram_buffer(2109) := X"00452021";
        ram_buffer(2110) := X"0064182A";
        ram_buffer(2111) := X"AFBF0024";
        ram_buffer(2112) := X"AFB40020";
        ram_buffer(2113) := X"AFB3001C";
        ram_buffer(2114) := X"AFB20018";
        ram_buffer(2115) := X"10600079";
        ram_buffer(2116) := X"AFB10014";
        ram_buffer(2117) := X"8E020130";
        ram_buffer(2118) := X"00000000";
        ram_buffer(2119) := X"14400037";
        ram_buffer(2120) := X"26120022";
        ram_buffer(2121) := X"8E110124";
        ram_buffer(2122) := X"2413002A";
        ram_buffer(2123) := X"2414FFFF";
        ram_buffer(2124) := X"02118821";
        ram_buffer(2125) := X"8222001E";
        ram_buffer(2126) := X"8E05000C";
        ram_buffer(2127) := X"A2020020";
        ram_buffer(2128) := X"8222001F";
        ram_buffer(2129) := X"00000000";
        ram_buffer(2130) := X"A2020021";
        ram_buffer(2131) := X"8CA20004";
        ram_buffer(2132) := X"00000000";
        ram_buffer(2133) := X"2442FFFF";
        ram_buffer(2134) := X"0440004D";
        ram_buffer(2135) := X"ACA20004";
        ram_buffer(2136) := X"8CA20000";
        ram_buffer(2137) := X"00000000";
        ram_buffer(2138) := X"24430001";
        ram_buffer(2139) := X"ACA30000";
        ram_buffer(2140) := X"90510000";
        ram_buffer(2141) := X"00000000";
        ram_buffer(2142) := X"1A200031";
        ram_buffer(2143) := X"02203021";
        ram_buffer(2144) := X"8E07000C";
        ram_buffer(2145) := X"24050001";
        ram_buffer(2146) := X"0C0272E9";
        ram_buffer(2147) := X"02402021";
        ram_buffer(2148) := X"12220009";
        ram_buffer(2149) := X"00000000";
        ram_buffer(2150) := X"8E040018";
        ram_buffer(2151) := X"00000000";
        ram_buffer(2152) := X"8C820000";
        ram_buffer(2153) := X"00000000";
        ram_buffer(2154) := X"8C430000";
        ram_buffer(2155) := X"00000000";
        ram_buffer(2156) := X"0060F809";
        ram_buffer(2157) := X"AC530014";
        ram_buffer(2158) := X"8E040128";
        ram_buffer(2159) := X"8E02012C";
        ram_buffer(2160) := X"8E050140";
        ram_buffer(2161) := X"00441023";
        ram_buffer(2162) := X"26310002";
        ram_buffer(2163) := X"24420010";
        ram_buffer(2164) := X"001118C0";
        ram_buffer(2165) := X"00A22021";
        ram_buffer(2166) := X"0064302A";
        ram_buffer(2167) := X"AE02012C";
        ram_buffer(2168) := X"AE110124";
        ram_buffer(2169) := X"10C00043";
        ram_buffer(2170) := X"AE030128";
        ram_buffer(2171) := X"8E020130";
        ram_buffer(2172) := X"00000000";
        ram_buffer(2173) := X"1040FFCF";
        ram_buffer(2174) := X"02118821";
        ram_buffer(2175) := X"8E040018";
        ram_buffer(2176) := X"24060400";
        ram_buffer(2177) := X"8C820000";
        ram_buffer(2178) := X"2405FFFF";
        ram_buffer(2179) := X"8C430004";
        ram_buffer(2180) := X"00000000";
        ram_buffer(2181) := X"0060F809";
        ram_buffer(2182) := X"AC460014";
        ram_buffer(2183) := X"8FBF0024";
        ram_buffer(2184) := X"8E02013C";
        ram_buffer(2185) := X"8FB40020";
        ram_buffer(2186) := X"8FB3001C";
        ram_buffer(2187) := X"8FB20018";
        ram_buffer(2188) := X"8FB10014";
        ram_buffer(2189) := X"8FB00010";
        ram_buffer(2190) := X"03E00008";
        ram_buffer(2191) := X"27BD0028";
        ram_buffer(2192) := X"1620FFDD";
        ram_buffer(2193) := X"24050001";
        ram_buffer(2194) := X"8E040018";
        ram_buffer(2195) := X"00000000";
        ram_buffer(2196) := X"8C820000";
        ram_buffer(2197) := X"24060400";
        ram_buffer(2198) := X"8C430004";
        ram_buffer(2199) := X"AE050130";
        ram_buffer(2200) := X"AC460014";
        ram_buffer(2201) := X"0060F809";
        ram_buffer(2202) := X"2405FFFF";
        ram_buffer(2203) := X"8FBF0024";
        ram_buffer(2204) := X"8E02013C";
        ram_buffer(2205) := X"8FB40020";
        ram_buffer(2206) := X"8FB3001C";
        ram_buffer(2207) := X"8FB20018";
        ram_buffer(2208) := X"8FB10014";
        ram_buffer(2209) := X"8FB00010";
        ram_buffer(2210) := X"03E00008";
        ram_buffer(2211) := X"27BD0028";
        ram_buffer(2212) := X"8F848098";
        ram_buffer(2213) := X"0C028350";
        ram_buffer(2214) := X"00000000";
        ram_buffer(2215) := X"1454FFB6";
        ram_buffer(2216) := X"00408821";
        ram_buffer(2217) := X"8E040018";
        ram_buffer(2218) := X"24110001";
        ram_buffer(2219) := X"8C820000";
        ram_buffer(2220) := X"00000000";
        ram_buffer(2221) := X"8C430000";
        ram_buffer(2222) := X"00000000";
        ram_buffer(2223) := X"0060F809";
        ram_buffer(2224) := X"AC530014";
        ram_buffer(2225) := X"8E040128";
        ram_buffer(2226) := X"8E02012C";
        ram_buffer(2227) := X"8E050140";
        ram_buffer(2228) := X"00441023";
        ram_buffer(2229) := X"24420010";
        ram_buffer(2230) := X"24030008";
        ram_buffer(2231) := X"00A22021";
        ram_buffer(2232) := X"0064302A";
        ram_buffer(2233) := X"AE02012C";
        ram_buffer(2234) := X"AE110124";
        ram_buffer(2235) := X"14C0FFBF";
        ram_buffer(2236) := X"AE030128";
        ram_buffer(2237) := X"000230C3";
        ram_buffer(2238) := X"02063021";
        ram_buffer(2239) := X"90C30022";
        ram_buffer(2240) := X"90C70021";
        ram_buffer(2241) := X"00031A00";
        ram_buffer(2242) := X"90C60020";
        ram_buffer(2243) := X"00E31825";
        ram_buffer(2244) := X"00031A00";
        ram_buffer(2245) := X"00C31825";
        ram_buffer(2246) := X"24060001";
        ram_buffer(2247) := X"8FBF0024";
        ram_buffer(2248) := X"30420007";
        ram_buffer(2249) := X"00A62804";
        ram_buffer(2250) := X"00431007";
        ram_buffer(2251) := X"24A5FFFF";
        ram_buffer(2252) := X"AE04012C";
        ram_buffer(2253) := X"8FB40020";
        ram_buffer(2254) := X"8FB3001C";
        ram_buffer(2255) := X"8FB20018";
        ram_buffer(2256) := X"8FB10014";
        ram_buffer(2257) := X"8FB00010";
        ram_buffer(2258) := X"00451024";
        ram_buffer(2259) := X"03E00008";
        ram_buffer(2260) := X"27BD0028";
        ram_buffer(2261) := X"8C830008";
        ram_buffer(2262) := X"8C82001C";
        ram_buffer(2263) := X"27BDFEB8";
        ram_buffer(2264) := X"AFBE0140";
        ram_buffer(2265) := X"AFBF0144";
        ram_buffer(2266) := X"AFB7013C";
        ram_buffer(2267) := X"AFB60138";
        ram_buffer(2268) := X"AFB50134";
        ram_buffer(2269) := X"AFB40130";
        ram_buffer(2270) := X"AFB3012C";
        ram_buffer(2271) := X"AFB20128";
        ram_buffer(2272) := X"AFB10124";
        ram_buffer(2273) := X"AFB00120";
        ram_buffer(2274) := X"AFA40148";
        ram_buffer(2275) := X"00A0F021";
        ram_buffer(2276) := X"104001C7";
        ram_buffer(2277) := X"AFA3011C";
        ram_buffer(2278) := X"AFA00118";
        ram_buffer(2279) := X"24150001";
        ram_buffer(2280) := X"24B00022";
        ram_buffer(2281) := X"8FA3011C";
        ram_buffer(2282) := X"00000000";
        ram_buffer(2283) := X"10600007";
        ram_buffer(2284) := X"00000000";
        ram_buffer(2285) := X"8FA40118";
        ram_buffer(2286) := X"8C650000";
        ram_buffer(2287) := X"AC640004";
        ram_buffer(2288) := X"8FA40148";
        ram_buffer(2289) := X"00A0F809";
        ram_buffer(2290) := X"AC620008";
        ram_buffer(2291) := X"8FA20148";
        ram_buffer(2292) := X"8FC5016C";
        ram_buffer(2293) := X"8C420004";
        ram_buffer(2294) := X"AFB50010";
        ram_buffer(2295) := X"8C42001C";
        ram_buffer(2296) := X"8FA60118";
        ram_buffer(2297) := X"8FA40148";
        ram_buffer(2298) := X"0040F809";
        ram_buffer(2299) := X"24070001";
        ram_buffer(2300) := X"8FA30148";
        ram_buffer(2301) := X"8C540000";
        ram_buffer(2302) := X"8C730018";
        ram_buffer(2303) := X"00000000";
        ram_buffer(2304) := X"1260007D";
        ram_buffer(2305) := X"2411002A";
        ram_buffer(2306) := X"8FC2014C";
        ram_buffer(2307) := X"00000000";
        ram_buffer(2308) := X"104000F0";
        ram_buffer(2309) := X"26940001";
        ram_buffer(2310) := X"8FC80138";
        ram_buffer(2311) := X"AFC0014C";
        ram_buffer(2312) := X"8FC20160";
        ram_buffer(2313) := X"8FC50134";
        ram_buffer(2314) := X"25040002";
        ram_buffer(2315) := X"AFC20164";
        ram_buffer(2316) := X"8FC2012C";
        ram_buffer(2317) := X"24A50001";
        ram_buffer(2318) := X"00083040";
        ram_buffer(2319) := X"AFC40148";
        ram_buffer(2320) := X"8FC40128";
        ram_buffer(2321) := X"AFC60144";
        ram_buffer(2322) := X"00453021";
        ram_buffer(2323) := X"0086202A";
        ram_buffer(2324) := X"AFC50140";
        ram_buffer(2325) := X"2412FFFF";
        ram_buffer(2326) := X"1080004E";
        ram_buffer(2327) := X"24160400";
        ram_buffer(2328) := X"8FC20130";
        ram_buffer(2329) := X"00000000";
        ram_buffer(2330) := X"14400036";
        ram_buffer(2331) := X"00000000";
        ram_buffer(2332) := X"8FC80124";
        ram_buffer(2333) := X"00000000";
        ram_buffer(2334) := X"03C84021";
        ram_buffer(2335) := X"8102001E";
        ram_buffer(2336) := X"8FC5000C";
        ram_buffer(2337) := X"A3C20020";
        ram_buffer(2338) := X"8102001F";
        ram_buffer(2339) := X"00000000";
        ram_buffer(2340) := X"A3C20021";
        ram_buffer(2341) := X"8CA20004";
        ram_buffer(2342) := X"00000000";
        ram_buffer(2343) := X"2442FFFF";
        ram_buffer(2344) := X"044000AF";
        ram_buffer(2345) := X"ACA20004";
        ram_buffer(2346) := X"8CA20000";
        ram_buffer(2347) := X"00000000";
        ram_buffer(2348) := X"24440001";
        ram_buffer(2349) := X"ACA40000";
        ram_buffer(2350) := X"90570000";
        ram_buffer(2351) := X"00000000";
        ram_buffer(2352) := X"1AE000A0";
        ram_buffer(2353) := X"02E03021";
        ram_buffer(2354) := X"8FC7000C";
        ram_buffer(2355) := X"24050001";
        ram_buffer(2356) := X"0C0272E9";
        ram_buffer(2357) := X"02002021";
        ram_buffer(2358) := X"12E20009";
        ram_buffer(2359) := X"00000000";
        ram_buffer(2360) := X"8FC40018";
        ram_buffer(2361) := X"00000000";
        ram_buffer(2362) := X"8C820000";
        ram_buffer(2363) := X"00000000";
        ram_buffer(2364) := X"8C450000";
        ram_buffer(2365) := X"00000000";
        ram_buffer(2366) := X"00A0F809";
        ram_buffer(2367) := X"AC510014";
        ram_buffer(2368) := X"8FC60128";
        ram_buffer(2369) := X"8FC2012C";
        ram_buffer(2370) := X"8FC50140";
        ram_buffer(2371) := X"00461023";
        ram_buffer(2372) := X"26E80002";
        ram_buffer(2373) := X"24420010";
        ram_buffer(2374) := X"000820C0";
        ram_buffer(2375) := X"00453021";
        ram_buffer(2376) := X"0086382A";
        ram_buffer(2377) := X"AFC2012C";
        ram_buffer(2378) := X"AFC80124";
        ram_buffer(2379) := X"10E000A6";
        ram_buffer(2380) := X"AFC40128";
        ram_buffer(2381) := X"8FC20130";
        ram_buffer(2382) := X"00000000";
        ram_buffer(2383) := X"1040FFCF";
        ram_buffer(2384) := X"03C84021";
        ram_buffer(2385) := X"8FC40018";
        ram_buffer(2386) := X"2405FFFF";
        ram_buffer(2387) := X"8C820000";
        ram_buffer(2388) := X"00000000";
        ram_buffer(2389) := X"8C460004";
        ram_buffer(2390) := X"00000000";
        ram_buffer(2391) := X"00C0F809";
        ram_buffer(2392) := X"AC560014";
        ram_buffer(2393) := X"8FC2013C";
        ram_buffer(2394) := X"8FC80138";
        ram_buffer(2395) := X"00000000";
        ram_buffer(2396) := X"15020018";
        ram_buffer(2397) := X"00000000";
        ram_buffer(2398) := X"8FC50140";
        ram_buffer(2399) := X"8FC2012C";
        ram_buffer(2400) := X"8FC40128";
        ram_buffer(2401) := X"00453021";
        ram_buffer(2402) := X"0086202A";
        ram_buffer(2403) := X"1480FFB4";
        ram_buffer(2404) := X"00000000";
        ram_buffer(2405) := X"000238C3";
        ram_buffer(2406) := X"03C73821";
        ram_buffer(2407) := X"90E40022";
        ram_buffer(2408) := X"90E90021";
        ram_buffer(2409) := X"00042200";
        ram_buffer(2410) := X"90E70020";
        ram_buffer(2411) := X"01242025";
        ram_buffer(2412) := X"00042200";
        ram_buffer(2413) := X"00E42025";
        ram_buffer(2414) := X"30420007";
        ram_buffer(2415) := X"00B52804";
        ram_buffer(2416) := X"00441007";
        ram_buffer(2417) := X"24A5FFFF";
        ram_buffer(2418) := X"00451024";
        ram_buffer(2419) := X"1102FFEA";
        ram_buffer(2420) := X"AFC6012C";
        ram_buffer(2421) := X"0102402A";
        ram_buffer(2422) := X"1500011E";
        ram_buffer(2423) := X"240303FD";
        ram_buffer(2424) := X"304400FF";
        ram_buffer(2425) := X"AFC20150";
        ram_buffer(2426) := X"AFC20154";
        ram_buffer(2427) := X"2673FFFF";
        ram_buffer(2428) := X"1660FF85";
        ram_buffer(2429) := X"A284FFFF";
        ram_buffer(2430) := X"8FA20148";
        ram_buffer(2431) := X"8FA30118";
        ram_buffer(2432) := X"8C42001C";
        ram_buffer(2433) := X"24630001";
        ram_buffer(2434) := X"0062202B";
        ram_buffer(2435) := X"1480FF65";
        ram_buffer(2436) := X"AFA30118";
        ram_buffer(2437) := X"24460007";
        ram_buffer(2438) := X"24440003";
        ram_buffer(2439) := X"000630C2";
        ram_buffer(2440) := X"24420001";
        ram_buffer(2441) := X"000420C2";
        ram_buffer(2442) := X"00862021";
        ram_buffer(2443) := X"00021082";
        ram_buffer(2444) := X"8FA3011C";
        ram_buffer(2445) := X"00441021";
        ram_buffer(2446) := X"10600005";
        ram_buffer(2447) := X"00000000";
        ram_buffer(2448) := X"8C650014";
        ram_buffer(2449) := X"00000000";
        ram_buffer(2450) := X"24A50001";
        ram_buffer(2451) := X"AC650014";
        ram_buffer(2452) := X"8FA30148";
        ram_buffer(2453) := X"8FC5016C";
        ram_buffer(2454) := X"8C670004";
        ram_buffer(2455) := X"AFA00010";
        ram_buffer(2456) := X"8CE8001C";
        ram_buffer(2457) := X"3C071008";
        ram_buffer(2458) := X"24E71D90";
        ram_buffer(2459) := X"AFC70004";
        ram_buffer(2460) := X"AFC60174";
        ram_buffer(2461) := X"AFC40178";
        ram_buffer(2462) := X"24070001";
        ram_buffer(2463) := X"00602021";
        ram_buffer(2464) := X"AFC00170";
        ram_buffer(2465) := X"AFC2017C";
        ram_buffer(2466) := X"8FD0001C";
        ram_buffer(2467) := X"0100F809";
        ram_buffer(2468) := X"00003021";
        ram_buffer(2469) := X"8FA30148";
        ram_buffer(2470) := X"8C440000";
        ram_buffer(2471) := X"8C650018";
        ram_buffer(2472) := X"8FC20010";
        ram_buffer(2473) := X"00000000";
        ram_buffer(2474) := X"8C420000";
        ram_buffer(2475) := X"10A00015";
        ram_buffer(2476) := X"00853821";
        ram_buffer(2477) := X"24840001";
        ram_buffer(2478) := X"9086FFFF";
        ram_buffer(2479) := X"8E050000";
        ram_buffer(2480) := X"24420003";
        ram_buffer(2481) := X"00A62821";
        ram_buffer(2482) := X"90A50000";
        ram_buffer(2483) := X"00000000";
        ram_buffer(2484) := X"A045FFFD";
        ram_buffer(2485) := X"8E050004";
        ram_buffer(2486) := X"00000000";
        ram_buffer(2487) := X"00A62821";
        ram_buffer(2488) := X"90A50000";
        ram_buffer(2489) := X"00000000";
        ram_buffer(2490) := X"A045FFFE";
        ram_buffer(2491) := X"8E050008";
        ram_buffer(2492) := X"00000000";
        ram_buffer(2493) := X"00A62821";
        ram_buffer(2494) := X"90A50000";
        ram_buffer(2495) := X"1487FFED";
        ram_buffer(2496) := X"A045FFFF";
        ram_buffer(2497) := X"8FC20170";
        ram_buffer(2498) := X"8FBF0144";
        ram_buffer(2499) := X"24420001";
        ram_buffer(2500) := X"AFC20170";
        ram_buffer(2501) := X"8FB7013C";
        ram_buffer(2502) := X"8FBE0140";
        ram_buffer(2503) := X"8FB60138";
        ram_buffer(2504) := X"8FB50134";
        ram_buffer(2505) := X"8FB40130";
        ram_buffer(2506) := X"8FB3012C";
        ram_buffer(2507) := X"8FB20128";
        ram_buffer(2508) := X"8FB10124";
        ram_buffer(2509) := X"8FB00120";
        ram_buffer(2510) := X"24020001";
        ram_buffer(2511) := X"03E00008";
        ram_buffer(2512) := X"27BD0148";
        ram_buffer(2513) := X"16E0FF6E";
        ram_buffer(2514) := X"2405FFFF";
        ram_buffer(2515) := X"8FC40018";
        ram_buffer(2516) := X"AFD50130";
        ram_buffer(2517) := X"8C820000";
        ram_buffer(2518) := X"1000FF7E";
        ram_buffer(2519) := X"00000000";
        ram_buffer(2520) := X"8F848098";
        ram_buffer(2521) := X"0C028350";
        ram_buffer(2522) := X"00000000";
        ram_buffer(2523) := X"1452FF54";
        ram_buffer(2524) := X"0040B821";
        ram_buffer(2525) := X"8FC40018";
        ram_buffer(2526) := X"00000000";
        ram_buffer(2527) := X"8C820000";
        ram_buffer(2528) := X"00000000";
        ram_buffer(2529) := X"8C450000";
        ram_buffer(2530) := X"00000000";
        ram_buffer(2531) := X"00A0F809";
        ram_buffer(2532) := X"AC510014";
        ram_buffer(2533) := X"8FC60128";
        ram_buffer(2534) := X"8FC2012C";
        ram_buffer(2535) := X"8FC50140";
        ram_buffer(2536) := X"00461023";
        ram_buffer(2537) := X"24420010";
        ram_buffer(2538) := X"24040008";
        ram_buffer(2539) := X"00453021";
        ram_buffer(2540) := X"24080001";
        ram_buffer(2541) := X"0086382A";
        ram_buffer(2542) := X"AFC2012C";
        ram_buffer(2543) := X"AFC80124";
        ram_buffer(2544) := X"14E0FF5C";
        ram_buffer(2545) := X"AFC40128";
        ram_buffer(2546) := X"8FC80138";
        ram_buffer(2547) := X"1000FF72";
        ram_buffer(2548) := X"000238C3";
        ram_buffer(2549) := X"8FC40164";
        ram_buffer(2550) := X"8FC20160";
        ram_buffer(2551) := X"00000000";
        ram_buffer(2552) := X"0044102B";
        ram_buffer(2553) := X"1040000F";
        ram_buffer(2554) := X"2482FFFF";
        ram_buffer(2555) := X"AFC20164";
        ram_buffer(2556) := X"9084FFFF";
        ram_buffer(2557) := X"2673FFFF";
        ram_buffer(2558) := X"1660FF03";
        ram_buffer(2559) := X"A284FFFF";
        ram_buffer(2560) := X"8FA20148";
        ram_buffer(2561) := X"8FA30118";
        ram_buffer(2562) := X"8C42001C";
        ram_buffer(2563) := X"24630001";
        ram_buffer(2564) := X"0062202B";
        ram_buffer(2565) := X"1480FEE3";
        ram_buffer(2566) := X"AFA30118";
        ram_buffer(2567) := X"1000FF7E";
        ram_buffer(2568) := X"24460007";
        ram_buffer(2569) := X"0C020837";
        ram_buffer(2570) := X"03C02021";
        ram_buffer(2571) := X"8FC40138";
        ram_buffer(2572) := X"00000000";
        ram_buffer(2573) := X"1044FEFA";
        ram_buffer(2574) := X"00804021";
        ram_buffer(2575) := X"8FC5013C";
        ram_buffer(2576) := X"00000000";
        ram_buffer(2577) := X"10450042";
        ram_buffer(2578) := X"00000000";
        ram_buffer(2579) := X"8FC50148";
        ram_buffer(2580) := X"00000000";
        ram_buffer(2581) := X"0045302A";
        ram_buffer(2582) := X"14C0001B";
        ram_buffer(2583) := X"00403821";
        ram_buffer(2584) := X"00A2282A";
        ram_buffer(2585) := X"14A00088";
        ram_buffer(2586) := X"240303FD";
        ram_buffer(2587) := X"8FC40164";
        ram_buffer(2588) := X"8FC50154";
        ram_buffer(2589) := X"24860001";
        ram_buffer(2590) := X"AFC60164";
        ram_buffer(2591) := X"A0850000";
        ram_buffer(2592) := X"00403821";
        ram_buffer(2593) := X"8FC40138";
        ram_buffer(2594) := X"8FC20150";
        ram_buffer(2595) := X"1000000F";
        ram_buffer(2596) := X"0044202A";
        ram_buffer(2597) := X"8FC50164";
        ram_buffer(2598) := X"8FC4015C";
        ram_buffer(2599) := X"24A60001";
        ram_buffer(2600) := X"AFC60164";
        ram_buffer(2601) := X"00822021";
        ram_buffer(2602) := X"90840000";
        ram_buffer(2603) := X"00021040";
        ram_buffer(2604) := X"A0A40000";
        ram_buffer(2605) := X"8FC50158";
        ram_buffer(2606) := X"8FC40138";
        ram_buffer(2607) := X"00A21021";
        ram_buffer(2608) := X"94420000";
        ram_buffer(2609) := X"00000000";
        ram_buffer(2610) := X"0044202A";
        ram_buffer(2611) := X"1080FFF1";
        ram_buffer(2612) := X"00000000";
        ram_buffer(2613) := X"8FC40148";
        ram_buffer(2614) := X"00000000";
        ram_buffer(2615) := X"28851000";
        ram_buffer(2616) := X"10A00018";
        ram_buffer(2617) := X"AFC20154";
        ram_buffer(2618) := X"8FC5015C";
        ram_buffer(2619) := X"8FC60158";
        ram_buffer(2620) := X"8FC80150";
        ram_buffer(2621) := X"00044840";
        ram_buffer(2622) := X"00C93021";
        ram_buffer(2623) := X"00A42021";
        ram_buffer(2624) := X"A4C80000";
        ram_buffer(2625) := X"A0820000";
        ram_buffer(2626) := X"8FC20148";
        ram_buffer(2627) := X"8FC40144";
        ram_buffer(2628) := X"24420001";
        ram_buffer(2629) := X"0044282A";
        ram_buffer(2630) := X"14A00009";
        ram_buffer(2631) := X"AFC20148";
        ram_buffer(2632) := X"8FC20140";
        ram_buffer(2633) := X"00000000";
        ram_buffer(2634) := X"2845000C";
        ram_buffer(2635) := X"10A00004";
        ram_buffer(2636) := X"24420001";
        ram_buffer(2637) := X"00042040";
        ram_buffer(2638) := X"AFC20140";
        ram_buffer(2639) := X"AFC40144";
        ram_buffer(2640) := X"8FC20154";
        ram_buffer(2641) := X"AFC70150";
        ram_buffer(2642) := X"1000FFAA";
        ram_buffer(2643) := X"304400FF";
        ram_buffer(2644) := X"8FC20130";
        ram_buffer(2645) := X"00000000";
        ram_buffer(2646) := X"14400034";
        ram_buffer(2647) := X"00000000";
        ram_buffer(2648) := X"2412FFFF";
        ram_buffer(2649) := X"8FC5000C";
        ram_buffer(2650) := X"00000000";
        ram_buffer(2651) := X"8CA20004";
        ram_buffer(2652) := X"00000000";
        ram_buffer(2653) := X"2442FFFF";
        ram_buffer(2654) := X"0440001E";
        ram_buffer(2655) := X"ACA20004";
        ram_buffer(2656) := X"8CA20000";
        ram_buffer(2657) := X"00000000";
        ram_buffer(2658) := X"24440001";
        ram_buffer(2659) := X"ACA40000";
        ram_buffer(2660) := X"90560000";
        ram_buffer(2661) := X"27A40018";
        ram_buffer(2662) := X"02C03021";
        ram_buffer(2663) := X"1AC00022";
        ram_buffer(2664) := X"24050001";
        ram_buffer(2665) := X"8FC7000C";
        ram_buffer(2666) := X"0C0272E9";
        ram_buffer(2667) := X"00000000";
        ram_buffer(2668) := X"12C2FFEC";
        ram_buffer(2669) := X"00000000";
        ram_buffer(2670) := X"8FC40018";
        ram_buffer(2671) := X"00000000";
        ram_buffer(2672) := X"8C820000";
        ram_buffer(2673) := X"00000000";
        ram_buffer(2674) := X"8C450000";
        ram_buffer(2675) := X"00000000";
        ram_buffer(2676) := X"00A0F809";
        ram_buffer(2677) := X"AC510014";
        ram_buffer(2678) := X"8FC5000C";
        ram_buffer(2679) := X"00000000";
        ram_buffer(2680) := X"8CA20004";
        ram_buffer(2681) := X"00000000";
        ram_buffer(2682) := X"2442FFFF";
        ram_buffer(2683) := X"0441FFE4";
        ram_buffer(2684) := X"ACA20004";
        ram_buffer(2685) := X"8F848098";
        ram_buffer(2686) := X"0C028350";
        ram_buffer(2687) := X"00000000";
        ram_buffer(2688) := X"1452FFE4";
        ram_buffer(2689) := X"0040B021";
        ram_buffer(2690) := X"8FC40018";
        ram_buffer(2691) := X"00000000";
        ram_buffer(2692) := X"8C820000";
        ram_buffer(2693) := X"00000000";
        ram_buffer(2694) := X"8C450000";
        ram_buffer(2695) := X"00000000";
        ram_buffer(2696) := X"00A0F809";
        ram_buffer(2697) := X"AC510014";
        ram_buffer(2698) := X"AFD50130";
        ram_buffer(2699) := X"8FC40018";
        ram_buffer(2700) := X"240303FF";
        ram_buffer(2701) := X"8C820000";
        ram_buffer(2702) := X"2405FFFF";
        ram_buffer(2703) := X"8C460004";
        ram_buffer(2704) := X"00000000";
        ram_buffer(2705) := X"00C0F809";
        ram_buffer(2706) := X"AC430014";
        ram_buffer(2707) := X"1000FF69";
        ram_buffer(2708) := X"00002021";
        ram_buffer(2709) := X"8FC40018";
        ram_buffer(2710) := X"00000000";
        ram_buffer(2711) := X"8C820000";
        ram_buffer(2712) := X"2405FFFF";
        ram_buffer(2713) := X"8C460004";
        ram_buffer(2714) := X"00000000";
        ram_buffer(2715) := X"00C0F809";
        ram_buffer(2716) := X"AC430014";
        ram_buffer(2717) := X"00001021";
        ram_buffer(2718) := X"00002021";
        ram_buffer(2719) := X"AFC20150";
        ram_buffer(2720) := X"1000FEDA";
        ram_buffer(2721) := X"AFC20154";
        ram_buffer(2722) := X"8FC40018";
        ram_buffer(2723) := X"00000000";
        ram_buffer(2724) := X"8C820000";
        ram_buffer(2725) := X"2405FFFF";
        ram_buffer(2726) := X"8C460004";
        ram_buffer(2727) := X"00000000";
        ram_buffer(2728) := X"00C0F809";
        ram_buffer(2729) := X"AC430014";
        ram_buffer(2730) := X"1000FF70";
        ram_buffer(2731) := X"00001021";
        ram_buffer(2732) := X"00002021";
        ram_buffer(2733) := X"1000FEE0";
        ram_buffer(2734) := X"00003021";
        ram_buffer(2735) := X"8C85000C";
        ram_buffer(2736) := X"27BDFED8";
        ram_buffer(2737) := X"8CA20004";
        ram_buffer(2738) := X"AFB10118";
        ram_buffer(2739) := X"2442FFFF";
        ram_buffer(2740) := X"AFBF0124";
        ram_buffer(2741) := X"AFB30120";
        ram_buffer(2742) := X"AFB2011C";
        ram_buffer(2743) := X"AFB00114";
        ram_buffer(2744) := X"00808821";
        ram_buffer(2745) := X"0440004B";
        ram_buffer(2746) := X"ACA20004";
        ram_buffer(2747) := X"8CA20000";
        ram_buffer(2748) := X"00000000";
        ram_buffer(2749) := X"24430001";
        ram_buffer(2750) := X"ACA30000";
        ram_buffer(2751) := X"90500000";
        ram_buffer(2752) := X"8E220018";
        ram_buffer(2753) := X"24050001";
        ram_buffer(2754) := X"8C430000";
        ram_buffer(2755) := X"240203FB";
        ram_buffer(2756) := X"AC700018";
        ram_buffer(2757) := X"8E240018";
        ram_buffer(2758) := X"AC620014";
        ram_buffer(2759) := X"8C820000";
        ram_buffer(2760) := X"2413FFFF";
        ram_buffer(2761) := X"8C420004";
        ram_buffer(2762) := X"00000000";
        ram_buffer(2763) := X"0040F809";
        ram_buffer(2764) := X"2412002A";
        ram_buffer(2765) := X"8E25000C";
        ram_buffer(2766) := X"00000000";
        ram_buffer(2767) := X"8CA20004";
        ram_buffer(2768) := X"00000000";
        ram_buffer(2769) := X"2442FFFF";
        ram_buffer(2770) := X"0440001E";
        ram_buffer(2771) := X"ACA20004";
        ram_buffer(2772) := X"8CA20000";
        ram_buffer(2773) := X"00000000";
        ram_buffer(2774) := X"24430001";
        ram_buffer(2775) := X"ACA30000";
        ram_buffer(2776) := X"90500000";
        ram_buffer(2777) := X"27A40010";
        ram_buffer(2778) := X"02003021";
        ram_buffer(2779) := X"1A000022";
        ram_buffer(2780) := X"24050001";
        ram_buffer(2781) := X"8E27000C";
        ram_buffer(2782) := X"0C0272E9";
        ram_buffer(2783) := X"00000000";
        ram_buffer(2784) := X"1202FFEC";
        ram_buffer(2785) := X"00000000";
        ram_buffer(2786) := X"8E240018";
        ram_buffer(2787) := X"00000000";
        ram_buffer(2788) := X"8C820000";
        ram_buffer(2789) := X"00000000";
        ram_buffer(2790) := X"8C430000";
        ram_buffer(2791) := X"00000000";
        ram_buffer(2792) := X"0060F809";
        ram_buffer(2793) := X"AC520014";
        ram_buffer(2794) := X"8E25000C";
        ram_buffer(2795) := X"00000000";
        ram_buffer(2796) := X"8CA20004";
        ram_buffer(2797) := X"00000000";
        ram_buffer(2798) := X"2442FFFF";
        ram_buffer(2799) := X"0441FFE4";
        ram_buffer(2800) := X"ACA20004";
        ram_buffer(2801) := X"8F848098";
        ram_buffer(2802) := X"0C028350";
        ram_buffer(2803) := X"00000000";
        ram_buffer(2804) := X"1453FFE4";
        ram_buffer(2805) := X"00408021";
        ram_buffer(2806) := X"8E240018";
        ram_buffer(2807) := X"2405002A";
        ram_buffer(2808) := X"8C820000";
        ram_buffer(2809) := X"00000000";
        ram_buffer(2810) := X"8C430000";
        ram_buffer(2811) := X"00000000";
        ram_buffer(2812) := X"0060F809";
        ram_buffer(2813) := X"AC450014";
        ram_buffer(2814) := X"8FBF0124";
        ram_buffer(2815) := X"8FB30120";
        ram_buffer(2816) := X"8FB2011C";
        ram_buffer(2817) := X"8FB10118";
        ram_buffer(2818) := X"8FB00114";
        ram_buffer(2819) := X"03E00008";
        ram_buffer(2820) := X"27BD0128";
        ram_buffer(2821) := X"8F848098";
        ram_buffer(2822) := X"0C028350";
        ram_buffer(2823) := X"00000000";
        ram_buffer(2824) := X"00408021";
        ram_buffer(2825) := X"2402FFFF";
        ram_buffer(2826) := X"1602FFB5";
        ram_buffer(2827) := X"2405002A";
        ram_buffer(2828) := X"8E240018";
        ram_buffer(2829) := X"00000000";
        ram_buffer(2830) := X"8C820000";
        ram_buffer(2831) := X"00000000";
        ram_buffer(2832) := X"8C430000";
        ram_buffer(2833) := X"00000000";
        ram_buffer(2834) := X"0060F809";
        ram_buffer(2835) := X"AC450014";
        ram_buffer(2836) := X"1000FFAB";
        ram_buffer(2837) := X"00000000";
        ram_buffer(2838) := X"8C820004";
        ram_buffer(2839) := X"27BDFFB0";
        ram_buffer(2840) := X"8C420008";
        ram_buffer(2841) := X"24070003";
        ram_buffer(2842) := X"AFBF004C";
        ram_buffer(2843) := X"AFB1002C";
        ram_buffer(2844) := X"AFB00028";
        ram_buffer(2845) := X"24060100";
        ram_buffer(2846) := X"00A08021";
        ram_buffer(2847) := X"AFBE0048";
        ram_buffer(2848) := X"24050001";
        ram_buffer(2849) := X"AFB70044";
        ram_buffer(2850) := X"AFB60040";
        ram_buffer(2851) := X"AFB5003C";
        ram_buffer(2852) := X"AFB40038";
        ram_buffer(2853) := X"AFB30034";
        ram_buffer(2854) := X"AFB20030";
        ram_buffer(2855) := X"0040F809";
        ram_buffer(2856) := X"00808821";
        ram_buffer(2857) := X"8E07000C";
        ram_buffer(2858) := X"AE02001C";
        ram_buffer(2859) := X"24060006";
        ram_buffer(2860) := X"24050001";
        ram_buffer(2861) := X"0C0272E9";
        ram_buffer(2862) := X"27A40018";
        ram_buffer(2863) := X"24030006";
        ram_buffer(2864) := X"10430007";
        ram_buffer(2865) := X"00000000";
        ram_buffer(2866) := X"8E220000";
        ram_buffer(2867) := X"240403F8";
        ram_buffer(2868) := X"8C430000";
        ram_buffer(2869) := X"AC440014";
        ram_buffer(2870) := X"0060F809";
        ram_buffer(2871) := X"02202021";
        ram_buffer(2872) := X"83A30018";
        ram_buffer(2873) := X"24020047";
        ram_buffer(2874) := X"106200FA";
        ram_buffer(2875) := X"24020049";
        ram_buffer(2876) := X"8E220000";
        ram_buffer(2877) := X"240403F8";
        ram_buffer(2878) := X"8C430000";
        ram_buffer(2879) := X"AC440014";
        ram_buffer(2880) := X"0060F809";
        ram_buffer(2881) := X"02202021";
        ram_buffer(2882) := X"83A3001B";
        ram_buffer(2883) := X"24020038";
        ram_buffer(2884) := X"83A4001C";
        ram_buffer(2885) := X"106200E5";
        ram_buffer(2886) := X"24020037";
        ram_buffer(2887) := X"83A5001D";
        ram_buffer(2888) := X"8E220000";
        ram_buffer(2889) := X"00000000";
        ram_buffer(2890) := X"AC430018";
        ram_buffer(2891) := X"8C460004";
        ram_buffer(2892) := X"240303FA";
        ram_buffer(2893) := X"AC44001C";
        ram_buffer(2894) := X"AC450020";
        ram_buffer(2895) := X"AC430014";
        ram_buffer(2896) := X"24050001";
        ram_buffer(2897) := X"00C0F809";
        ram_buffer(2898) := X"02202021";
        ram_buffer(2899) := X"8E07000C";
        ram_buffer(2900) := X"24060007";
        ram_buffer(2901) := X"24050001";
        ram_buffer(2902) := X"0C0272E9";
        ram_buffer(2903) := X"27A40018";
        ram_buffer(2904) := X"24030007";
        ram_buffer(2905) := X"10430007";
        ram_buffer(2906) := X"2404002A";
        ram_buffer(2907) := X"8E220000";
        ram_buffer(2908) := X"00000000";
        ram_buffer(2909) := X"8C430000";
        ram_buffer(2910) := X"AC440014";
        ram_buffer(2911) := X"0060F809";
        ram_buffer(2912) := X"02202021";
        ram_buffer(2913) := X"83A2001C";
        ram_buffer(2914) := X"93A3001E";
        ram_buffer(2915) := X"30440007";
        ram_buffer(2916) := X"24130002";
        ram_buffer(2917) := X"1060000C";
        ram_buffer(2918) := X"00939804";
        ram_buffer(2919) := X"24040031";
        ram_buffer(2920) := X"10640009";
        ram_buffer(2921) := X"24050001";
        ram_buffer(2922) := X"8E220000";
        ram_buffer(2923) := X"240403FC";
        ram_buffer(2924) := X"8C430004";
        ram_buffer(2925) := X"AC440014";
        ram_buffer(2926) := X"0060F809";
        ram_buffer(2927) := X"02202021";
        ram_buffer(2928) := X"83A2001C";
        ram_buffer(2929) := X"00000000";
        ram_buffer(2930) := X"04400119";
        ram_buffer(2931) := X"02602821";
        ram_buffer(2932) := X"241603FE";
        ram_buffer(2933) := X"2412003B";
        ram_buffer(2934) := X"24140021";
        ram_buffer(2935) := X"2415002C";
        ram_buffer(2936) := X"241703F7";
        ram_buffer(2937) := X"8E05000C";
        ram_buffer(2938) := X"00000000";
        ram_buffer(2939) := X"8CA20004";
        ram_buffer(2940) := X"00000000";
        ram_buffer(2941) := X"2442FFFF";
        ram_buffer(2942) := X"04400092";
        ram_buffer(2943) := X"ACA20004";
        ram_buffer(2944) := X"8CA20000";
        ram_buffer(2945) := X"00000000";
        ram_buffer(2946) := X"24430001";
        ram_buffer(2947) := X"ACA30000";
        ram_buffer(2948) := X"905E0000";
        ram_buffer(2949) := X"00000000";
        ram_buffer(2950) := X"13D200BC";
        ram_buffer(2951) := X"00000000";
        ram_buffer(2952) := X"13D400B6";
        ram_buffer(2953) := X"00000000";
        ram_buffer(2954) := X"17D50095";
        ram_buffer(2955) := X"24060009";
        ram_buffer(2956) := X"8E07000C";
        ram_buffer(2957) := X"24050001";
        ram_buffer(2958) := X"0C0272E9";
        ram_buffer(2959) := X"27A40018";
        ram_buffer(2960) := X"24030009";
        ram_buffer(2961) := X"10430007";
        ram_buffer(2962) := X"2404002A";
        ram_buffer(2963) := X"8E220000";
        ram_buffer(2964) := X"00000000";
        ram_buffer(2965) := X"8C430000";
        ram_buffer(2966) := X"AC440014";
        ram_buffer(2967) := X"0060F809";
        ram_buffer(2968) := X"02202021";
        ram_buffer(2969) := X"97A3001C";
        ram_buffer(2970) := X"97A2001E";
        ram_buffer(2971) := X"83A40020";
        ram_buffer(2972) := X"3072FFFF";
        ram_buffer(2973) := X"3054FFFF";
        ram_buffer(2974) := X"00031A00";
        ram_buffer(2975) := X"00021200";
        ram_buffer(2976) := X"00129202";
        ram_buffer(2977) := X"0014A202";
        ram_buffer(2978) := X"308500FF";
        ram_buffer(2979) := X"0054A025";
        ram_buffer(2980) := X"00729025";
        ram_buffer(2981) := X"30A20040";
        ram_buffer(2982) := X"3252FFFF";
        ram_buffer(2983) := X"3294FFFF";
        ram_buffer(2984) := X"048000DA";
        ram_buffer(2985) := X"AE020168";
        ram_buffer(2986) := X"8E05000C";
        ram_buffer(2987) := X"00000000";
        ram_buffer(2988) := X"8CA20004";
        ram_buffer(2989) := X"00000000";
        ram_buffer(2990) := X"2442FFFF";
        ram_buffer(2991) := X"044000B8";
        ram_buffer(2992) := X"ACA20004";
        ram_buffer(2993) := X"8CA20000";
        ram_buffer(2994) := X"00000000";
        ram_buffer(2995) := X"24430001";
        ram_buffer(2996) := X"ACA30000";
        ram_buffer(2997) := X"90550000";
        ram_buffer(2998) := X"00000000";
        ram_buffer(2999) := X"26A2FFFE";
        ram_buffer(3000) := X"2C42000A";
        ram_buffer(3001) := X"104000BE";
        ram_buffer(3002) := X"AE150134";
        ram_buffer(3003) := X"8E220004";
        ram_buffer(3004) := X"02202021";
        ram_buffer(3005) := X"8C420004";
        ram_buffer(3006) := X"24062000";
        ram_buffer(3007) := X"0040F809";
        ram_buffer(3008) := X"24050001";
        ram_buffer(3009) := X"8E230004";
        ram_buffer(3010) := X"02202021";
        ram_buffer(3011) := X"8C630004";
        ram_buffer(3012) := X"24061000";
        ram_buffer(3013) := X"24050001";
        ram_buffer(3014) := X"0060F809";
        ram_buffer(3015) := X"AE020158";
        ram_buffer(3016) := X"8E230004";
        ram_buffer(3017) := X"AE02015C";
        ram_buffer(3018) := X"8C620004";
        ram_buffer(3019) := X"24061000";
        ram_buffer(3020) := X"24050001";
        ram_buffer(3021) := X"0040F809";
        ram_buffer(3022) := X"02202021";
        ram_buffer(3023) := X"8E030134";
        ram_buffer(3024) := X"24050001";
        ram_buffer(3025) := X"00652004";
        ram_buffer(3026) := X"8E060168";
        ram_buffer(3027) := X"24890001";
        ram_buffer(3028) := X"24630001";
        ram_buffer(3029) := X"00044040";
        ram_buffer(3030) := X"24870002";
        ram_buffer(3031) := X"240A0002";
        ram_buffer(3032) := X"AE020160";
        ram_buffer(3033) := X"AE0A0124";
        ram_buffer(3034) := X"AE000128";
        ram_buffer(3035) := X"AE00012C";
        ram_buffer(3036) := X"AE000130";
        ram_buffer(3037) := X"AE040138";
        ram_buffer(3038) := X"AE09013C";
        ram_buffer(3039) := X"AE05014C";
        ram_buffer(3040) := X"AE030140";
        ram_buffer(3041) := X"AE080144";
        ram_buffer(3042) := X"AE070148";
        ram_buffer(3043) := X"14C00070";
        ram_buffer(3044) := X"AE020164";
        ram_buffer(3045) := X"3C021008";
        ram_buffer(3046) := X"24423244";
        ram_buffer(3047) := X"AE020004";
        ram_buffer(3048) := X"8E220004";
        ram_buffer(3049) := X"00123040";
        ram_buffer(3050) := X"8C420008";
        ram_buffer(3051) := X"02202021";
        ram_buffer(3052) := X"00D23021";
        ram_buffer(3053) := X"24050001";
        ram_buffer(3054) := X"0040F809";
        ram_buffer(3055) := X"24070001";
        ram_buffer(3056) := X"8E230000";
        ram_buffer(3057) := X"02202021";
        ram_buffer(3058) := X"8C660004";
        ram_buffer(3059) := X"AE020010";
        ram_buffer(3060) := X"24020001";
        ram_buffer(3061) := X"AE020014";
        ram_buffer(3062) := X"24020002";
        ram_buffer(3063) := X"AE220024";
        ram_buffer(3064) := X"24020003";
        ram_buffer(3065) := X"AE220020";
        ram_buffer(3066) := X"24020008";
        ram_buffer(3067) := X"AE220030";
        ram_buffer(3068) := X"240203F9";
        ram_buffer(3069) := X"AE320018";
        ram_buffer(3070) := X"AE34001C";
        ram_buffer(3071) := X"24050001";
        ram_buffer(3072) := X"AC720018";
        ram_buffer(3073) := X"AC74001C";
        ram_buffer(3074) := X"AC730020";
        ram_buffer(3075) := X"00C0F809";
        ram_buffer(3076) := X"AC620014";
        ram_buffer(3077) := X"8FBF004C";
        ram_buffer(3078) := X"8FBE0048";
        ram_buffer(3079) := X"8FB70044";
        ram_buffer(3080) := X"8FB60040";
        ram_buffer(3081) := X"8FB5003C";
        ram_buffer(3082) := X"8FB40038";
        ram_buffer(3083) := X"8FB30034";
        ram_buffer(3084) := X"8FB20030";
        ram_buffer(3085) := X"8FB1002C";
        ram_buffer(3086) := X"8FB00028";
        ram_buffer(3087) := X"03E00008";
        ram_buffer(3088) := X"27BD0050";
        ram_buffer(3089) := X"8F848098";
        ram_buffer(3090) := X"0C028350";
        ram_buffer(3091) := X"00000000";
        ram_buffer(3092) := X"0040F021";
        ram_buffer(3093) := X"2402FFFF";
        ram_buffer(3094) := X"17C2FF6F";
        ram_buffer(3095) := X"2405002A";
        ram_buffer(3096) := X"8E040018";
        ram_buffer(3097) := X"00000000";
        ram_buffer(3098) := X"8C820000";
        ram_buffer(3099) := X"00000000";
        ram_buffer(3100) := X"8C430000";
        ram_buffer(3101) := X"00000000";
        ram_buffer(3102) := X"0060F809";
        ram_buffer(3103) := X"AC450014";
        ram_buffer(3104) := X"8E220000";
        ram_buffer(3105) := X"2405FFFF";
        ram_buffer(3106) := X"AC5E0018";
        ram_buffer(3107) := X"8E230000";
        ram_buffer(3108) := X"AC560014";
        ram_buffer(3109) := X"8C620004";
        ram_buffer(3110) := X"00000000";
        ram_buffer(3111) := X"0040F809";
        ram_buffer(3112) := X"02202021";
        ram_buffer(3113) := X"1000FF4F";
        ram_buffer(3114) := X"00000000";
        ram_buffer(3115) := X"83A5001D";
        ram_buffer(3116) := X"10820003";
        ram_buffer(3117) := X"24020039";
        ram_buffer(3118) := X"1482FF19";
        ram_buffer(3119) := X"00000000";
        ram_buffer(3120) := X"24020061";
        ram_buffer(3121) := X"14A2FF16";
        ram_buffer(3122) := X"00000000";
        ram_buffer(3123) := X"1000FF1F";
        ram_buffer(3124) := X"00000000";
        ram_buffer(3125) := X"83A30019";
        ram_buffer(3126) := X"00000000";
        ram_buffer(3127) := X"1462FF04";
        ram_buffer(3128) := X"24020046";
        ram_buffer(3129) := X"83A3001A";
        ram_buffer(3130) := X"00000000";
        ram_buffer(3131) := X"1462FF00";
        ram_buffer(3132) := X"00000000";
        ram_buffer(3133) := X"1000FF04";
        ram_buffer(3134) := X"00000000";
        ram_buffer(3135) := X"0C020AAF";
        ram_buffer(3136) := X"02002021";
        ram_buffer(3137) := X"1000FF37";
        ram_buffer(3138) := X"00000000";
        ram_buffer(3139) := X"8E220000";
        ram_buffer(3140) := X"02202021";
        ram_buffer(3141) := X"8C430000";
        ram_buffer(3142) := X"00000000";
        ram_buffer(3143) := X"0060F809";
        ram_buffer(3144) := X"AC570014";
        ram_buffer(3145) := X"8E220000";
        ram_buffer(3146) := X"2405FFFF";
        ram_buffer(3147) := X"AC5E0018";
        ram_buffer(3148) := X"8E230000";
        ram_buffer(3149) := X"AC560014";
        ram_buffer(3150) := X"8C620004";
        ram_buffer(3151) := X"00000000";
        ram_buffer(3152) := X"0040F809";
        ram_buffer(3153) := X"02202021";
        ram_buffer(3154) := X"1000FF26";
        ram_buffer(3155) := X"00000000";
        ram_buffer(3156) := X"8E220004";
        ram_buffer(3157) := X"AFA50014";
        ram_buffer(3158) := X"AFB40010";
        ram_buffer(3159) := X"8C420010";
        ram_buffer(3160) := X"02403821";
        ram_buffer(3161) := X"00003021";
        ram_buffer(3162) := X"0040F809";
        ram_buffer(3163) := X"02202021";
        ram_buffer(3164) := X"8E230008";
        ram_buffer(3165) := X"00000000";
        ram_buffer(3166) := X"10600005";
        ram_buffer(3167) := X"AE02016C";
        ram_buffer(3168) := X"8C620018";
        ram_buffer(3169) := X"00000000";
        ram_buffer(3170) := X"24420001";
        ram_buffer(3171) := X"AC620018";
        ram_buffer(3172) := X"3C021008";
        ram_buffer(3173) := X"24422354";
        ram_buffer(3174) := X"1000FF81";
        ram_buffer(3175) := X"AE020004";
        ram_buffer(3176) := X"8F848098";
        ram_buffer(3177) := X"0C028350";
        ram_buffer(3178) := X"00000000";
        ram_buffer(3179) := X"0040A821";
        ram_buffer(3180) := X"2402FFFF";
        ram_buffer(3181) := X"16A2FF49";
        ram_buffer(3182) := X"2405002A";
        ram_buffer(3183) := X"8E040018";
        ram_buffer(3184) := X"00000000";
        ram_buffer(3185) := X"8C820000";
        ram_buffer(3186) := X"00000000";
        ram_buffer(3187) := X"8C430000";
        ram_buffer(3188) := X"00000000";
        ram_buffer(3189) := X"0060F809";
        ram_buffer(3190) := X"AC450014";
        ram_buffer(3191) := X"AE150134";
        ram_buffer(3192) := X"8E220000";
        ram_buffer(3193) := X"240403F5";
        ram_buffer(3194) := X"AC550018";
        ram_buffer(3195) := X"8E230000";
        ram_buffer(3196) := X"AC440014";
        ram_buffer(3197) := X"8C620000";
        ram_buffer(3198) := X"00000000";
        ram_buffer(3199) := X"0040F809";
        ram_buffer(3200) := X"02202021";
        ram_buffer(3201) := X"1000FF39";
        ram_buffer(3202) := X"00000000";
        ram_buffer(3203) := X"30A50007";
        ram_buffer(3204) := X"24130002";
        ram_buffer(3205) := X"00B39804";
        ram_buffer(3206) := X"8E06001C";
        ram_buffer(3207) := X"02602821";
        ram_buffer(3208) := X"0C0207B4";
        ram_buffer(3209) := X"02002021";
        ram_buffer(3210) := X"1000FF1F";
        ram_buffer(3211) := X"00000000";
        ram_buffer(3212) := X"8E06001C";
        ram_buffer(3213) := X"0C0207B4";
        ram_buffer(3214) := X"02002021";
        ram_buffer(3215) := X"1000FEE5";
        ram_buffer(3216) := X"241603FE";
        ram_buffer(3217) := X"27BDFEC8";
        ram_buffer(3218) := X"8CA20010";
        ram_buffer(3219) := X"AFB40120";
        ram_buffer(3220) := X"8C940018";
        ram_buffer(3221) := X"AFB50124";
        ram_buffer(3222) := X"AFB20118";
        ram_buffer(3223) := X"AFBF0134";
        ram_buffer(3224) := X"AFBE0130";
        ram_buffer(3225) := X"AFB7012C";
        ram_buffer(3226) := X"AFB60128";
        ram_buffer(3227) := X"AFB3011C";
        ram_buffer(3228) := X"AFB10114";
        ram_buffer(3229) := X"AFB00110";
        ram_buffer(3230) := X"8CB5001C";
        ram_buffer(3231) := X"8C520000";
        ram_buffer(3232) := X"128000BB";
        ram_buffer(3233) := X"00A0F021";
        ram_buffer(3234) := X"2411002A";
        ram_buffer(3235) := X"24B00022";
        ram_buffer(3236) := X"8FC2014C";
        ram_buffer(3237) := X"00000000";
        ram_buffer(3238) := X"1040009B";
        ram_buffer(3239) := X"00000000";
        ram_buffer(3240) := X"8FC80138";
        ram_buffer(3241) := X"AFC0014C";
        ram_buffer(3242) := X"8FC20160";
        ram_buffer(3243) := X"8FC50134";
        ram_buffer(3244) := X"25040002";
        ram_buffer(3245) := X"AFC20164";
        ram_buffer(3246) := X"8FC2012C";
        ram_buffer(3247) := X"24A50001";
        ram_buffer(3248) := X"00083040";
        ram_buffer(3249) := X"AFC40148";
        ram_buffer(3250) := X"8FC40128";
        ram_buffer(3251) := X"AFC60144";
        ram_buffer(3252) := X"00453021";
        ram_buffer(3253) := X"0086202A";
        ram_buffer(3254) := X"AFC50140";
        ram_buffer(3255) := X"24160001";
        ram_buffer(3256) := X"1080004E";
        ram_buffer(3257) := X"2413FFFF";
        ram_buffer(3258) := X"8FC20130";
        ram_buffer(3259) := X"00000000";
        ram_buffer(3260) := X"14400036";
        ram_buffer(3261) := X"00000000";
        ram_buffer(3262) := X"8FC80124";
        ram_buffer(3263) := X"00000000";
        ram_buffer(3264) := X"03C84021";
        ram_buffer(3265) := X"8102001E";
        ram_buffer(3266) := X"8FC5000C";
        ram_buffer(3267) := X"A3C20020";
        ram_buffer(3268) := X"8102001F";
        ram_buffer(3269) := X"00000000";
        ram_buffer(3270) := X"A3C20021";
        ram_buffer(3271) := X"8CA20004";
        ram_buffer(3272) := X"00000000";
        ram_buffer(3273) := X"2442FFFF";
        ram_buffer(3274) := X"0440005A";
        ram_buffer(3275) := X"ACA20004";
        ram_buffer(3276) := X"8CA20000";
        ram_buffer(3277) := X"00000000";
        ram_buffer(3278) := X"24440001";
        ram_buffer(3279) := X"ACA40000";
        ram_buffer(3280) := X"90570000";
        ram_buffer(3281) := X"00000000";
        ram_buffer(3282) := X"1AE0004B";
        ram_buffer(3283) := X"02E03021";
        ram_buffer(3284) := X"8FC7000C";
        ram_buffer(3285) := X"24050001";
        ram_buffer(3286) := X"0C0272E9";
        ram_buffer(3287) := X"02002021";
        ram_buffer(3288) := X"12E20009";
        ram_buffer(3289) := X"00000000";
        ram_buffer(3290) := X"8FC40018";
        ram_buffer(3291) := X"00000000";
        ram_buffer(3292) := X"8C820000";
        ram_buffer(3293) := X"00000000";
        ram_buffer(3294) := X"8C450000";
        ram_buffer(3295) := X"00000000";
        ram_buffer(3296) := X"00A0F809";
        ram_buffer(3297) := X"AC510014";
        ram_buffer(3298) := X"8FC60128";
        ram_buffer(3299) := X"8FC2012C";
        ram_buffer(3300) := X"8FC50140";
        ram_buffer(3301) := X"00461023";
        ram_buffer(3302) := X"26E80002";
        ram_buffer(3303) := X"24420010";
        ram_buffer(3304) := X"000820C0";
        ram_buffer(3305) := X"00453021";
        ram_buffer(3306) := X"0086382A";
        ram_buffer(3307) := X"AFC2012C";
        ram_buffer(3308) := X"AFC80124";
        ram_buffer(3309) := X"10E00051";
        ram_buffer(3310) := X"AFC40128";
        ram_buffer(3311) := X"8FC20130";
        ram_buffer(3312) := X"00000000";
        ram_buffer(3313) := X"1040FFCF";
        ram_buffer(3314) := X"03C84021";
        ram_buffer(3315) := X"8FC40018";
        ram_buffer(3316) := X"2405FFFF";
        ram_buffer(3317) := X"8C820000";
        ram_buffer(3318) := X"24030400";
        ram_buffer(3319) := X"8C460004";
        ram_buffer(3320) := X"00000000";
        ram_buffer(3321) := X"00C0F809";
        ram_buffer(3322) := X"AC430014";
        ram_buffer(3323) := X"8FC4013C";
        ram_buffer(3324) := X"8FC80138";
        ram_buffer(3325) := X"00000000";
        ram_buffer(3326) := X"15040018";
        ram_buffer(3327) := X"00000000";
        ram_buffer(3328) := X"8FC50140";
        ram_buffer(3329) := X"8FC2012C";
        ram_buffer(3330) := X"8FC40128";
        ram_buffer(3331) := X"00453021";
        ram_buffer(3332) := X"0086202A";
        ram_buffer(3333) := X"1480FFB4";
        ram_buffer(3334) := X"00000000";
        ram_buffer(3335) := X"000238C3";
        ram_buffer(3336) := X"03C73821";
        ram_buffer(3337) := X"90E40022";
        ram_buffer(3338) := X"90E90021";
        ram_buffer(3339) := X"00042200";
        ram_buffer(3340) := X"90E70020";
        ram_buffer(3341) := X"01242025";
        ram_buffer(3342) := X"00042200";
        ram_buffer(3343) := X"00E42025";
        ram_buffer(3344) := X"30420007";
        ram_buffer(3345) := X"00B62804";
        ram_buffer(3346) := X"00441007";
        ram_buffer(3347) := X"24A4FFFF";
        ram_buffer(3348) := X"00442024";
        ram_buffer(3349) := X"1104FFEA";
        ram_buffer(3350) := X"AFC6012C";
        ram_buffer(3351) := X"0104402A";
        ram_buffer(3352) := X"150000DC";
        ram_buffer(3353) := X"240303FD";
        ram_buffer(3354) := X"00801021";
        ram_buffer(3355) := X"AFC40150";
        ram_buffer(3356) := X"1000002D";
        ram_buffer(3357) := X"AFC40154";
        ram_buffer(3358) := X"16E0FFC3";
        ram_buffer(3359) := X"2405FFFF";
        ram_buffer(3360) := X"8FC40018";
        ram_buffer(3361) := X"AFD60130";
        ram_buffer(3362) := X"8C820000";
        ram_buffer(3363) := X"1000FFD3";
        ram_buffer(3364) := X"24030400";
        ram_buffer(3365) := X"8F848098";
        ram_buffer(3366) := X"0C028350";
        ram_buffer(3367) := X"00000000";
        ram_buffer(3368) := X"1453FFA9";
        ram_buffer(3369) := X"0040B821";
        ram_buffer(3370) := X"8FC40018";
        ram_buffer(3371) := X"00000000";
        ram_buffer(3372) := X"8C820000";
        ram_buffer(3373) := X"00000000";
        ram_buffer(3374) := X"8C450000";
        ram_buffer(3375) := X"00000000";
        ram_buffer(3376) := X"00A0F809";
        ram_buffer(3377) := X"AC510014";
        ram_buffer(3378) := X"8FC60128";
        ram_buffer(3379) := X"8FC2012C";
        ram_buffer(3380) := X"8FC50140";
        ram_buffer(3381) := X"00461023";
        ram_buffer(3382) := X"24420010";
        ram_buffer(3383) := X"24040008";
        ram_buffer(3384) := X"00453021";
        ram_buffer(3385) := X"24080001";
        ram_buffer(3386) := X"0086382A";
        ram_buffer(3387) := X"AFC2012C";
        ram_buffer(3388) := X"AFC80124";
        ram_buffer(3389) := X"14E0FFB1";
        ram_buffer(3390) := X"AFC40128";
        ram_buffer(3391) := X"8FC80138";
        ram_buffer(3392) := X"1000FFC7";
        ram_buffer(3393) := X"000238C3";
        ram_buffer(3394) := X"8FC40164";
        ram_buffer(3395) := X"8FC20160";
        ram_buffer(3396) := X"00000000";
        ram_buffer(3397) := X"0044102B";
        ram_buffer(3398) := X"10400022";
        ram_buffer(3399) := X"2482FFFF";
        ram_buffer(3400) := X"AFC20164";
        ram_buffer(3401) := X"9082FFFF";
        ram_buffer(3402) := X"8EA40000";
        ram_buffer(3403) := X"26520003";
        ram_buffer(3404) := X"00822021";
        ram_buffer(3405) := X"90840000";
        ram_buffer(3406) := X"2694FFFF";
        ram_buffer(3407) := X"A244FFFD";
        ram_buffer(3408) := X"8EA40004";
        ram_buffer(3409) := X"00000000";
        ram_buffer(3410) := X"00822021";
        ram_buffer(3411) := X"90840000";
        ram_buffer(3412) := X"00000000";
        ram_buffer(3413) := X"A244FFFE";
        ram_buffer(3414) := X"8EA40008";
        ram_buffer(3415) := X"00000000";
        ram_buffer(3416) := X"00821021";
        ram_buffer(3417) := X"90420000";
        ram_buffer(3418) := X"1680FF49";
        ram_buffer(3419) := X"A242FFFF";
        ram_buffer(3420) := X"8FBF0134";
        ram_buffer(3421) := X"8FBE0130";
        ram_buffer(3422) := X"8FB7012C";
        ram_buffer(3423) := X"8FB60128";
        ram_buffer(3424) := X"8FB50124";
        ram_buffer(3425) := X"8FB40120";
        ram_buffer(3426) := X"8FB3011C";
        ram_buffer(3427) := X"8FB20118";
        ram_buffer(3428) := X"8FB10114";
        ram_buffer(3429) := X"8FB00110";
        ram_buffer(3430) := X"24020001";
        ram_buffer(3431) := X"03E00008";
        ram_buffer(3432) := X"27BD0138";
        ram_buffer(3433) := X"0C020837";
        ram_buffer(3434) := X"03C02021";
        ram_buffer(3435) := X"8FC40138";
        ram_buffer(3436) := X"00000000";
        ram_buffer(3437) := X"1044FF3C";
        ram_buffer(3438) := X"00804021";
        ram_buffer(3439) := X"8FC5013C";
        ram_buffer(3440) := X"00000000";
        ram_buffer(3441) := X"10450041";
        ram_buffer(3442) := X"00000000";
        ram_buffer(3443) := X"8FC50148";
        ram_buffer(3444) := X"00000000";
        ram_buffer(3445) := X"0045302A";
        ram_buffer(3446) := X"14C0001B";
        ram_buffer(3447) := X"00403821";
        ram_buffer(3448) := X"00A2282A";
        ram_buffer(3449) := X"14A00088";
        ram_buffer(3450) := X"240303FD";
        ram_buffer(3451) := X"8FC40164";
        ram_buffer(3452) := X"8FC50154";
        ram_buffer(3453) := X"24860001";
        ram_buffer(3454) := X"AFC60164";
        ram_buffer(3455) := X"A0850000";
        ram_buffer(3456) := X"00403821";
        ram_buffer(3457) := X"8FC40138";
        ram_buffer(3458) := X"8FC20150";
        ram_buffer(3459) := X"1000000F";
        ram_buffer(3460) := X"0044202A";
        ram_buffer(3461) := X"8FC50164";
        ram_buffer(3462) := X"8FC4015C";
        ram_buffer(3463) := X"24A60001";
        ram_buffer(3464) := X"AFC60164";
        ram_buffer(3465) := X"00822021";
        ram_buffer(3466) := X"90840000";
        ram_buffer(3467) := X"00021040";
        ram_buffer(3468) := X"A0A40000";
        ram_buffer(3469) := X"8FC50158";
        ram_buffer(3470) := X"8FC40138";
        ram_buffer(3471) := X"00A21021";
        ram_buffer(3472) := X"94420000";
        ram_buffer(3473) := X"00000000";
        ram_buffer(3474) := X"0044202A";
        ram_buffer(3475) := X"1080FFF1";
        ram_buffer(3476) := X"00000000";
        ram_buffer(3477) := X"8FC40148";
        ram_buffer(3478) := X"00000000";
        ram_buffer(3479) := X"28851000";
        ram_buffer(3480) := X"10A00018";
        ram_buffer(3481) := X"AFC20154";
        ram_buffer(3482) := X"8FC5015C";
        ram_buffer(3483) := X"8FC60158";
        ram_buffer(3484) := X"8FC80150";
        ram_buffer(3485) := X"00044840";
        ram_buffer(3486) := X"00C93021";
        ram_buffer(3487) := X"00A42021";
        ram_buffer(3488) := X"A4C80000";
        ram_buffer(3489) := X"A0820000";
        ram_buffer(3490) := X"8FC20148";
        ram_buffer(3491) := X"8FC40144";
        ram_buffer(3492) := X"24420001";
        ram_buffer(3493) := X"0044282A";
        ram_buffer(3494) := X"14A00009";
        ram_buffer(3495) := X"AFC20148";
        ram_buffer(3496) := X"8FC20140";
        ram_buffer(3497) := X"00000000";
        ram_buffer(3498) := X"2845000C";
        ram_buffer(3499) := X"10A00004";
        ram_buffer(3500) := X"00042040";
        ram_buffer(3501) := X"24420001";
        ram_buffer(3502) := X"AFC20140";
        ram_buffer(3503) := X"AFC40144";
        ram_buffer(3504) := X"8FC20154";
        ram_buffer(3505) := X"1000FF98";
        ram_buffer(3506) := X"AFC70150";
        ram_buffer(3507) := X"8FC20130";
        ram_buffer(3508) := X"00000000";
        ram_buffer(3509) := X"14400035";
        ram_buffer(3510) := X"00000000";
        ram_buffer(3511) := X"2413FFFF";
        ram_buffer(3512) := X"8FC5000C";
        ram_buffer(3513) := X"00000000";
        ram_buffer(3514) := X"8CA20004";
        ram_buffer(3515) := X"00000000";
        ram_buffer(3516) := X"2442FFFF";
        ram_buffer(3517) := X"0440001E";
        ram_buffer(3518) := X"ACA20004";
        ram_buffer(3519) := X"8CA20000";
        ram_buffer(3520) := X"00000000";
        ram_buffer(3521) := X"24440001";
        ram_buffer(3522) := X"ACA40000";
        ram_buffer(3523) := X"90560000";
        ram_buffer(3524) := X"27A40010";
        ram_buffer(3525) := X"02C03021";
        ram_buffer(3526) := X"1AC00022";
        ram_buffer(3527) := X"24050001";
        ram_buffer(3528) := X"8FC7000C";
        ram_buffer(3529) := X"0C0272E9";
        ram_buffer(3530) := X"00000000";
        ram_buffer(3531) := X"12C2FFEC";
        ram_buffer(3532) := X"00000000";
        ram_buffer(3533) := X"8FC40018";
        ram_buffer(3534) := X"00000000";
        ram_buffer(3535) := X"8C820000";
        ram_buffer(3536) := X"00000000";
        ram_buffer(3537) := X"8C450000";
        ram_buffer(3538) := X"00000000";
        ram_buffer(3539) := X"00A0F809";
        ram_buffer(3540) := X"AC510014";
        ram_buffer(3541) := X"8FC5000C";
        ram_buffer(3542) := X"00000000";
        ram_buffer(3543) := X"8CA20004";
        ram_buffer(3544) := X"00000000";
        ram_buffer(3545) := X"2442FFFF";
        ram_buffer(3546) := X"0441FFE4";
        ram_buffer(3547) := X"ACA20004";
        ram_buffer(3548) := X"8F848098";
        ram_buffer(3549) := X"0C028350";
        ram_buffer(3550) := X"00000000";
        ram_buffer(3551) := X"1453FFE4";
        ram_buffer(3552) := X"0040B021";
        ram_buffer(3553) := X"8FC40018";
        ram_buffer(3554) := X"00000000";
        ram_buffer(3555) := X"8C820000";
        ram_buffer(3556) := X"00000000";
        ram_buffer(3557) := X"8C450000";
        ram_buffer(3558) := X"00000000";
        ram_buffer(3559) := X"00A0F809";
        ram_buffer(3560) := X"AC510014";
        ram_buffer(3561) := X"24020001";
        ram_buffer(3562) := X"AFC20130";
        ram_buffer(3563) := X"8FC40018";
        ram_buffer(3564) := X"240303FF";
        ram_buffer(3565) := X"8C820000";
        ram_buffer(3566) := X"2405FFFF";
        ram_buffer(3567) := X"8C460004";
        ram_buffer(3568) := X"00000000";
        ram_buffer(3569) := X"00C0F809";
        ram_buffer(3570) := X"AC430014";
        ram_buffer(3571) := X"1000FF56";
        ram_buffer(3572) := X"00001021";
        ram_buffer(3573) := X"8FC40018";
        ram_buffer(3574) := X"00000000";
        ram_buffer(3575) := X"8C820000";
        ram_buffer(3576) := X"2405FFFF";
        ram_buffer(3577) := X"8C460004";
        ram_buffer(3578) := X"00000000";
        ram_buffer(3579) := X"00C0F809";
        ram_buffer(3580) := X"AC430014";
        ram_buffer(3581) := X"00002021";
        ram_buffer(3582) := X"00001021";
        ram_buffer(3583) := X"AFC40150";
        ram_buffer(3584) := X"1000FF49";
        ram_buffer(3585) := X"AFC40154";
        ram_buffer(3586) := X"8FC40018";
        ram_buffer(3587) := X"00000000";
        ram_buffer(3588) := X"8C820000";
        ram_buffer(3589) := X"2405FFFF";
        ram_buffer(3590) := X"8C460004";
        ram_buffer(3591) := X"00000000";
        ram_buffer(3592) := X"00C0F809";
        ram_buffer(3593) := X"AC430014";
        ram_buffer(3594) := X"1000FF70";
        ram_buffer(3595) := X"00001021";
        ram_buffer(3596) := X"8C820004";
        ram_buffer(3597) := X"27BDFFE8";
        ram_buffer(3598) := X"8C420000";
        ram_buffer(3599) := X"24060180";
        ram_buffer(3600) := X"AFBF0014";
        ram_buffer(3601) := X"AFB00010";
        ram_buffer(3602) := X"24050001";
        ram_buffer(3603) := X"0040F809";
        ram_buffer(3604) := X"00808021";
        ram_buffer(3605) := X"3C041008";
        ram_buffer(3606) := X"24842C58";
        ram_buffer(3607) := X"AC440000";
        ram_buffer(3608) := X"8FBF0014";
        ram_buffer(3609) := X"3C041008";
        ram_buffer(3610) := X"24841EC8";
        ram_buffer(3611) := X"AC500018";
        ram_buffer(3612) := X"AC440008";
        ram_buffer(3613) := X"8FB00010";
        ram_buffer(3614) := X"03E00008";
        ram_buffer(3615) := X"27BD0018";
        ram_buffer(3616) := X"27BDFFE0";
        ram_buffer(3617) := X"8CA20010";
        ram_buffer(3618) := X"AFB00010";
        ram_buffer(3619) := X"8C900018";
        ram_buffer(3620) := X"AFB20018";
        ram_buffer(3621) := X"AFBF001C";
        ram_buffer(3622) := X"AFB10014";
        ram_buffer(3623) := X"8C520000";
        ram_buffer(3624) := X"1200000A";
        ram_buffer(3625) := X"00A08821";
        ram_buffer(3626) := X"8E220028";
        ram_buffer(3627) := X"00000000";
        ram_buffer(3628) := X"0040F809";
        ram_buffer(3629) := X"02202021";
        ram_buffer(3630) := X"9222002C";
        ram_buffer(3631) := X"26520001";
        ram_buffer(3632) := X"2610FFFF";
        ram_buffer(3633) := X"1600FFF8";
        ram_buffer(3634) := X"A242FFFF";
        ram_buffer(3635) := X"8FBF001C";
        ram_buffer(3636) := X"8FB20018";
        ram_buffer(3637) := X"8FB10014";
        ram_buffer(3638) := X"8FB00010";
        ram_buffer(3639) := X"24020001";
        ram_buffer(3640) := X"03E00008";
        ram_buffer(3641) := X"27BD0020";
        ram_buffer(3642) := X"27BDFFD8";
        ram_buffer(3643) := X"8CA20010";
        ram_buffer(3644) := X"AFB2001C";
        ram_buffer(3645) := X"8C920018";
        ram_buffer(3646) := X"AFB30020";
        ram_buffer(3647) := X"AFB00014";
        ram_buffer(3648) := X"AFBF0024";
        ram_buffer(3649) := X"AFB10018";
        ram_buffer(3650) := X"8CB3001C";
        ram_buffer(3651) := X"8C500000";
        ram_buffer(3652) := X"12400018";
        ram_buffer(3653) := X"00A08821";
        ram_buffer(3654) := X"8E220028";
        ram_buffer(3655) := X"00000000";
        ram_buffer(3656) := X"0040F809";
        ram_buffer(3657) := X"02202021";
        ram_buffer(3658) := X"9223002C";
        ram_buffer(3659) := X"8E620000";
        ram_buffer(3660) := X"26100003";
        ram_buffer(3661) := X"00431021";
        ram_buffer(3662) := X"90420000";
        ram_buffer(3663) := X"2652FFFF";
        ram_buffer(3664) := X"A202FFFD";
        ram_buffer(3665) := X"8E620004";
        ram_buffer(3666) := X"00000000";
        ram_buffer(3667) := X"00431021";
        ram_buffer(3668) := X"90420000";
        ram_buffer(3669) := X"00000000";
        ram_buffer(3670) := X"A202FFFE";
        ram_buffer(3671) := X"8E620008";
        ram_buffer(3672) := X"00000000";
        ram_buffer(3673) := X"00431021";
        ram_buffer(3674) := X"90420000";
        ram_buffer(3675) := X"1640FFEA";
        ram_buffer(3676) := X"A202FFFF";
        ram_buffer(3677) := X"8FBF0024";
        ram_buffer(3678) := X"8FB30020";
        ram_buffer(3679) := X"8FB2001C";
        ram_buffer(3680) := X"8FB10018";
        ram_buffer(3681) := X"8FB00014";
        ram_buffer(3682) := X"24020001";
        ram_buffer(3683) := X"03E00008";
        ram_buffer(3684) := X"27BD0028";
        ram_buffer(3685) := X"27BDFFD8";
        ram_buffer(3686) := X"8CA20010";
        ram_buffer(3687) := X"AFB30020";
        ram_buffer(3688) := X"8C930018";
        ram_buffer(3689) := X"AFB00014";
        ram_buffer(3690) := X"AFBF0024";
        ram_buffer(3691) := X"AFB2001C";
        ram_buffer(3692) := X"AFB10018";
        ram_buffer(3693) := X"8C500000";
        ram_buffer(3694) := X"1260001C";
        ram_buffer(3695) := X"3C12100D";
        ram_buffer(3696) := X"00A08821";
        ram_buffer(3697) := X"265282E8";
        ram_buffer(3698) := X"8E220028";
        ram_buffer(3699) := X"00000000";
        ram_buffer(3700) := X"0040F809";
        ram_buffer(3701) := X"02202021";
        ram_buffer(3702) := X"9222002D";
        ram_buffer(3703) := X"9223002C";
        ram_buffer(3704) := X"00021200";
        ram_buffer(3705) := X"00431021";
        ram_buffer(3706) := X"00022143";
        ram_buffer(3707) := X"00021A83";
        ram_buffer(3708) := X"3084001F";
        ram_buffer(3709) := X"3042001F";
        ram_buffer(3710) := X"3063001F";
        ram_buffer(3711) := X"02421021";
        ram_buffer(3712) := X"02442021";
        ram_buffer(3713) := X"02431821";
        ram_buffer(3714) := X"90450000";
        ram_buffer(3715) := X"90840000";
        ram_buffer(3716) := X"90620000";
        ram_buffer(3717) := X"2673FFFF";
        ram_buffer(3718) := X"A2050002";
        ram_buffer(3719) := X"A2040001";
        ram_buffer(3720) := X"A2020000";
        ram_buffer(3721) := X"1660FFE8";
        ram_buffer(3722) := X"26100003";
        ram_buffer(3723) := X"8FBF0024";
        ram_buffer(3724) := X"8FB30020";
        ram_buffer(3725) := X"8FB2001C";
        ram_buffer(3726) := X"8FB10018";
        ram_buffer(3727) := X"8FB00014";
        ram_buffer(3728) := X"24020001";
        ram_buffer(3729) := X"03E00008";
        ram_buffer(3730) := X"27BD0028";
        ram_buffer(3731) := X"27BDFFE0";
        ram_buffer(3732) := X"8CA20010";
        ram_buffer(3733) := X"AFB20018";
        ram_buffer(3734) := X"8C920018";
        ram_buffer(3735) := X"AFB10014";
        ram_buffer(3736) := X"AFBF001C";
        ram_buffer(3737) := X"AFB00010";
        ram_buffer(3738) := X"8C510000";
        ram_buffer(3739) := X"1240000E";
        ram_buffer(3740) := X"00A08021";
        ram_buffer(3741) := X"8E020028";
        ram_buffer(3742) := X"00000000";
        ram_buffer(3743) := X"0040F809";
        ram_buffer(3744) := X"02002021";
        ram_buffer(3745) := X"9202002E";
        ram_buffer(3746) := X"26310003";
        ram_buffer(3747) := X"A222FFFD";
        ram_buffer(3748) := X"9202002D";
        ram_buffer(3749) := X"2652FFFF";
        ram_buffer(3750) := X"A222FFFE";
        ram_buffer(3751) := X"9202002C";
        ram_buffer(3752) := X"1640FFF4";
        ram_buffer(3753) := X"A222FFFF";
        ram_buffer(3754) := X"8FBF001C";
        ram_buffer(3755) := X"8FB20018";
        ram_buffer(3756) := X"8FB10014";
        ram_buffer(3757) := X"8FB00010";
        ram_buffer(3758) := X"24020001";
        ram_buffer(3759) := X"03E00008";
        ram_buffer(3760) := X"27BD0020";
        ram_buffer(3761) := X"27BDFFE0";
        ram_buffer(3762) := X"8C830004";
        ram_buffer(3763) := X"8C82001C";
        ram_buffer(3764) := X"8CA60024";
        ram_buffer(3765) := X"AFB00018";
        ram_buffer(3766) := X"00A08021";
        ram_buffer(3767) := X"8CA50020";
        ram_buffer(3768) := X"AFA00010";
        ram_buffer(3769) := X"2442FFFF";
        ram_buffer(3770) := X"8C63001C";
        ram_buffer(3771) := X"AFBF001C";
        ram_buffer(3772) := X"24070001";
        ram_buffer(3773) := X"0060F809";
        ram_buffer(3774) := X"00463023";
        ram_buffer(3775) := X"8E030024";
        ram_buffer(3776) := X"8FBF001C";
        ram_buffer(3777) := X"24630001";
        ram_buffer(3778) := X"AE020010";
        ram_buffer(3779) := X"AE030024";
        ram_buffer(3780) := X"24020001";
        ram_buffer(3781) := X"8FB00018";
        ram_buffer(3782) := X"03E00008";
        ram_buffer(3783) := X"27BD0020";
        ram_buffer(3784) := X"8C86001C";
        ram_buffer(3785) := X"27BDFFD0";
        ram_buffer(3786) := X"AFB30024";
        ram_buffer(3787) := X"AFB1001C";
        ram_buffer(3788) := X"AFB00018";
        ram_buffer(3789) := X"AFBF002C";
        ram_buffer(3790) := X"AFB40028";
        ram_buffer(3791) := X"AFB20020";
        ram_buffer(3792) := X"00808021";
        ram_buffer(3793) := X"8C930008";
        ram_buffer(3794) := X"10C0004E";
        ram_buffer(3795) := X"00A08821";
        ram_buffer(3796) := X"00009021";
        ram_buffer(3797) := X"12600037";
        ram_buffer(3798) := X"24140001";
        ram_buffer(3799) := X"8E620000";
        ram_buffer(3800) := X"AE720004";
        ram_buffer(3801) := X"AE660008";
        ram_buffer(3802) := X"0040F809";
        ram_buffer(3803) := X"02002021";
        ram_buffer(3804) := X"8E020004";
        ram_buffer(3805) := X"8E250020";
        ram_buffer(3806) := X"AFB40010";
        ram_buffer(3807) := X"8C42001C";
        ram_buffer(3808) := X"02403021";
        ram_buffer(3809) := X"02002021";
        ram_buffer(3810) := X"0040F809";
        ram_buffer(3811) := X"24070001";
        ram_buffer(3812) := X"8E23003C";
        ram_buffer(3813) := X"AE220010";
        ram_buffer(3814) := X"02202821";
        ram_buffer(3815) := X"0060F809";
        ram_buffer(3816) := X"02002021";
        ram_buffer(3817) := X"8E06001C";
        ram_buffer(3818) := X"26520001";
        ram_buffer(3819) := X"0246102B";
        ram_buffer(3820) := X"1440FFEA";
        ram_buffer(3821) := X"00000000";
        ram_buffer(3822) := X"24C6FFFF";
        ram_buffer(3823) := X"12600005";
        ram_buffer(3824) := X"00000000";
        ram_buffer(3825) := X"8E620014";
        ram_buffer(3826) := X"00000000";
        ram_buffer(3827) := X"24420001";
        ram_buffer(3828) := X"AE620014";
        ram_buffer(3829) := X"8E020004";
        ram_buffer(3830) := X"8E250020";
        ram_buffer(3831) := X"AFA00010";
        ram_buffer(3832) := X"8C43001C";
        ram_buffer(3833) := X"3C021008";
        ram_buffer(3834) := X"24423AC4";
        ram_buffer(3835) := X"AE220004";
        ram_buffer(3836) := X"AE200024";
        ram_buffer(3837) := X"02002021";
        ram_buffer(3838) := X"0060F809";
        ram_buffer(3839) := X"24070001";
        ram_buffer(3840) := X"8E230024";
        ram_buffer(3841) := X"8FBF002C";
        ram_buffer(3842) := X"24630001";
        ram_buffer(3843) := X"AE220010";
        ram_buffer(3844) := X"AE230024";
        ram_buffer(3845) := X"8FB40028";
        ram_buffer(3846) := X"8FB30024";
        ram_buffer(3847) := X"8FB20020";
        ram_buffer(3848) := X"8FB1001C";
        ram_buffer(3849) := X"8FB00018";
        ram_buffer(3850) := X"24020001";
        ram_buffer(3851) := X"03E00008";
        ram_buffer(3852) := X"27BD0030";
        ram_buffer(3853) := X"8E020004";
        ram_buffer(3854) := X"8E250020";
        ram_buffer(3855) := X"AFB40010";
        ram_buffer(3856) := X"8C42001C";
        ram_buffer(3857) := X"02403021";
        ram_buffer(3858) := X"02002021";
        ram_buffer(3859) := X"0040F809";
        ram_buffer(3860) := X"24070001";
        ram_buffer(3861) := X"8E23003C";
        ram_buffer(3862) := X"AE220010";
        ram_buffer(3863) := X"02202821";
        ram_buffer(3864) := X"0060F809";
        ram_buffer(3865) := X"02002021";
        ram_buffer(3866) := X"8E06001C";
        ram_buffer(3867) := X"26520001";
        ram_buffer(3868) := X"0246102B";
        ram_buffer(3869) := X"1440FFEF";
        ram_buffer(3870) := X"24C6FFFF";
        ram_buffer(3871) := X"1000FFCF";
        ram_buffer(3872) := X"00000000";
        ram_buffer(3873) := X"1000FFCD";
        ram_buffer(3874) := X"2406FFFF";
        ram_buffer(3875) := X"03E00008";
        ram_buffer(3876) := X"00000000";
        ram_buffer(3877) := X"8C830030";
        ram_buffer(3878) := X"00000000";
        ram_buffer(3879) := X"18600047";
        ram_buffer(3880) := X"00000000";
        ram_buffer(3881) := X"27BDFFE0";
        ram_buffer(3882) := X"AFB00014";
        ram_buffer(3883) := X"8C90000C";
        ram_buffer(3884) := X"AFB10018";
        ram_buffer(3885) := X"8E020004";
        ram_buffer(3886) := X"AFBF001C";
        ram_buffer(3887) := X"2442FFFF";
        ram_buffer(3888) := X"00808821";
        ram_buffer(3889) := X"0440003F";
        ram_buffer(3890) := X"AE020004";
        ram_buffer(3891) := X"8E020000";
        ram_buffer(3892) := X"00000000";
        ram_buffer(3893) := X"24440001";
        ram_buffer(3894) := X"AE040000";
        ram_buffer(3895) := X"90440000";
        ram_buffer(3896) := X"28620002";
        ram_buffer(3897) := X"14400031";
        ram_buffer(3898) := X"A224002C";
        ram_buffer(3899) := X"8E020004";
        ram_buffer(3900) := X"00000000";
        ram_buffer(3901) := X"2442FFFF";
        ram_buffer(3902) := X"04400038";
        ram_buffer(3903) := X"AE020004";
        ram_buffer(3904) := X"8E020000";
        ram_buffer(3905) := X"00000000";
        ram_buffer(3906) := X"24440001";
        ram_buffer(3907) := X"AE040000";
        ram_buffer(3908) := X"90440000";
        ram_buffer(3909) := X"28620003";
        ram_buffer(3910) := X"14400024";
        ram_buffer(3911) := X"A224002D";
        ram_buffer(3912) := X"8E020004";
        ram_buffer(3913) := X"00000000";
        ram_buffer(3914) := X"2442FFFF";
        ram_buffer(3915) := X"04400031";
        ram_buffer(3916) := X"AE020004";
        ram_buffer(3917) := X"8E020000";
        ram_buffer(3918) := X"00000000";
        ram_buffer(3919) := X"24440001";
        ram_buffer(3920) := X"AE040000";
        ram_buffer(3921) := X"90440000";
        ram_buffer(3922) := X"28620004";
        ram_buffer(3923) := X"14400017";
        ram_buffer(3924) := X"A224002E";
        ram_buffer(3925) := X"8E020004";
        ram_buffer(3926) := X"00000000";
        ram_buffer(3927) := X"2442FFFF";
        ram_buffer(3928) := X"0440002A";
        ram_buffer(3929) := X"AE020004";
        ram_buffer(3930) := X"8E020000";
        ram_buffer(3931) := X"00000000";
        ram_buffer(3932) := X"24440001";
        ram_buffer(3933) := X"AE040000";
        ram_buffer(3934) := X"90420000";
        ram_buffer(3935) := X"28630005";
        ram_buffer(3936) := X"1460000A";
        ram_buffer(3937) := X"A222002F";
        ram_buffer(3938) := X"8E020004";
        ram_buffer(3939) := X"00000000";
        ram_buffer(3940) := X"2442FFFF";
        ram_buffer(3941) := X"04400023";
        ram_buffer(3942) := X"AE020004";
        ram_buffer(3943) := X"8E020000";
        ram_buffer(3944) := X"00000000";
        ram_buffer(3945) := X"24420001";
        ram_buffer(3946) := X"AE020000";
        ram_buffer(3947) := X"8FBF001C";
        ram_buffer(3948) := X"8FB10018";
        ram_buffer(3949) := X"8FB00014";
        ram_buffer(3950) := X"27BD0020";
        ram_buffer(3951) := X"03E00008";
        ram_buffer(3952) := X"00000000";
        ram_buffer(3953) := X"8F848098";
        ram_buffer(3954) := X"0C028350";
        ram_buffer(3955) := X"02002821";
        ram_buffer(3956) := X"8E230030";
        ram_buffer(3957) := X"1000FFC2";
        ram_buffer(3958) := X"304400FF";
        ram_buffer(3959) := X"8F848098";
        ram_buffer(3960) := X"0C028350";
        ram_buffer(3961) := X"02002821";
        ram_buffer(3962) := X"8E230030";
        ram_buffer(3963) := X"1000FFC9";
        ram_buffer(3964) := X"304400FF";
        ram_buffer(3965) := X"8F848098";
        ram_buffer(3966) := X"0C028350";
        ram_buffer(3967) := X"02002821";
        ram_buffer(3968) := X"8E230030";
        ram_buffer(3969) := X"1000FFD0";
        ram_buffer(3970) := X"304400FF";
        ram_buffer(3971) := X"8F848098";
        ram_buffer(3972) := X"0C028350";
        ram_buffer(3973) := X"02002821";
        ram_buffer(3974) := X"8E230030";
        ram_buffer(3975) := X"1000FFD7";
        ram_buffer(3976) := X"304200FF";
        ram_buffer(3977) := X"8F848098";
        ram_buffer(3978) := X"0C028350";
        ram_buffer(3979) := X"02002821";
        ram_buffer(3980) := X"8C820038";
        ram_buffer(3981) := X"00000000";
        ram_buffer(3982) := X"18400003";
        ram_buffer(3983) := X"2442FFFF";
        ram_buffer(3984) := X"03E00008";
        ram_buffer(3985) := X"AC820038";
        ram_buffer(3986) := X"8C820034";
        ram_buffer(3987) := X"27BDFFE0";
        ram_buffer(3988) := X"2442FFFF";
        ram_buffer(3989) := X"AFB10018";
        ram_buffer(3990) := X"AFB00014";
        ram_buffer(3991) := X"AFBF001C";
        ram_buffer(3992) := X"00808021";
        ram_buffer(3993) := X"8C91000C";
        ram_buffer(3994) := X"04400047";
        ram_buffer(3995) := X"AC820034";
        ram_buffer(3996) := X"8E030030";
        ram_buffer(3997) := X"00000000";
        ram_buffer(3998) := X"1860003E";
        ram_buffer(3999) := X"00000000";
        ram_buffer(4000) := X"8E220004";
        ram_buffer(4001) := X"00000000";
        ram_buffer(4002) := X"2442FFFF";
        ram_buffer(4003) := X"0440004E";
        ram_buffer(4004) := X"AE220004";
        ram_buffer(4005) := X"8E220000";
        ram_buffer(4006) := X"00000000";
        ram_buffer(4007) := X"24440001";
        ram_buffer(4008) := X"AE240000";
        ram_buffer(4009) := X"90440000";
        ram_buffer(4010) := X"28620002";
        ram_buffer(4011) := X"14400031";
        ram_buffer(4012) := X"A204002C";
        ram_buffer(4013) := X"8E220004";
        ram_buffer(4014) := X"00000000";
        ram_buffer(4015) := X"2442FFFF";
        ram_buffer(4016) := X"04400047";
        ram_buffer(4017) := X"AE220004";
        ram_buffer(4018) := X"8E220000";
        ram_buffer(4019) := X"00000000";
        ram_buffer(4020) := X"24440001";
        ram_buffer(4021) := X"AE240000";
        ram_buffer(4022) := X"90440000";
        ram_buffer(4023) := X"28620003";
        ram_buffer(4024) := X"14400024";
        ram_buffer(4025) := X"A204002D";
        ram_buffer(4026) := X"8E220004";
        ram_buffer(4027) := X"00000000";
        ram_buffer(4028) := X"2442FFFF";
        ram_buffer(4029) := X"04400040";
        ram_buffer(4030) := X"AE220004";
        ram_buffer(4031) := X"8E220000";
        ram_buffer(4032) := X"00000000";
        ram_buffer(4033) := X"24440001";
        ram_buffer(4034) := X"AE240000";
        ram_buffer(4035) := X"90440000";
        ram_buffer(4036) := X"28620004";
        ram_buffer(4037) := X"14400017";
        ram_buffer(4038) := X"A204002E";
        ram_buffer(4039) := X"8E220004";
        ram_buffer(4040) := X"00000000";
        ram_buffer(4041) := X"2442FFFF";
        ram_buffer(4042) := X"04400039";
        ram_buffer(4043) := X"AE220004";
        ram_buffer(4044) := X"8E220000";
        ram_buffer(4045) := X"00000000";
        ram_buffer(4046) := X"24440001";
        ram_buffer(4047) := X"AE240000";
        ram_buffer(4048) := X"90420000";
        ram_buffer(4049) := X"28630005";
        ram_buffer(4050) := X"1460000A";
        ram_buffer(4051) := X"A202002F";
        ram_buffer(4052) := X"8E220004";
        ram_buffer(4053) := X"00000000";
        ram_buffer(4054) := X"2442FFFF";
        ram_buffer(4055) := X"04400032";
        ram_buffer(4056) := X"AE220004";
        ram_buffer(4057) := X"8E220000";
        ram_buffer(4058) := X"00000000";
        ram_buffer(4059) := X"24420001";
        ram_buffer(4060) := X"AE220000";
        ram_buffer(4061) := X"8FBF001C";
        ram_buffer(4062) := X"8FB10018";
        ram_buffer(4063) := X"8FB00014";
        ram_buffer(4064) := X"03E00008";
        ram_buffer(4065) := X"27BD0020";
        ram_buffer(4066) := X"8E220004";
        ram_buffer(4067) := X"00000000";
        ram_buffer(4068) := X"2442FFFF";
        ram_buffer(4069) := X"04400027";
        ram_buffer(4070) := X"AE220004";
        ram_buffer(4071) := X"8E220000";
        ram_buffer(4072) := X"00000000";
        ram_buffer(4073) := X"24430001";
        ram_buffer(4074) := X"AE230000";
        ram_buffer(4075) := X"90420000";
        ram_buffer(4076) := X"00000000";
        ram_buffer(4077) := X"30430080";
        ram_buffer(4078) := X"1460002D";
        ram_buffer(4079) := X"3042007F";
        ram_buffer(4080) := X"1000FFAB";
        ram_buffer(4081) := X"AE020034";
        ram_buffer(4082) := X"8F848098";
        ram_buffer(4083) := X"0C028350";
        ram_buffer(4084) := X"02202821";
        ram_buffer(4085) := X"8E030030";
        ram_buffer(4086) := X"1000FFB3";
        ram_buffer(4087) := X"304400FF";
        ram_buffer(4088) := X"8F848098";
        ram_buffer(4089) := X"0C028350";
        ram_buffer(4090) := X"02202821";
        ram_buffer(4091) := X"8E030030";
        ram_buffer(4092) := X"1000FFBA";
        ram_buffer(4093) := X"304400FF";
        ram_buffer(4094) := X"8F848098";
        ram_buffer(4095) := X"0C028350";
        ram_buffer(4096) := X"02202821";
        ram_buffer(4097) := X"8E030030";
        ram_buffer(4098) := X"1000FFC1";
        ram_buffer(4099) := X"304400FF";
        ram_buffer(4100) := X"8F848098";
        ram_buffer(4101) := X"0C028350";
        ram_buffer(4102) := X"02202821";
        ram_buffer(4103) := X"8E030030";
        ram_buffer(4104) := X"1000FFC8";
        ram_buffer(4105) := X"304200FF";
        ram_buffer(4106) := X"8F848098";
        ram_buffer(4107) := X"0C028350";
        ram_buffer(4108) := X"02202821";
        ram_buffer(4109) := X"8F848098";
        ram_buffer(4110) := X"0C028350";
        ram_buffer(4111) := X"02202821";
        ram_buffer(4112) := X"2403FFFF";
        ram_buffer(4113) := X"1443FFDB";
        ram_buffer(4114) := X"2405002A";
        ram_buffer(4115) := X"8E040018";
        ram_buffer(4116) := X"00000000";
        ram_buffer(4117) := X"8C820000";
        ram_buffer(4118) := X"00000000";
        ram_buffer(4119) := X"8C430000";
        ram_buffer(4120) := X"00000000";
        ram_buffer(4121) := X"0060F809";
        ram_buffer(4122) := X"AC450014";
        ram_buffer(4123) := X"2402007F";
        ram_buffer(4124) := X"AE020038";
        ram_buffer(4125) := X"1000FF7E";
        ram_buffer(4126) := X"AE000034";
        ram_buffer(4127) := X"27BDFFA0";
        ram_buffer(4128) := X"8CA7000C";
        ram_buffer(4129) := X"24060012";
        ram_buffer(4130) := X"AFBE0058";
        ram_buffer(4131) := X"AFB00038";
        ram_buffer(4132) := X"00A0F021";
        ram_buffer(4133) := X"00808021";
        ram_buffer(4134) := X"24050001";
        ram_buffer(4135) := X"27A40018";
        ram_buffer(4136) := X"AFBF005C";
        ram_buffer(4137) := X"AFB70054";
        ram_buffer(4138) := X"AFB60050";
        ram_buffer(4139) := X"AFB5004C";
        ram_buffer(4140) := X"AFB40048";
        ram_buffer(4141) := X"AFB30044";
        ram_buffer(4142) := X"AFB20040";
        ram_buffer(4143) := X"0C0272E9";
        ram_buffer(4144) := X"AFB1003C";
        ram_buffer(4145) := X"24040012";
        ram_buffer(4146) := X"10440007";
        ram_buffer(4147) := X"2404002A";
        ram_buffer(4148) := X"8E020000";
        ram_buffer(4149) := X"00000000";
        ram_buffer(4150) := X"8C450000";
        ram_buffer(4151) := X"AC440014";
        ram_buffer(4152) := X"00A0F809";
        ram_buffer(4153) := X"02002021";
        ram_buffer(4154) := X"93A70028";
        ram_buffer(4155) := X"2402000F";
        ram_buffer(4156) := X"10E20170";
        ram_buffer(4157) := X"24020010";
        ram_buffer(4158) := X"000710C2";
        ram_buffer(4159) := X"00405021";
        ram_buffer(4160) := X"93B60019";
        ram_buffer(4161) := X"93A6001E";
        ram_buffer(4162) := X"93A50025";
        ram_buffer(4163) := X"93A40027";
        ram_buffer(4164) := X"93A80029";
        ram_buffer(4165) := X"93B2001D";
        ram_buffer(4166) := X"93B30024";
        ram_buffer(4167) := X"93B40026";
        ram_buffer(4168) := X"00063200";
        ram_buffer(4169) := X"00052A00";
        ram_buffer(4170) := X"00042200";
        ram_buffer(4171) := X"31150020";
        ram_buffer(4172) := X"2AC90002";
        ram_buffer(4173) := X"93B10018";
        ram_buffer(4174) := X"93B7001A";
        ram_buffer(4175) := X"00D29021";
        ram_buffer(4176) := X"00B39821";
        ram_buffer(4177) := X"0094A021";
        ram_buffer(4178) := X"AFCA0030";
        ram_buffer(4179) := X"1520014F";
        ram_buffer(4180) := X"32B500FF";
        ram_buffer(4181) := X"8E020000";
        ram_buffer(4182) := X"24040409";
        ram_buffer(4183) := X"8C450000";
        ram_buffer(4184) := X"AC440014";
        ram_buffer(4185) := X"00A0F809";
        ram_buffer(4186) := X"02002021";
        ram_buffer(4187) := X"2AE20009";
        ram_buffer(4188) := X"144000ED";
        ram_buffer(4189) := X"3C021008";
        ram_buffer(4190) := X"3C021008";
        ram_buffer(4191) := X"24423E30";
        ram_buffer(4192) := X"24040002";
        ram_buffer(4193) := X"26F7FFF8";
        ram_buffer(4194) := X"AFC00038";
        ram_buffer(4195) := X"AFC00034";
        ram_buffer(4196) := X"AFC20028";
        ram_buffer(4197) := X"12E400E9";
        ram_buffer(4198) := X"AE040024";
        ram_buffer(4199) := X"24020003";
        ram_buffer(4200) := X"12E20149";
        ram_buffer(4201) := X"24020001";
        ram_buffer(4202) := X"12E200F9";
        ram_buffer(4203) := X"24040409";
        ram_buffer(4204) := X"8E020000";
        ram_buffer(4205) := X"00000000";
        ram_buffer(4206) := X"8C450000";
        ram_buffer(4207) := X"AC440014";
        ram_buffer(4208) := X"00A0F809";
        ram_buffer(4209) := X"02002021";
        ram_buffer(4210) := X"24020003";
        ram_buffer(4211) := X"24060003";
        ram_buffer(4212) := X"AFA20034";
        ram_buffer(4213) := X"16A00109";
        ram_buffer(4214) := X"02660018";
        ram_buffer(4215) := X"8E020004";
        ram_buffer(4216) := X"24040001";
        ram_buffer(4217) := X"AFA40014";
        ram_buffer(4218) := X"AFB40010";
        ram_buffer(4219) := X"8C420010";
        ram_buffer(4220) := X"02002021";
        ram_buffer(4221) := X"00003021";
        ram_buffer(4222) := X"00003812";
        ram_buffer(4223) := X"0040F809";
        ram_buffer(4224) := X"24050001";
        ram_buffer(4225) := X"8E040008";
        ram_buffer(4226) := X"00000000";
        ram_buffer(4227) := X"10800005";
        ram_buffer(4228) := X"AFC20020";
        ram_buffer(4229) := X"8C820018";
        ram_buffer(4230) := X"00000000";
        ram_buffer(4231) := X"24420001";
        ram_buffer(4232) := X"AC820018";
        ram_buffer(4233) := X"24020001";
        ram_buffer(4234) := X"AFC20014";
        ram_buffer(4235) := X"3C021008";
        ram_buffer(4236) := X"24423B20";
        ram_buffer(4237) := X"AFC20004";
        ram_buffer(4238) := X"0000B821";
        ram_buffer(4239) := X"2415002A";
        ram_buffer(4240) := X"1237000F";
        ram_buffer(4241) := X"00000000";
        ram_buffer(4242) := X"8FC5000C";
        ram_buffer(4243) := X"00000000";
        ram_buffer(4244) := X"8CA20004";
        ram_buffer(4245) := X"00000000";
        ram_buffer(4246) := X"2442FFFF";
        ram_buffer(4247) := X"044000F7";
        ram_buffer(4248) := X"ACA20004";
        ram_buffer(4249) := X"8CA20000";
        ram_buffer(4250) := X"00000000";
        ram_buffer(4251) := X"24420001";
        ram_buffer(4252) := X"ACA20000";
        ram_buffer(4253) := X"26F70001";
        ram_buffer(4254) := X"1637FFF3";
        ram_buffer(4255) := X"00000000";
        ram_buffer(4256) := X"124000FE";
        ram_buffer(4257) := X"2E420101";
        ram_buffer(4258) := X"10400007";
        ram_buffer(4259) := X"00000000";
        ram_buffer(4260) := X"93A2001C";
        ram_buffer(4261) := X"93A4001B";
        ram_buffer(4262) := X"00021200";
        ram_buffer(4263) := X"00441021";
        ram_buffer(4264) := X"10400007";
        ram_buffer(4265) := X"00000000";
        ram_buffer(4266) := X"8E020000";
        ram_buffer(4267) := X"24040408";
        ram_buffer(4268) := X"8C450000";
        ram_buffer(4269) := X"AC440014";
        ram_buffer(4270) := X"00A0F809";
        ram_buffer(4271) := X"02002021";
        ram_buffer(4272) := X"8E020004";
        ram_buffer(4273) := X"24050001";
        ram_buffer(4274) := X"8C420008";
        ram_buffer(4275) := X"02002021";
        ram_buffer(4276) := X"24070003";
        ram_buffer(4277) := X"0040F809";
        ram_buffer(4278) := X"02403021";
        ram_buffer(4279) := X"93A5001F";
        ram_buffer(4280) := X"24040018";
        ram_buffer(4281) := X"10A4000A";
        ram_buffer(4282) := X"AFC2001C";
        ram_buffer(4283) := X"8FC40018";
        ram_buffer(4284) := X"24060408";
        ram_buffer(4285) := X"8C820000";
        ram_buffer(4286) := X"00000000";
        ram_buffer(4287) := X"8C450000";
        ram_buffer(4288) := X"00000000";
        ram_buffer(4289) := X"00A0F809";
        ram_buffer(4290) := X"AC460014";
        ram_buffer(4291) := X"8FC2001C";
        ram_buffer(4292) := X"00008821";
        ram_buffer(4293) := X"2416FFFF";
        ram_buffer(4294) := X"10000029";
        ram_buffer(4295) := X"2415002A";
        ram_buffer(4296) := X"8CA20000";
        ram_buffer(4297) := X"00000000";
        ram_buffer(4298) := X"24440001";
        ram_buffer(4299) := X"ACA40000";
        ram_buffer(4300) := X"90420000";
        ram_buffer(4301) := X"00000000";
        ram_buffer(4302) := X"A2E20000";
        ram_buffer(4303) := X"8FC5000C";
        ram_buffer(4304) := X"8FC4001C";
        ram_buffer(4305) := X"8CA20004";
        ram_buffer(4306) := X"8C970004";
        ram_buffer(4307) := X"2442FFFF";
        ram_buffer(4308) := X"02F1B821";
        ram_buffer(4309) := X"04400039";
        ram_buffer(4310) := X"ACA20004";
        ram_buffer(4311) := X"8CA20000";
        ram_buffer(4312) := X"00000000";
        ram_buffer(4313) := X"24440001";
        ram_buffer(4314) := X"ACA40000";
        ram_buffer(4315) := X"90420000";
        ram_buffer(4316) := X"00000000";
        ram_buffer(4317) := X"A2E20000";
        ram_buffer(4318) := X"8FC5000C";
        ram_buffer(4319) := X"8FC4001C";
        ram_buffer(4320) := X"8CA20004";
        ram_buffer(4321) := X"8C970000";
        ram_buffer(4322) := X"2442FFFF";
        ram_buffer(4323) := X"02F1B821";
        ram_buffer(4324) := X"04400042";
        ram_buffer(4325) := X"ACA20004";
        ram_buffer(4326) := X"8CA20000";
        ram_buffer(4327) := X"00000000";
        ram_buffer(4328) := X"24440001";
        ram_buffer(4329) := X"ACA40000";
        ram_buffer(4330) := X"90420000";
        ram_buffer(4331) := X"26310001";
        ram_buffer(4332) := X"0232202A";
        ram_buffer(4333) := X"1080004A";
        ram_buffer(4334) := X"A2E20000";
        ram_buffer(4335) := X"8FC2001C";
        ram_buffer(4336) := X"8FC5000C";
        ram_buffer(4337) := X"8C570008";
        ram_buffer(4338) := X"8CA20004";
        ram_buffer(4339) := X"02F1B821";
        ram_buffer(4340) := X"2442FFFF";
        ram_buffer(4341) := X"0441FFD2";
        ram_buffer(4342) := X"ACA20004";
        ram_buffer(4343) := X"8F848098";
        ram_buffer(4344) := X"0C028350";
        ram_buffer(4345) := X"00000000";
        ram_buffer(4346) := X"1456FFD3";
        ram_buffer(4347) := X"00000000";
        ram_buffer(4348) := X"8FC40018";
        ram_buffer(4349) := X"AFA20030";
        ram_buffer(4350) := X"8C850000";
        ram_buffer(4351) := X"00000000";
        ram_buffer(4352) := X"8CA60000";
        ram_buffer(4353) := X"00000000";
        ram_buffer(4354) := X"00C0F809";
        ram_buffer(4355) := X"ACB50014";
        ram_buffer(4356) := X"8FA20030";
        ram_buffer(4357) := X"00000000";
        ram_buffer(4358) := X"A2E20000";
        ram_buffer(4359) := X"8FC5000C";
        ram_buffer(4360) := X"8FC4001C";
        ram_buffer(4361) := X"8CA20004";
        ram_buffer(4362) := X"8C970004";
        ram_buffer(4363) := X"2442FFFF";
        ram_buffer(4364) := X"02F1B821";
        ram_buffer(4365) := X"0441FFC9";
        ram_buffer(4366) := X"ACA20004";
        ram_buffer(4367) := X"8F848098";
        ram_buffer(4368) := X"0C028350";
        ram_buffer(4369) := X"00000000";
        ram_buffer(4370) := X"1456FFCA";
        ram_buffer(4371) := X"00000000";
        ram_buffer(4372) := X"8FC40018";
        ram_buffer(4373) := X"AFA20030";
        ram_buffer(4374) := X"8C850000";
        ram_buffer(4375) := X"00000000";
        ram_buffer(4376) := X"8CA60000";
        ram_buffer(4377) := X"00000000";
        ram_buffer(4378) := X"00C0F809";
        ram_buffer(4379) := X"ACB50014";
        ram_buffer(4380) := X"8FA20030";
        ram_buffer(4381) := X"00000000";
        ram_buffer(4382) := X"A2E20000";
        ram_buffer(4383) := X"8FC5000C";
        ram_buffer(4384) := X"8FC4001C";
        ram_buffer(4385) := X"8CA20004";
        ram_buffer(4386) := X"8C970000";
        ram_buffer(4387) := X"2442FFFF";
        ram_buffer(4388) := X"02F1B821";
        ram_buffer(4389) := X"0441FFC0";
        ram_buffer(4390) := X"ACA20004";
        ram_buffer(4391) := X"8F848098";
        ram_buffer(4392) := X"0C028350";
        ram_buffer(4393) := X"00000000";
        ram_buffer(4394) := X"1456FFC0";
        ram_buffer(4395) := X"00000000";
        ram_buffer(4396) := X"8FC40018";
        ram_buffer(4397) := X"AFA20030";
        ram_buffer(4398) := X"8C850000";
        ram_buffer(4399) := X"26310001";
        ram_buffer(4400) := X"8CA60000";
        ram_buffer(4401) := X"00000000";
        ram_buffer(4402) := X"00C0F809";
        ram_buffer(4403) := X"ACB50014";
        ram_buffer(4404) := X"8FA20030";
        ram_buffer(4405) := X"0232202A";
        ram_buffer(4406) := X"1480FFB8";
        ram_buffer(4407) := X"A2E20000";
        ram_buffer(4408) := X"8FA20034";
        ram_buffer(4409) := X"8FBF005C";
        ram_buffer(4410) := X"AE020020";
        ram_buffer(4411) := X"24020008";
        ram_buffer(4412) := X"AE130018";
        ram_buffer(4413) := X"AE14001C";
        ram_buffer(4414) := X"AE020030";
        ram_buffer(4415) := X"8FBE0058";
        ram_buffer(4416) := X"8FB70054";
        ram_buffer(4417) := X"8FB60050";
        ram_buffer(4418) := X"8FB5004C";
        ram_buffer(4419) := X"8FB40048";
        ram_buffer(4420) := X"8FB30044";
        ram_buffer(4421) := X"8FB20040";
        ram_buffer(4422) := X"8FB1003C";
        ram_buffer(4423) := X"8FB00038";
        ram_buffer(4424) := X"03E00008";
        ram_buffer(4425) := X"27BD0060";
        ram_buffer(4426) := X"24423C94";
        ram_buffer(4427) := X"24040002";
        ram_buffer(4428) := X"AFC20028";
        ram_buffer(4429) := X"16E4FF19";
        ram_buffer(4430) := X"AE040024";
        ram_buffer(4431) := X"8FC20030";
        ram_buffer(4432) := X"24040003";
        ram_buffer(4433) := X"1044008B";
        ram_buffer(4434) := X"00000000";
        ram_buffer(4435) := X"24040004";
        ram_buffer(4436) := X"10440088";
        ram_buffer(4437) := X"00000000";
        ram_buffer(4438) := X"1057008A";
        ram_buffer(4439) := X"00000000";
        ram_buffer(4440) := X"8E020000";
        ram_buffer(4441) := X"24040409";
        ram_buffer(4442) := X"8C450000";
        ram_buffer(4443) := X"AC440014";
        ram_buffer(4444) := X"00A0F809";
        ram_buffer(4445) := X"02002021";
        ram_buffer(4446) := X"8E020000";
        ram_buffer(4447) := X"00000000";
        ram_buffer(4448) := X"AC530018";
        ram_buffer(4449) := X"8E040000";
        ram_buffer(4450) := X"1000000F";
        ram_buffer(4451) := X"2405040B";
        ram_buffer(4452) := X"8FC20030";
        ram_buffer(4453) := X"00000000";
        ram_buffer(4454) := X"10570071";
        ram_buffer(4455) := X"00000000";
        ram_buffer(4456) := X"8E020000";
        ram_buffer(4457) := X"24040409";
        ram_buffer(4458) := X"8C450000";
        ram_buffer(4459) := X"AC440014";
        ram_buffer(4460) := X"00A0F809";
        ram_buffer(4461) := X"02002021";
        ram_buffer(4462) := X"8E020000";
        ram_buffer(4463) := X"2405040D";
        ram_buffer(4464) := X"AC530018";
        ram_buffer(4465) := X"8E040000";
        ram_buffer(4466) := X"AC450014";
        ram_buffer(4467) := X"AC94001C";
        ram_buffer(4468) := X"8E020000";
        ram_buffer(4469) := X"24050001";
        ram_buffer(4470) := X"8C420004";
        ram_buffer(4471) := X"00000000";
        ram_buffer(4472) := X"0040F809";
        ram_buffer(4473) := X"02002021";
        ram_buffer(4474) := X"24060003";
        ram_buffer(4475) := X"24020003";
        ram_buffer(4476) := X"AFA20034";
        ram_buffer(4477) := X"12A0FEF9";
        ram_buffer(4478) := X"02660018";
        ram_buffer(4479) := X"8E020004";
        ram_buffer(4480) := X"02002021";
        ram_buffer(4481) := X"8C420008";
        ram_buffer(4482) := X"AFC00020";
        ram_buffer(4483) := X"24070001";
        ram_buffer(4484) := X"24050001";
        ram_buffer(4485) := X"0000B821";
        ram_buffer(4486) := X"00003012";
        ram_buffer(4487) := X"0040F809";
        ram_buffer(4488) := X"2415002A";
        ram_buffer(4489) := X"8FC4003C";
        ram_buffer(4490) := X"AFC20010";
        ram_buffer(4491) := X"24020001";
        ram_buffer(4492) := X"AFC20014";
        ram_buffer(4493) := X"1000FF02";
        ram_buffer(4494) := X"AFC40004";
        ram_buffer(4495) := X"8F848098";
        ram_buffer(4496) := X"0C028350";
        ram_buffer(4497) := X"00000000";
        ram_buffer(4498) := X"2403FFFF";
        ram_buffer(4499) := X"1443FF09";
        ram_buffer(4500) := X"00000000";
        ram_buffer(4501) := X"8FC40018";
        ram_buffer(4502) := X"26F70001";
        ram_buffer(4503) := X"8C820000";
        ram_buffer(4504) := X"00000000";
        ram_buffer(4505) := X"8C450000";
        ram_buffer(4506) := X"00000000";
        ram_buffer(4507) := X"00A0F809";
        ram_buffer(4508) := X"AC550014";
        ram_buffer(4509) := X"1000FF00";
        ram_buffer(4510) := X"00000000";
        ram_buffer(4511) := X"16C0002C";
        ram_buffer(4512) := X"24040409";
        ram_buffer(4513) := X"1000FF96";
        ram_buffer(4514) := X"AFC0001C";
        ram_buffer(4515) := X"2442FFFF";
        ram_buffer(4516) := X"2C420004";
        ram_buffer(4517) := X"1040FEAF";
        ram_buffer(4518) := X"30E70007";
        ram_buffer(4519) := X"14E0FEAD";
        ram_buffer(4520) := X"00084183";
        ram_buffer(4521) := X"1100FEB2";
        ram_buffer(4522) := X"2AE20009";
        ram_buffer(4523) := X"1000FEA9";
        ram_buffer(4524) := X"00000000";
        ram_buffer(4525) := X"A3A20028";
        ram_buffer(4526) := X"240A0002";
        ram_buffer(4527) := X"24020002";
        ram_buffer(4528) := X"1000FE8F";
        ram_buffer(4529) := X"24070010";
        ram_buffer(4530) := X"8FC40030";
        ram_buffer(4531) := X"00000000";
        ram_buffer(4532) := X"1082001F";
        ram_buffer(4533) := X"AE020024";
        ram_buffer(4534) := X"8E020000";
        ram_buffer(4535) := X"24040409";
        ram_buffer(4536) := X"8C450000";
        ram_buffer(4537) := X"AC440014";
        ram_buffer(4538) := X"00A0F809";
        ram_buffer(4539) := X"02002021";
        ram_buffer(4540) := X"8E020000";
        ram_buffer(4541) := X"2405040C";
        ram_buffer(4542) := X"AC530018";
        ram_buffer(4543) := X"8E040000";
        ram_buffer(4544) := X"AC450014";
        ram_buffer(4545) := X"AC94001C";
        ram_buffer(4546) := X"8E020000";
        ram_buffer(4547) := X"24050001";
        ram_buffer(4548) := X"8C420004";
        ram_buffer(4549) := X"00000000";
        ram_buffer(4550) := X"0040F809";
        ram_buffer(4551) := X"02002021";
        ram_buffer(4552) := X"24020001";
        ram_buffer(4553) := X"24060001";
        ram_buffer(4554) := X"1000FEAA";
        ram_buffer(4555) := X"AFA20034";
        ram_buffer(4556) := X"8E020000";
        ram_buffer(4557) := X"00000000";
        ram_buffer(4558) := X"8C450000";
        ram_buffer(4559) := X"AC440014";
        ram_buffer(4560) := X"00A0F809";
        ram_buffer(4561) := X"02002021";
        ram_buffer(4562) := X"1000FF65";
        ram_buffer(4563) := X"AFC0001C";
        ram_buffer(4564) := X"3C021008";
        ram_buffer(4565) := X"24423880";
        ram_buffer(4566) := X"1000FFE5";
        ram_buffer(4567) := X"AFC2003C";
        ram_buffer(4568) := X"16D7FF8F";
        ram_buffer(4569) := X"3C021008";
        ram_buffer(4570) := X"244238E8";
        ram_buffer(4571) := X"1000FF92";
        ram_buffer(4572) := X"AFC2003C";
        ram_buffer(4573) := X"3C021008";
        ram_buffer(4574) := X"24423A4C";
        ram_buffer(4575) := X"1000FF7E";
        ram_buffer(4576) := X"AFC2003C";
        ram_buffer(4577) := X"3C021008";
        ram_buffer(4578) := X"24423994";
        ram_buffer(4579) := X"1000FF7A";
        ram_buffer(4580) := X"AFC2003C";
        ram_buffer(4581) := X"8C820004";
        ram_buffer(4582) := X"27BDFFE8";
        ram_buffer(4583) := X"8C420000";
        ram_buffer(4584) := X"24060040";
        ram_buffer(4585) := X"AFBF0014";
        ram_buffer(4586) := X"AFB00010";
        ram_buffer(4587) := X"24050001";
        ram_buffer(4588) := X"0040F809";
        ram_buffer(4589) := X"00808021";
        ram_buffer(4590) := X"3C041008";
        ram_buffer(4591) := X"2484407C";
        ram_buffer(4592) := X"AC440000";
        ram_buffer(4593) := X"8FBF0014";
        ram_buffer(4594) := X"3C041008";
        ram_buffer(4595) := X"24843C8C";
        ram_buffer(4596) := X"AC500018";
        ram_buffer(4597) := X"AC440008";
        ram_buffer(4598) := X"8FB00010";
        ram_buffer(4599) := X"03E00008";
        ram_buffer(4600) := X"27BD0018";
        ram_buffer(4601) := X"27BDFFD8";
        ram_buffer(4602) := X"8CA60024";
        ram_buffer(4603) := X"8C820004";
        ram_buffer(4604) := X"AFB1001C";
        ram_buffer(4605) := X"00A08821";
        ram_buffer(4606) := X"8CA50020";
        ram_buffer(4607) := X"AFA00010";
        ram_buffer(4608) := X"24C6FFFF";
        ram_buffer(4609) := X"8C42001C";
        ram_buffer(4610) := X"AFB20020";
        ram_buffer(4611) := X"AFB00018";
        ram_buffer(4612) := X"AFBF0024";
        ram_buffer(4613) := X"24070001";
        ram_buffer(4614) := X"AE260024";
        ram_buffer(4615) := X"8E30001C";
        ram_buffer(4616) := X"0040F809";
        ram_buffer(4617) := X"00809021";
        ram_buffer(4618) := X"8C430000";
        ram_buffer(4619) := X"8E440018";
        ram_buffer(4620) := X"8E220010";
        ram_buffer(4621) := X"00000000";
        ram_buffer(4622) := X"8C420000";
        ram_buffer(4623) := X"10800015";
        ram_buffer(4624) := X"00643021";
        ram_buffer(4625) := X"24630001";
        ram_buffer(4626) := X"9065FFFF";
        ram_buffer(4627) := X"8E040000";
        ram_buffer(4628) := X"24420003";
        ram_buffer(4629) := X"00852021";
        ram_buffer(4630) := X"90840000";
        ram_buffer(4631) := X"00000000";
        ram_buffer(4632) := X"A044FFFD";
        ram_buffer(4633) := X"8E040004";
        ram_buffer(4634) := X"00000000";
        ram_buffer(4635) := X"00852021";
        ram_buffer(4636) := X"90840000";
        ram_buffer(4637) := X"00000000";
        ram_buffer(4638) := X"A044FFFE";
        ram_buffer(4639) := X"8E040008";
        ram_buffer(4640) := X"00000000";
        ram_buffer(4641) := X"00852021";
        ram_buffer(4642) := X"90840000";
        ram_buffer(4643) := X"1466FFED";
        ram_buffer(4644) := X"A044FFFF";
        ram_buffer(4645) := X"8FBF0024";
        ram_buffer(4646) := X"8FB20020";
        ram_buffer(4647) := X"8FB1001C";
        ram_buffer(4648) := X"8FB00018";
        ram_buffer(4649) := X"24020001";
        ram_buffer(4650) := X"03E00008";
        ram_buffer(4651) := X"27BD0028";
        ram_buffer(4652) := X"27BDFFD8";
        ram_buffer(4653) := X"8CA60024";
        ram_buffer(4654) := X"8C820004";
        ram_buffer(4655) := X"AFB0001C";
        ram_buffer(4656) := X"00A08021";
        ram_buffer(4657) := X"8CA50020";
        ram_buffer(4658) := X"AFA00010";
        ram_buffer(4659) := X"24C6FFFF";
        ram_buffer(4660) := X"8C42001C";
        ram_buffer(4661) := X"AFB10020";
        ram_buffer(4662) := X"AFBF0024";
        ram_buffer(4663) := X"00808821";
        ram_buffer(4664) := X"AE060024";
        ram_buffer(4665) := X"0040F809";
        ram_buffer(4666) := X"24070001";
        ram_buffer(4667) := X"8E030010";
        ram_buffer(4668) := X"8E250018";
        ram_buffer(4669) := X"8C420000";
        ram_buffer(4670) := X"8C630000";
        ram_buffer(4671) := X"10A0000D";
        ram_buffer(4672) := X"00000000";
        ram_buffer(4673) := X"00052040";
        ram_buffer(4674) := X"00852821";
        ram_buffer(4675) := X"00452821";
        ram_buffer(4676) := X"90440000";
        ram_buffer(4677) := X"24420003";
        ram_buffer(4678) := X"A0640002";
        ram_buffer(4679) := X"9044FFFE";
        ram_buffer(4680) := X"24630003";
        ram_buffer(4681) := X"A064FFFE";
        ram_buffer(4682) := X"9044FFFF";
        ram_buffer(4683) := X"14A2FFF8";
        ram_buffer(4684) := X"A064FFFD";
        ram_buffer(4685) := X"8FBF0024";
        ram_buffer(4686) := X"8FB10020";
        ram_buffer(4687) := X"8FB0001C";
        ram_buffer(4688) := X"24020001";
        ram_buffer(4689) := X"03E00008";
        ram_buffer(4690) := X"27BD0028";
        ram_buffer(4691) := X"03E00008";
        ram_buffer(4692) := X"00000000";
        ram_buffer(4693) := X"8C82001C";
        ram_buffer(4694) := X"27BDFFC0";
        ram_buffer(4695) := X"AFB70034";
        ram_buffer(4696) := X"AFB30024";
        ram_buffer(4697) := X"AFB20020";
        ram_buffer(4698) := X"AFB00018";
        ram_buffer(4699) := X"AFBF003C";
        ram_buffer(4700) := X"AFBE0038";
        ram_buffer(4701) := X"AFB60030";
        ram_buffer(4702) := X"AFB5002C";
        ram_buffer(4703) := X"AFB40028";
        ram_buffer(4704) := X"AFB1001C";
        ram_buffer(4705) := X"00808021";
        ram_buffer(4706) := X"8CB7000C";
        ram_buffer(4707) := X"8C920008";
        ram_buffer(4708) := X"1040003B";
        ram_buffer(4709) := X"00A09821";
        ram_buffer(4710) := X"00008821";
        ram_buffer(4711) := X"2414002A";
        ram_buffer(4712) := X"12400006";
        ram_buffer(4713) := X"00000000";
        ram_buffer(4714) := X"8E430000";
        ram_buffer(4715) := X"AE510004";
        ram_buffer(4716) := X"AE420008";
        ram_buffer(4717) := X"0060F809";
        ram_buffer(4718) := X"02002021";
        ram_buffer(4719) := X"8E020004";
        ram_buffer(4720) := X"24030001";
        ram_buffer(4721) := X"8E650020";
        ram_buffer(4722) := X"AFA30010";
        ram_buffer(4723) := X"8C42001C";
        ram_buffer(4724) := X"24070001";
        ram_buffer(4725) := X"02203021";
        ram_buffer(4726) := X"0040F809";
        ram_buffer(4727) := X"02002021";
        ram_buffer(4728) := X"8E7E0028";
        ram_buffer(4729) := X"8C560000";
        ram_buffer(4730) := X"17C0000C";
        ram_buffer(4731) := X"00000000";
        ram_buffer(4732) := X"1000001E";
        ram_buffer(4733) := X"00000000";
        ram_buffer(4734) := X"8EE20000";
        ram_buffer(4735) := X"00000000";
        ram_buffer(4736) := X"24440001";
        ram_buffer(4737) := X"AEE40000";
        ram_buffer(4738) := X"90550000";
        ram_buffer(4739) := X"26D60001";
        ram_buffer(4740) := X"27DEFFFF";
        ram_buffer(4741) := X"13C00015";
        ram_buffer(4742) := X"A2D5FFFF";
        ram_buffer(4743) := X"8EE20004";
        ram_buffer(4744) := X"00000000";
        ram_buffer(4745) := X"2442FFFF";
        ram_buffer(4746) := X"0441FFF3";
        ram_buffer(4747) := X"AEE20004";
        ram_buffer(4748) := X"8F848098";
        ram_buffer(4749) := X"0C028350";
        ram_buffer(4750) := X"02E02821";
        ram_buffer(4751) := X"0040A821";
        ram_buffer(4752) := X"2402FFFF";
        ram_buffer(4753) := X"16A2FFF1";
        ram_buffer(4754) := X"02002021";
        ram_buffer(4755) := X"8E050000";
        ram_buffer(4756) := X"26D60001";
        ram_buffer(4757) := X"8CA60000";
        ram_buffer(4758) := X"ACB40014";
        ram_buffer(4759) := X"00C0F809";
        ram_buffer(4760) := X"27DEFFFF";
        ram_buffer(4761) := X"17C0FFED";
        ram_buffer(4762) := X"A2D5FFFF";
        ram_buffer(4763) := X"8E02001C";
        ram_buffer(4764) := X"26310001";
        ram_buffer(4765) := X"0222182B";
        ram_buffer(4766) := X"1460FFC9";
        ram_buffer(4767) := X"00000000";
        ram_buffer(4768) := X"12400005";
        ram_buffer(4769) := X"00000000";
        ram_buffer(4770) := X"8E430014";
        ram_buffer(4771) := X"00000000";
        ram_buffer(4772) := X"24630001";
        ram_buffer(4773) := X"AE430014";
        ram_buffer(4774) := X"8E63002C";
        ram_buffer(4775) := X"24040008";
        ram_buffer(4776) := X"1064001E";
        ram_buffer(4777) := X"24040018";
        ram_buffer(4778) := X"10640019";
        ram_buffer(4779) := X"3C191008";
        ram_buffer(4780) := X"8E020000";
        ram_buffer(4781) := X"240403EA";
        ram_buffer(4782) := X"8C430000";
        ram_buffer(4783) := X"AC440014";
        ram_buffer(4784) := X"0060F809";
        ram_buffer(4785) := X"02002021";
        ram_buffer(4786) := X"8E790004";
        ram_buffer(4787) := X"8E02001C";
        ram_buffer(4788) := X"00000000";
        ram_buffer(4789) := X"AE620024";
        ram_buffer(4790) := X"8FBF003C";
        ram_buffer(4791) := X"8FBE0038";
        ram_buffer(4792) := X"8FB70034";
        ram_buffer(4793) := X"8FB60030";
        ram_buffer(4794) := X"8FB5002C";
        ram_buffer(4795) := X"8FB40028";
        ram_buffer(4796) := X"8FB20020";
        ram_buffer(4797) := X"8FB1001C";
        ram_buffer(4798) := X"02602821";
        ram_buffer(4799) := X"02002021";
        ram_buffer(4800) := X"8FB30024";
        ram_buffer(4801) := X"8FB00018";
        ram_buffer(4802) := X"03200008";
        ram_buffer(4803) := X"27BD0040";
        ram_buffer(4804) := X"273948B0";
        ram_buffer(4805) := X"1000FFEF";
        ram_buffer(4806) := X"AE790004";
        ram_buffer(4807) := X"3C191008";
        ram_buffer(4808) := X"273947E4";
        ram_buffer(4809) := X"1000FFEB";
        ram_buffer(4810) := X"AE790004";
        ram_buffer(4811) := X"27BDFF58";
        ram_buffer(4812) := X"8CA7000C";
        ram_buffer(4813) := X"2406000E";
        ram_buffer(4814) := X"AFB20088";
        ram_buffer(4815) := X"AFB00080";
        ram_buffer(4816) := X"00809021";
        ram_buffer(4817) := X"00A08021";
        ram_buffer(4818) := X"27A40058";
        ram_buffer(4819) := X"24050001";
        ram_buffer(4820) := X"AFBF00A4";
        ram_buffer(4821) := X"AFBE00A0";
        ram_buffer(4822) := X"AFB7009C";
        ram_buffer(4823) := X"AFB60098";
        ram_buffer(4824) := X"AFB50094";
        ram_buffer(4825) := X"AFB40090";
        ram_buffer(4826) := X"AFB3008C";
        ram_buffer(4827) := X"0C0272E9";
        ram_buffer(4828) := X"AFB10084";
        ram_buffer(4829) := X"2403000E";
        ram_buffer(4830) := X"10430007";
        ram_buffer(4831) := X"00000000";
        ram_buffer(4832) := X"8E420000";
        ram_buffer(4833) := X"2404002A";
        ram_buffer(4834) := X"8C430000";
        ram_buffer(4835) := X"AC440014";
        ram_buffer(4836) := X"0060F809";
        ram_buffer(4837) := X"02402021";
        ram_buffer(4838) := X"93A20059";
        ram_buffer(4839) := X"93A30058";
        ram_buffer(4840) := X"00021200";
        ram_buffer(4841) := X"00431021";
        ram_buffer(4842) := X"24034D42";
        ram_buffer(4843) := X"10430007";
        ram_buffer(4844) := X"240403EF";
        ram_buffer(4845) := X"8E420000";
        ram_buffer(4846) := X"00000000";
        ram_buffer(4847) := X"8C430000";
        ram_buffer(4848) := X"AC440014";
        ram_buffer(4849) := X"0060F809";
        ram_buffer(4850) := X"02402021";
        ram_buffer(4851) := X"93A30063";
        ram_buffer(4852) := X"93A40062";
        ram_buffer(4853) := X"93A20064";
        ram_buffer(4854) := X"93B30065";
        ram_buffer(4855) := X"00031A00";
        ram_buffer(4856) := X"00641821";
        ram_buffer(4857) := X"00021400";
        ram_buffer(4858) := X"8E07000C";
        ram_buffer(4859) := X"00621021";
        ram_buffer(4860) := X"00139E00";
        ram_buffer(4861) := X"24060004";
        ram_buffer(4862) := X"24050001";
        ram_buffer(4863) := X"27A40018";
        ram_buffer(4864) := X"0C0272E9";
        ram_buffer(4865) := X"00539821";
        ram_buffer(4866) := X"24030004";
        ram_buffer(4867) := X"10430007";
        ram_buffer(4868) := X"2404002A";
        ram_buffer(4869) := X"8E420000";
        ram_buffer(4870) := X"00000000";
        ram_buffer(4871) := X"8C430000";
        ram_buffer(4872) := X"AC440014";
        ram_buffer(4873) := X"0060F809";
        ram_buffer(4874) := X"02402021";
        ram_buffer(4875) := X"93A30019";
        ram_buffer(4876) := X"93A40018";
        ram_buffer(4877) := X"93A2001A";
        ram_buffer(4878) := X"00031A00";
        ram_buffer(4879) := X"93B1001B";
        ram_buffer(4880) := X"00641821";
        ram_buffer(4881) := X"00021400";
        ram_buffer(4882) := X"00621021";
        ram_buffer(4883) := X"00118E00";
        ram_buffer(4884) := X"00518821";
        ram_buffer(4885) := X"2622FFF4";
        ram_buffer(4886) := X"2C420035";
        ram_buffer(4887) := X"104001DF";
        ram_buffer(4888) := X"240403EB";
        ram_buffer(4889) := X"2634FFFC";
        ram_buffer(4890) := X"8E07000C";
        ram_buffer(4891) := X"02803021";
        ram_buffer(4892) := X"24050001";
        ram_buffer(4893) := X"0C0272E9";
        ram_buffer(4894) := X"27A4001C";
        ram_buffer(4895) := X"12820008";
        ram_buffer(4896) := X"24020028";
        ram_buffer(4897) := X"8E420000";
        ram_buffer(4898) := X"2404002A";
        ram_buffer(4899) := X"8C430000";
        ram_buffer(4900) := X"AC440014";
        ram_buffer(4901) := X"0060F809";
        ram_buffer(4902) := X"02402021";
        ram_buffer(4903) := X"24020028";
        ram_buffer(4904) := X"12220099";
        ram_buffer(4905) := X"24020040";
        ram_buffer(4906) := X"12220097";
        ram_buffer(4907) := X"2402000C";
        ram_buffer(4908) := X"1222005A";
        ram_buffer(4909) := X"240403EB";
        ram_buffer(4910) := X"8E420000";
        ram_buffer(4911) := X"00000000";
        ram_buffer(4912) := X"8C430000";
        ram_buffer(4913) := X"02719823";
        ram_buffer(4914) := X"AC440014";
        ram_buffer(4915) := X"2673FFF2";
        ram_buffer(4916) := X"0060F809";
        ram_buffer(4917) := X"02402021";
        ram_buffer(4918) := X"0000A021";
        ram_buffer(4919) := X"0000A821";
        ram_buffer(4920) := X"066001C8";
        ram_buffer(4921) := X"0000F021";
        ram_buffer(4922) := X"2417FFFF";
        ram_buffer(4923) := X"2416002A";
        ram_buffer(4924) := X"2673FFFF";
        ram_buffer(4925) := X"0660000D";
        ram_buffer(4926) := X"00000000";
        ram_buffer(4927) := X"8E05000C";
        ram_buffer(4928) := X"00000000";
        ram_buffer(4929) := X"8CA20004";
        ram_buffer(4930) := X"00000000";
        ram_buffer(4931) := X"2442FFFF";
        ram_buffer(4932) := X"0440006E";
        ram_buffer(4933) := X"ACA20004";
        ram_buffer(4934) := X"8CA20000";
        ram_buffer(4935) := X"2673FFFF";
        ram_buffer(4936) := X"24420001";
        ram_buffer(4937) := X"0661FFF5";
        ram_buffer(4938) := X"ACA20000";
        ram_buffer(4939) := X"8E03002C";
        ram_buffer(4940) := X"24020018";
        ram_buffer(4941) := X"106201B1";
        ram_buffer(4942) := X"00000000";
        ram_buffer(4943) := X"10000001";
        ram_buffer(4944) := X"03C03821";
        ram_buffer(4945) := X"30E20003";
        ram_buffer(4946) := X"1440FFFE";
        ram_buffer(4947) := X"24E70001";
        ram_buffer(4948) := X"24E7FFFF";
        ram_buffer(4949) := X"8E420004";
        ram_buffer(4950) := X"24030001";
        ram_buffer(4951) := X"AFA30014";
        ram_buffer(4952) := X"AFB40010";
        ram_buffer(4953) := X"8C420010";
        ram_buffer(4954) := X"00003021";
        ram_buffer(4955) := X"AE070028";
        ram_buffer(4956) := X"24050001";
        ram_buffer(4957) := X"0040F809";
        ram_buffer(4958) := X"02402021";
        ram_buffer(4959) := X"8E430008";
        ram_buffer(4960) := X"AE020020";
        ram_buffer(4961) := X"3C021008";
        ram_buffer(4962) := X"24424954";
        ram_buffer(4963) := X"10600005";
        ram_buffer(4964) := X"AE020004";
        ram_buffer(4965) := X"8C620018";
        ram_buffer(4966) := X"00000000";
        ram_buffer(4967) := X"24420001";
        ram_buffer(4968) := X"AC620018";
        ram_buffer(4969) := X"8E420004";
        ram_buffer(4970) := X"02A03021";
        ram_buffer(4971) := X"8C420008";
        ram_buffer(4972) := X"02402021";
        ram_buffer(4973) := X"24070001";
        ram_buffer(4974) := X"0040F809";
        ram_buffer(4975) := X"24050001";
        ram_buffer(4976) := X"AE020010";
        ram_buffer(4977) := X"24020001";
        ram_buffer(4978) := X"AE020014";
        ram_buffer(4979) := X"24020002";
        ram_buffer(4980) := X"AE420024";
        ram_buffer(4981) := X"8FBF00A4";
        ram_buffer(4982) := X"24020003";
        ram_buffer(4983) := X"AE420020";
        ram_buffer(4984) := X"24020008";
        ram_buffer(4985) := X"AE5E0018";
        ram_buffer(4986) := X"AE54001C";
        ram_buffer(4987) := X"AE420030";
        ram_buffer(4988) := X"8FBE00A0";
        ram_buffer(4989) := X"8FB7009C";
        ram_buffer(4990) := X"8FB60098";
        ram_buffer(4991) := X"8FB50094";
        ram_buffer(4992) := X"8FB40090";
        ram_buffer(4993) := X"8FB3008C";
        ram_buffer(4994) := X"8FB20088";
        ram_buffer(4995) := X"8FB10084";
        ram_buffer(4996) := X"8FB00080";
        ram_buffer(4997) := X"03E00008";
        ram_buffer(4998) := X"27BD00A8";
        ram_buffer(4999) := X"93A5001F";
        ram_buffer(5000) := X"93A20023";
        ram_buffer(5001) := X"93A30021";
        ram_buffer(5002) := X"93A4001D";
        ram_buffer(5003) := X"93B4001E";
        ram_buffer(5004) := X"93A60022";
        ram_buffer(5005) := X"93B10020";
        ram_buffer(5006) := X"00031A00";
        ram_buffer(5007) := X"93BE001C";
        ram_buffer(5008) := X"00052A00";
        ram_buffer(5009) := X"00021200";
        ram_buffer(5010) := X"00042200";
        ram_buffer(5011) := X"00B4A021";
        ram_buffer(5012) := X"00461021";
        ram_buffer(5013) := X"00718821";
        ram_buffer(5014) := X"24030008";
        ram_buffer(5015) := X"009EF021";
        ram_buffer(5016) := X"0280B821";
        ram_buffer(5017) := X"104301A2";
        ram_buffer(5018) := X"AE02002C";
        ram_buffer(5019) := X"24030018";
        ram_buffer(5020) := X"1043017C";
        ram_buffer(5021) := X"24050001";
        ram_buffer(5022) := X"8E420000";
        ram_buffer(5023) := X"240403EA";
        ram_buffer(5024) := X"8C430000";
        ram_buffer(5025) := X"AC440014";
        ram_buffer(5026) := X"0060F809";
        ram_buffer(5027) := X"02402021";
        ram_buffer(5028) := X"24020001";
        ram_buffer(5029) := X"12220007";
        ram_buffer(5030) := X"00000000";
        ram_buffer(5031) := X"8E420000";
        ram_buffer(5032) := X"240403EC";
        ram_buffer(5033) := X"8C430000";
        ram_buffer(5034) := X"AC440014";
        ram_buffer(5035) := X"0060F809";
        ram_buffer(5036) := X"02402021";
        ram_buffer(5037) := X"001EA840";
        ram_buffer(5038) := X"2673FFE6";
        ram_buffer(5039) := X"0661FF8A";
        ram_buffer(5040) := X"02BEA821";
        ram_buffer(5041) := X"1000014F";
        ram_buffer(5042) := X"00000000";
        ram_buffer(5043) := X"8F848098";
        ram_buffer(5044) := X"0C028350";
        ram_buffer(5045) := X"00000000";
        ram_buffer(5046) := X"1457FF85";
        ram_buffer(5047) := X"00000000";
        ram_buffer(5048) := X"8E040018";
        ram_buffer(5049) := X"00000000";
        ram_buffer(5050) := X"8C820000";
        ram_buffer(5051) := X"00000000";
        ram_buffer(5052) := X"8C430000";
        ram_buffer(5053) := X"00000000";
        ram_buffer(5054) := X"0060F809";
        ram_buffer(5055) := X"AC560014";
        ram_buffer(5056) := X"1000FF7C";
        ram_buffer(5057) := X"2673FFFF";
        ram_buffer(5058) := X"93A2001E";
        ram_buffer(5059) := X"93AB001D";
        ram_buffer(5060) := X"AFA20068";
        ram_buffer(5061) := X"93A2003B";
        ram_buffer(5062) := X"93BE001C";
        ram_buffer(5063) := X"AFA2006C";
        ram_buffer(5064) := X"93A90029";
        ram_buffer(5065) := X"8FA20068";
        ram_buffer(5066) := X"93B60028";
        ram_buffer(5067) := X"93A30039";
        ram_buffer(5068) := X"93A6002A";
        ram_buffer(5069) := X"000B5A00";
        ram_buffer(5070) := X"93B40038";
        ram_buffer(5071) := X"93B8003A";
        ram_buffer(5072) := X"93AD002B";
        ram_buffer(5073) := X"017E5821";
        ram_buffer(5074) := X"00021400";
        ram_buffer(5075) := X"00094A00";
        ram_buffer(5076) := X"01625821";
        ram_buffer(5077) := X"00031A00";
        ram_buffer(5078) := X"8FA2006C";
        ram_buffer(5079) := X"01364821";
        ram_buffer(5080) := X"00063400";
        ram_buffer(5081) := X"00741821";
        ram_buffer(5082) := X"93A70027";
        ram_buffer(5083) := X"0018A400";
        ram_buffer(5084) := X"0126B021";
        ram_buffer(5085) := X"000D6E00";
        ram_buffer(5086) := X"93AA0021";
        ram_buffer(5087) := X"93BF0026";
        ram_buffer(5088) := X"0074A021";
        ram_buffer(5089) := X"00021E00";
        ram_buffer(5090) := X"02CD1021";
        ram_buffer(5091) := X"93B70020";
        ram_buffer(5092) := X"93A50022";
        ram_buffer(5093) := X"AFA20068";
        ram_buffer(5094) := X"00073A00";
        ram_buffer(5095) := X"93A20034";
        ram_buffer(5096) := X"000A5200";
        ram_buffer(5097) := X"00FF3821";
        ram_buffer(5098) := X"93B50030";
        ram_buffer(5099) := X"93A40031";
        ram_buffer(5100) := X"93B90032";
        ram_buffer(5101) := X"93AF001F";
        ram_buffer(5102) := X"93AE0023";
        ram_buffer(5103) := X"93A80025";
        ram_buffer(5104) := X"93AC0033";
        ram_buffer(5105) := X"01575021";
        ram_buffer(5106) := X"AE07002C";
        ram_buffer(5107) := X"0005BC00";
        ram_buffer(5108) := X"AFA2006C";
        ram_buffer(5109) := X"93A50024";
        ram_buffer(5110) := X"93A20035";
        ram_buffer(5111) := X"00042200";
        ram_buffer(5112) := X"AFA20070";
        ram_buffer(5113) := X"93A20036";
        ram_buffer(5114) := X"00952021";
        ram_buffer(5115) := X"AFA20074";
        ram_buffer(5116) := X"93A20037";
        ram_buffer(5117) := X"0019CC00";
        ram_buffer(5118) := X"000F7E00";
        ram_buffer(5119) := X"0157B821";
        ram_buffer(5120) := X"000E7600";
        ram_buffer(5121) := X"00084200";
        ram_buffer(5122) := X"0099A821";
        ram_buffer(5123) := X"000C6600";
        ram_buffer(5124) := X"AFA20078";
        ram_buffer(5125) := X"24020008";
        ram_buffer(5126) := X"016FF021";
        ram_buffer(5127) := X"02EEB821";
        ram_buffer(5128) := X"01054021";
        ram_buffer(5129) := X"02ACA821";
        ram_buffer(5130) := X"10E201D1";
        ram_buffer(5131) := X"0283A021";
        ram_buffer(5132) := X"24020018";
        ram_buffer(5133) := X"10E200FB";
        ram_buffer(5134) := X"240403F0";
        ram_buffer(5135) := X"8E420000";
        ram_buffer(5136) := X"240403EA";
        ram_buffer(5137) := X"8C430000";
        ram_buffer(5138) := X"AC440014";
        ram_buffer(5139) := X"02402021";
        ram_buffer(5140) := X"0060F809";
        ram_buffer(5141) := X"AFA8007C";
        ram_buffer(5142) := X"8FA8007C";
        ram_buffer(5143) := X"0000B021";
        ram_buffer(5144) := X"24020001";
        ram_buffer(5145) := X"11020007";
        ram_buffer(5146) := X"00000000";
        ram_buffer(5147) := X"8E420000";
        ram_buffer(5148) := X"240403EC";
        ram_buffer(5149) := X"8C450000";
        ram_buffer(5150) := X"AC440014";
        ram_buffer(5151) := X"00A0F809";
        ram_buffer(5152) := X"02402021";
        ram_buffer(5153) := X"8FA20068";
        ram_buffer(5154) := X"00000000";
        ram_buffer(5155) := X"14400103";
        ram_buffer(5156) := X"00000000";
        ram_buffer(5157) := X"1AA0001B";
        ram_buffer(5158) := X"00000000";
        ram_buffer(5159) := X"8FA20070";
        ram_buffer(5160) := X"8FA3006C";
        ram_buffer(5161) := X"00021200";
        ram_buffer(5162) := X"00431021";
        ram_buffer(5163) := X"8FA30074";
        ram_buffer(5164) := X"00000000";
        ram_buffer(5165) := X"00032400";
        ram_buffer(5166) := X"8FA30078";
        ram_buffer(5167) := X"00441021";
        ram_buffer(5168) := X"00032600";
        ram_buffer(5169) := X"00441021";
        ram_buffer(5170) := X"1840000E";
        ram_buffer(5171) := X"24040064";
        ram_buffer(5172) := X"14800002";
        ram_buffer(5173) := X"02A4001A";
        ram_buffer(5174) := X"0007000D";
        ram_buffer(5175) := X"24050002";
        ram_buffer(5176) := X"A24500CC";
        ram_buffer(5177) := X"0000A812";
        ram_buffer(5178) := X"A65500CE";
        ram_buffer(5179) := X"00000000";
        ram_buffer(5180) := X"14800002";
        ram_buffer(5181) := X"0044001A";
        ram_buffer(5182) := X"0007000D";
        ram_buffer(5183) := X"00001012";
        ram_buffer(5184) := X"A64200D0";
        ram_buffer(5185) := X"02719823";
        ram_buffer(5186) := X"12C001A9";
        ram_buffer(5187) := X"2673FFF2";
        ram_buffer(5188) := X"1A8001AD";
        ram_buffer(5189) := X"2A820101";
        ram_buffer(5190) := X"1040018A";
        ram_buffer(5191) := X"02D40018";
        ram_buffer(5192) := X"02803021";
        ram_buffer(5193) := X"00001012";
        ram_buffer(5194) := X"AFA20068";
        ram_buffer(5195) := X"8E420004";
        ram_buffer(5196) := X"02402021";
        ram_buffer(5197) := X"8C420008";
        ram_buffer(5198) := X"24070003";
        ram_buffer(5199) := X"0040F809";
        ram_buffer(5200) := X"24050001";
        ram_buffer(5201) := X"24040003";
        ram_buffer(5202) := X"12C4010A";
        ram_buffer(5203) := X"AE02001C";
        ram_buffer(5204) := X"12C000DA";
        ram_buffer(5205) := X"240503E9";
        ram_buffer(5206) := X"0000B021";
        ram_buffer(5207) := X"10000035";
        ram_buffer(5208) := X"2411002A";
        ram_buffer(5209) := X"8CA20000";
        ram_buffer(5210) := X"00000000";
        ram_buffer(5211) := X"24440001";
        ram_buffer(5212) := X"ACA40000";
        ram_buffer(5213) := X"90420000";
        ram_buffer(5214) := X"00000000";
        ram_buffer(5215) := X"A2A20000";
        ram_buffer(5216) := X"8E05000C";
        ram_buffer(5217) := X"8E04001C";
        ram_buffer(5218) := X"8CA20004";
        ram_buffer(5219) := X"8C860004";
        ram_buffer(5220) := X"2442FFFF";
        ram_buffer(5221) := X"00D6A821";
        ram_buffer(5222) := X"04400046";
        ram_buffer(5223) := X"ACA20004";
        ram_buffer(5224) := X"8CA20000";
        ram_buffer(5225) := X"00000000";
        ram_buffer(5226) := X"24440001";
        ram_buffer(5227) := X"ACA40000";
        ram_buffer(5228) := X"90420000";
        ram_buffer(5229) := X"00000000";
        ram_buffer(5230) := X"A2A20000";
        ram_buffer(5231) := X"8E05000C";
        ram_buffer(5232) := X"8E04001C";
        ram_buffer(5233) := X"8CA20004";
        ram_buffer(5234) := X"8C860000";
        ram_buffer(5235) := X"2442FFFF";
        ram_buffer(5236) := X"00D6A821";
        ram_buffer(5237) := X"04400050";
        ram_buffer(5238) := X"ACA20004";
        ram_buffer(5239) := X"8CA20000";
        ram_buffer(5240) := X"00000000";
        ram_buffer(5241) := X"24440001";
        ram_buffer(5242) := X"ACA40000";
        ram_buffer(5243) := X"90420000";
        ram_buffer(5244) := X"00000000";
        ram_buffer(5245) := X"A2A20000";
        ram_buffer(5246) := X"8E05000C";
        ram_buffer(5247) := X"00000000";
        ram_buffer(5248) := X"8CA20004";
        ram_buffer(5249) := X"00000000";
        ram_buffer(5250) := X"2442FFFF";
        ram_buffer(5251) := X"0440005A";
        ram_buffer(5252) := X"ACA20004";
        ram_buffer(5253) := X"8CA20000";
        ram_buffer(5254) := X"00000000";
        ram_buffer(5255) := X"24420001";
        ram_buffer(5256) := X"ACA20000";
        ram_buffer(5257) := X"26D60001";
        ram_buffer(5258) := X"12960063";
        ram_buffer(5259) := X"00000000";
        ram_buffer(5260) := X"8E02001C";
        ram_buffer(5261) := X"8E05000C";
        ram_buffer(5262) := X"8C460008";
        ram_buffer(5263) := X"8CA20004";
        ram_buffer(5264) := X"00D6A821";
        ram_buffer(5265) := X"2442FFFF";
        ram_buffer(5266) := X"0441FFC6";
        ram_buffer(5267) := X"ACA20004";
        ram_buffer(5268) := X"8F848098";
        ram_buffer(5269) := X"0C028350";
        ram_buffer(5270) := X"00000000";
        ram_buffer(5271) := X"2403FFFF";
        ram_buffer(5272) := X"1443FFC6";
        ram_buffer(5273) := X"00000000";
        ram_buffer(5274) := X"8E040018";
        ram_buffer(5275) := X"AFA2006C";
        ram_buffer(5276) := X"8C850000";
        ram_buffer(5277) := X"00000000";
        ram_buffer(5278) := X"8CA70000";
        ram_buffer(5279) := X"00000000";
        ram_buffer(5280) := X"00E0F809";
        ram_buffer(5281) := X"ACB10014";
        ram_buffer(5282) := X"8FA2006C";
        ram_buffer(5283) := X"00000000";
        ram_buffer(5284) := X"A2A20000";
        ram_buffer(5285) := X"8E05000C";
        ram_buffer(5286) := X"8E04001C";
        ram_buffer(5287) := X"8CA20004";
        ram_buffer(5288) := X"8C860004";
        ram_buffer(5289) := X"2442FFFF";
        ram_buffer(5290) := X"00D6A821";
        ram_buffer(5291) := X"0441FFBC";
        ram_buffer(5292) := X"ACA20004";
        ram_buffer(5293) := X"8F848098";
        ram_buffer(5294) := X"0C028350";
        ram_buffer(5295) := X"00000000";
        ram_buffer(5296) := X"2403FFFF";
        ram_buffer(5297) := X"1443FFBC";
        ram_buffer(5298) := X"00000000";
        ram_buffer(5299) := X"8E040018";
        ram_buffer(5300) := X"AFA2006C";
        ram_buffer(5301) := X"8C850000";
        ram_buffer(5302) := X"00000000";
        ram_buffer(5303) := X"8CA70000";
        ram_buffer(5304) := X"00000000";
        ram_buffer(5305) := X"00E0F809";
        ram_buffer(5306) := X"ACB10014";
        ram_buffer(5307) := X"8FA2006C";
        ram_buffer(5308) := X"00000000";
        ram_buffer(5309) := X"A2A20000";
        ram_buffer(5310) := X"8E05000C";
        ram_buffer(5311) := X"8E04001C";
        ram_buffer(5312) := X"8CA20004";
        ram_buffer(5313) := X"8C860000";
        ram_buffer(5314) := X"2442FFFF";
        ram_buffer(5315) := X"00D6A821";
        ram_buffer(5316) := X"0441FFB2";
        ram_buffer(5317) := X"ACA20004";
        ram_buffer(5318) := X"8F848098";
        ram_buffer(5319) := X"0C028350";
        ram_buffer(5320) := X"00000000";
        ram_buffer(5321) := X"2403FFFF";
        ram_buffer(5322) := X"1443FFB2";
        ram_buffer(5323) := X"00000000";
        ram_buffer(5324) := X"8E040018";
        ram_buffer(5325) := X"AFA2006C";
        ram_buffer(5326) := X"8C850000";
        ram_buffer(5327) := X"00000000";
        ram_buffer(5328) := X"8CA70000";
        ram_buffer(5329) := X"00000000";
        ram_buffer(5330) := X"00E0F809";
        ram_buffer(5331) := X"ACB10014";
        ram_buffer(5332) := X"8FA2006C";
        ram_buffer(5333) := X"00000000";
        ram_buffer(5334) := X"A2A20000";
        ram_buffer(5335) := X"8E05000C";
        ram_buffer(5336) := X"00000000";
        ram_buffer(5337) := X"8CA20004";
        ram_buffer(5338) := X"00000000";
        ram_buffer(5339) := X"2442FFFF";
        ram_buffer(5340) := X"0441FFA8";
        ram_buffer(5341) := X"ACA20004";
        ram_buffer(5342) := X"8F848098";
        ram_buffer(5343) := X"0C028350";
        ram_buffer(5344) := X"00000000";
        ram_buffer(5345) := X"2403FFFF";
        ram_buffer(5346) := X"1443FFA6";
        ram_buffer(5347) := X"00000000";
        ram_buffer(5348) := X"8E040018";
        ram_buffer(5349) := X"26D60001";
        ram_buffer(5350) := X"8C820000";
        ram_buffer(5351) := X"00000000";
        ram_buffer(5352) := X"8C450000";
        ram_buffer(5353) := X"00000000";
        ram_buffer(5354) := X"00A0F809";
        ram_buffer(5355) := X"AC510014";
        ram_buffer(5356) := X"1696FF9F";
        ram_buffer(5357) := X"00000000";
        ram_buffer(5358) := X"8FA20068";
        ram_buffer(5359) := X"001EA840";
        ram_buffer(5360) := X"02629823";
        ram_buffer(5361) := X"02E0A021";
        ram_buffer(5362) := X"02BEA821";
        ram_buffer(5363) := X"0661FE46";
        ram_buffer(5364) := X"00000000";
        ram_buffer(5365) := X"1000000B";
        ram_buffer(5366) := X"00000000";
        ram_buffer(5367) := X"8E420000";
        ram_buffer(5368) := X"00000000";
        ram_buffer(5369) := X"8C430000";
        ram_buffer(5370) := X"AC440014";
        ram_buffer(5371) := X"0060F809";
        ram_buffer(5372) := X"02402021";
        ram_buffer(5373) := X"1000FE1C";
        ram_buffer(5374) := X"2634FFFC";
        ram_buffer(5375) := X"1000FE51";
        ram_buffer(5376) := X"02A03821";
        ram_buffer(5377) := X"8E420000";
        ram_buffer(5378) := X"240403EB";
        ram_buffer(5379) := X"8C430000";
        ram_buffer(5380) := X"AC440014";
        ram_buffer(5381) := X"0060F809";
        ram_buffer(5382) := X"02402021";
        ram_buffer(5383) := X"1000FE33";
        ram_buffer(5384) := X"2417FFFF";
        ram_buffer(5385) := X"8E420000";
        ram_buffer(5386) := X"00000000";
        ram_buffer(5387) := X"AC5E0018";
        ram_buffer(5388) := X"8E430000";
        ram_buffer(5389) := X"AC440014";
        ram_buffer(5390) := X"AC77001C";
        ram_buffer(5391) := X"8E420000";
        ram_buffer(5392) := X"24050001";
        ram_buffer(5393) := X"8C420004";
        ram_buffer(5394) := X"02402021";
        ram_buffer(5395) := X"AFA8007C";
        ram_buffer(5396) := X"0040F809";
        ram_buffer(5397) := X"0000B021";
        ram_buffer(5398) := X"8FA8007C";
        ram_buffer(5399) := X"1000FF01";
        ram_buffer(5400) := X"24020001";
        ram_buffer(5401) := X"8E420000";
        ram_buffer(5402) := X"240403F2";
        ram_buffer(5403) := X"AC5E0018";
        ram_buffer(5404) := X"8E430000";
        ram_buffer(5405) := X"AC440014";
        ram_buffer(5406) := X"AC74001C";
        ram_buffer(5407) := X"8E420000";
        ram_buffer(5408) := X"00000000";
        ram_buffer(5409) := X"8C420004";
        ram_buffer(5410) := X"00000000";
        ram_buffer(5411) := X"0040F809";
        ram_buffer(5412) := X"02402021";
        ram_buffer(5413) := X"1000FE7F";
        ram_buffer(5414) := X"24020001";
        ram_buffer(5415) := X"8E420000";
        ram_buffer(5416) := X"240403EE";
        ram_buffer(5417) := X"8C450000";
        ram_buffer(5418) := X"AC440014";
        ram_buffer(5419) := X"00A0F809";
        ram_buffer(5420) := X"02402021";
        ram_buffer(5421) := X"1000FEF7";
        ram_buffer(5422) := X"00000000";
        ram_buffer(5423) := X"8E040018";
        ram_buffer(5424) := X"00000000";
        ram_buffer(5425) := X"8C820000";
        ram_buffer(5426) := X"001EA840";
        ram_buffer(5427) := X"8C430000";
        ram_buffer(5428) := X"00000000";
        ram_buffer(5429) := X"0060F809";
        ram_buffer(5430) := X"AC450014";
        ram_buffer(5431) := X"8FA20068";
        ram_buffer(5432) := X"02E0A021";
        ram_buffer(5433) := X"02629823";
        ram_buffer(5434) := X"1000FFB8";
        ram_buffer(5435) := X"02BEA821";
        ram_buffer(5436) := X"8E420000";
        ram_buffer(5437) := X"240403F3";
        ram_buffer(5438) := X"AC5E0018";
        ram_buffer(5439) := X"8E430000";
        ram_buffer(5440) := X"AC440014";
        ram_buffer(5441) := X"AC74001C";
        ram_buffer(5442) := X"8E420000";
        ram_buffer(5443) := X"24050001";
        ram_buffer(5444) := X"8C420004";
        ram_buffer(5445) := X"00000000";
        ram_buffer(5446) := X"0040F809";
        ram_buffer(5447) := X"02402021";
        ram_buffer(5448) := X"24020001";
        ram_buffer(5449) := X"12220007";
        ram_buffer(5450) := X"240503EC";
        ram_buffer(5451) := X"8E420000";
        ram_buffer(5452) := X"00000000";
        ram_buffer(5453) := X"8C430000";
        ram_buffer(5454) := X"02402021";
        ram_buffer(5455) := X"0060F809";
        ram_buffer(5456) := X"AC450014";
        ram_buffer(5457) := X"8E420004";
        ram_buffer(5458) := X"24070003";
        ram_buffer(5459) := X"8C420008";
        ram_buffer(5460) := X"24060100";
        ram_buffer(5461) := X"24050001";
        ram_buffer(5462) := X"0040F809";
        ram_buffer(5463) := X"02402021";
        ram_buffer(5464) := X"24030300";
        ram_buffer(5465) := X"2673FFE6";
        ram_buffer(5466) := X"AE02001C";
        ram_buffer(5467) := X"AFA30068";
        ram_buffer(5468) := X"24140100";
        ram_buffer(5469) := X"0000A821";
        ram_buffer(5470) := X"10000028";
        ram_buffer(5471) := X"2411002A";
        ram_buffer(5472) := X"8CA20000";
        ram_buffer(5473) := X"00000000";
        ram_buffer(5474) := X"24440001";
        ram_buffer(5475) := X"ACA40000";
        ram_buffer(5476) := X"90420000";
        ram_buffer(5477) := X"00000000";
        ram_buffer(5478) := X"A2C20000";
        ram_buffer(5479) := X"8E05000C";
        ram_buffer(5480) := X"8E04001C";
        ram_buffer(5481) := X"8CA20004";
        ram_buffer(5482) := X"8C860004";
        ram_buffer(5483) := X"2442FFFF";
        ram_buffer(5484) := X"00D5B021";
        ram_buffer(5485) := X"04400039";
        ram_buffer(5486) := X"ACA20004";
        ram_buffer(5487) := X"8CA20000";
        ram_buffer(5488) := X"00000000";
        ram_buffer(5489) := X"24440001";
        ram_buffer(5490) := X"ACA40000";
        ram_buffer(5491) := X"90420000";
        ram_buffer(5492) := X"00000000";
        ram_buffer(5493) := X"A2C20000";
        ram_buffer(5494) := X"8E05000C";
        ram_buffer(5495) := X"8E04001C";
        ram_buffer(5496) := X"8CA20004";
        ram_buffer(5497) := X"8C860000";
        ram_buffer(5498) := X"2442FFFF";
        ram_buffer(5499) := X"00D5B021";
        ram_buffer(5500) := X"04400043";
        ram_buffer(5501) := X"ACA20004";
        ram_buffer(5502) := X"8CA20000";
        ram_buffer(5503) := X"00000000";
        ram_buffer(5504) := X"24440001";
        ram_buffer(5505) := X"ACA40000";
        ram_buffer(5506) := X"90420000";
        ram_buffer(5507) := X"26B50001";
        ram_buffer(5508) := X"12B4FF69";
        ram_buffer(5509) := X"A2C20000";
        ram_buffer(5510) := X"8E02001C";
        ram_buffer(5511) := X"8E05000C";
        ram_buffer(5512) := X"8C460008";
        ram_buffer(5513) := X"8CA20004";
        ram_buffer(5514) := X"00D5B021";
        ram_buffer(5515) := X"2442FFFF";
        ram_buffer(5516) := X"0441FFD3";
        ram_buffer(5517) := X"ACA20004";
        ram_buffer(5518) := X"8F848098";
        ram_buffer(5519) := X"0C028350";
        ram_buffer(5520) := X"00000000";
        ram_buffer(5521) := X"2403FFFF";
        ram_buffer(5522) := X"1443FFD3";
        ram_buffer(5523) := X"00000000";
        ram_buffer(5524) := X"8E040018";
        ram_buffer(5525) := X"AFA2006C";
        ram_buffer(5526) := X"8C850000";
        ram_buffer(5527) := X"00000000";
        ram_buffer(5528) := X"8CA70000";
        ram_buffer(5529) := X"00000000";
        ram_buffer(5530) := X"00E0F809";
        ram_buffer(5531) := X"ACB10014";
        ram_buffer(5532) := X"8FA2006C";
        ram_buffer(5533) := X"00000000";
        ram_buffer(5534) := X"A2C20000";
        ram_buffer(5535) := X"8E05000C";
        ram_buffer(5536) := X"8E04001C";
        ram_buffer(5537) := X"8CA20004";
        ram_buffer(5538) := X"8C860004";
        ram_buffer(5539) := X"2442FFFF";
        ram_buffer(5540) := X"00D5B021";
        ram_buffer(5541) := X"0441FFC9";
        ram_buffer(5542) := X"ACA20004";
        ram_buffer(5543) := X"8F848098";
        ram_buffer(5544) := X"0C028350";
        ram_buffer(5545) := X"00000000";
        ram_buffer(5546) := X"2403FFFF";
        ram_buffer(5547) := X"1443FFC9";
        ram_buffer(5548) := X"00000000";
        ram_buffer(5549) := X"8E040018";
        ram_buffer(5550) := X"AFA2006C";
        ram_buffer(5551) := X"8C850000";
        ram_buffer(5552) := X"00000000";
        ram_buffer(5553) := X"8CA70000";
        ram_buffer(5554) := X"00000000";
        ram_buffer(5555) := X"00E0F809";
        ram_buffer(5556) := X"ACB10014";
        ram_buffer(5557) := X"8FA2006C";
        ram_buffer(5558) := X"00000000";
        ram_buffer(5559) := X"A2C20000";
        ram_buffer(5560) := X"8E05000C";
        ram_buffer(5561) := X"8E04001C";
        ram_buffer(5562) := X"8CA20004";
        ram_buffer(5563) := X"8C860000";
        ram_buffer(5564) := X"2442FFFF";
        ram_buffer(5565) := X"00D5B021";
        ram_buffer(5566) := X"0441FFBF";
        ram_buffer(5567) := X"ACA20004";
        ram_buffer(5568) := X"8F848098";
        ram_buffer(5569) := X"0C028350";
        ram_buffer(5570) := X"00000000";
        ram_buffer(5571) := X"2403FFFF";
        ram_buffer(5572) := X"1443FFBE";
        ram_buffer(5573) := X"00000000";
        ram_buffer(5574) := X"8E040018";
        ram_buffer(5575) := X"AFA2006C";
        ram_buffer(5576) := X"8C850000";
        ram_buffer(5577) := X"00000000";
        ram_buffer(5578) := X"8CA70000";
        ram_buffer(5579) := X"00000000";
        ram_buffer(5580) := X"00E0F809";
        ram_buffer(5581) := X"ACB10014";
        ram_buffer(5582) := X"8FA2006C";
        ram_buffer(5583) := X"1000FFB4";
        ram_buffer(5584) := X"26B50001";
        ram_buffer(5585) := X"8E420000";
        ram_buffer(5586) := X"240403E9";
        ram_buffer(5587) := X"8C450000";
        ram_buffer(5588) := X"AC440014";
        ram_buffer(5589) := X"00A0F809";
        ram_buffer(5590) := X"02402021";
        ram_buffer(5591) := X"02D40018";
        ram_buffer(5592) := X"02803021";
        ram_buffer(5593) := X"00001012";
        ram_buffer(5594) := X"1000FE70";
        ram_buffer(5595) := X"AFA20068";
        ram_buffer(5596) := X"8E420000";
        ram_buffer(5597) := X"240403F1";
        ram_buffer(5598) := X"AC5E0018";
        ram_buffer(5599) := X"8E430000";
        ram_buffer(5600) := X"AC440014";
        ram_buffer(5601) := X"AC77001C";
        ram_buffer(5602) := X"8E420000";
        ram_buffer(5603) := X"24050001";
        ram_buffer(5604) := X"8C420004";
        ram_buffer(5605) := X"02402021";
        ram_buffer(5606) := X"AFA8007C";
        ram_buffer(5607) := X"0040F809";
        ram_buffer(5608) := X"24160004";
        ram_buffer(5609) := X"8FA8007C";
        ram_buffer(5610) := X"1000FE2E";
        ram_buffer(5611) := X"24020001";
        ram_buffer(5612) := X"001EA840";
        ram_buffer(5613) := X"02E0A021";
        ram_buffer(5614) := X"0661FD4B";
        ram_buffer(5615) := X"02BEA821";
        ram_buffer(5616) := X"1000FF10";
        ram_buffer(5617) := X"00000000";
        ram_buffer(5618) := X"00161200";
        ram_buffer(5619) := X"AFA20068";
        ram_buffer(5620) := X"24060100";
        ram_buffer(5621) := X"1000FE55";
        ram_buffer(5622) := X"24140100";
        ram_buffer(5623) := X"8C820004";
        ram_buffer(5624) := X"27BDFFE8";
        ram_buffer(5625) := X"8C420000";
        ram_buffer(5626) := X"24060030";
        ram_buffer(5627) := X"AFBF0014";
        ram_buffer(5628) := X"AFB00010";
        ram_buffer(5629) := X"24050001";
        ram_buffer(5630) := X"0040F809";
        ram_buffer(5631) := X"00808021";
        ram_buffer(5632) := X"3C041008";
        ram_buffer(5633) := X"24844B2C";
        ram_buffer(5634) := X"AC440000";
        ram_buffer(5635) := X"8FBF0014";
        ram_buffer(5636) := X"3C041008";
        ram_buffer(5637) := X"2484494C";
        ram_buffer(5638) := X"AC500018";
        ram_buffer(5639) := X"AC440008";
        ram_buffer(5640) := X"8FB00010";
        ram_buffer(5641) := X"03E00008";
        ram_buffer(5642) := X"27BD0018";
        ram_buffer(5643) := X"27BDFFD0";
        ram_buffer(5644) := X"AFB50024";
        ram_buffer(5645) := X"AFB40020";
        ram_buffer(5646) := X"AFB3001C";
        ram_buffer(5647) := X"AFB20018";
        ram_buffer(5648) := X"AFB10014";
        ram_buffer(5649) := X"AFB00010";
        ram_buffer(5650) := X"AFBF002C";
        ram_buffer(5651) := X"AFB60028";
        ram_buffer(5652) := X"00808021";
        ram_buffer(5653) := X"00A09821";
        ram_buffer(5654) := X"00C09021";
        ram_buffer(5655) := X"2415000A";
        ram_buffer(5656) := X"2414FFFF";
        ram_buffer(5657) := X"24110023";
        ram_buffer(5658) := X"8E020004";
        ram_buffer(5659) := X"00000000";
        ram_buffer(5660) := X"2442FFFF";
        ram_buffer(5661) := X"04400053";
        ram_buffer(5662) := X"AE020004";
        ram_buffer(5663) := X"8E030000";
        ram_buffer(5664) := X"00000000";
        ram_buffer(5665) := X"24640001";
        ram_buffer(5666) := X"AE040000";
        ram_buffer(5667) := X"90630000";
        ram_buffer(5668) := X"00000000";
        ram_buffer(5669) := X"1071003F";
        ram_buffer(5670) := X"2442FFFF";
        ram_buffer(5671) := X"24620001";
        ram_buffer(5672) := X"8F848090";
        ram_buffer(5673) := X"00000000";
        ram_buffer(5674) := X"00821021";
        ram_buffer(5675) := X"90420000";
        ram_buffer(5676) := X"00000000";
        ram_buffer(5677) := X"30450008";
        ram_buffer(5678) := X"14A0FFEB";
        ram_buffer(5679) := X"30420004";
        ram_buffer(5680) := X"10400075";
        ram_buffer(5681) := X"2471FFD0";
        ram_buffer(5682) := X"8E020004";
        ram_buffer(5683) := X"00000000";
        ram_buffer(5684) := X"2442FFFF";
        ram_buffer(5685) := X"2416000A";
        ram_buffer(5686) := X"2415FFFF";
        ram_buffer(5687) := X"24140023";
        ram_buffer(5688) := X"04400019";
        ram_buffer(5689) := X"AE020004";
        ram_buffer(5690) := X"8E030000";
        ram_buffer(5691) := X"00000000";
        ram_buffer(5692) := X"24650001";
        ram_buffer(5693) := X"AE050000";
        ram_buffer(5694) := X"90650000";
        ram_buffer(5695) := X"00000000";
        ram_buffer(5696) := X"10B40050";
        ram_buffer(5697) := X"2442FFFF";
        ram_buffer(5698) := X"24A20001";
        ram_buffer(5699) := X"00821021";
        ram_buffer(5700) := X"90420000";
        ram_buffer(5701) := X"00000000";
        ram_buffer(5702) := X"30420004";
        ram_buffer(5703) := X"10400056";
        ram_buffer(5704) := X"00000000";
        ram_buffer(5705) := X"00111040";
        ram_buffer(5706) := X"001118C0";
        ram_buffer(5707) := X"00431821";
        ram_buffer(5708) := X"8E020004";
        ram_buffer(5709) := X"24A5FFD0";
        ram_buffer(5710) := X"2442FFFF";
        ram_buffer(5711) := X"00A38821";
        ram_buffer(5712) := X"0441FFE9";
        ram_buffer(5713) := X"AE020004";
        ram_buffer(5714) := X"8F848098";
        ram_buffer(5715) := X"0C028350";
        ram_buffer(5716) := X"02002821";
        ram_buffer(5717) := X"10540044";
        ram_buffer(5718) := X"00402821";
        ram_buffer(5719) := X"10550045";
        ram_buffer(5720) := X"00000000";
        ram_buffer(5721) := X"8F848090";
        ram_buffer(5722) := X"1000FFE8";
        ram_buffer(5723) := X"24A20001";
        ram_buffer(5724) := X"8E030000";
        ram_buffer(5725) := X"00000000";
        ram_buffer(5726) := X"24640001";
        ram_buffer(5727) := X"AE040000";
        ram_buffer(5728) := X"90630000";
        ram_buffer(5729) := X"00000000";
        ram_buffer(5730) := X"10750022";
        ram_buffer(5731) := X"00000000";
        ram_buffer(5732) := X"2442FFFF";
        ram_buffer(5733) := X"0441FFF6";
        ram_buffer(5734) := X"AE020004";
        ram_buffer(5735) := X"8F848098";
        ram_buffer(5736) := X"0C028350";
        ram_buffer(5737) := X"02002821";
        ram_buffer(5738) := X"1055001A";
        ram_buffer(5739) := X"00000000";
        ram_buffer(5740) := X"1054000B";
        ram_buffer(5741) := X"00000000";
        ram_buffer(5742) := X"8E020004";
        ram_buffer(5743) := X"1000FFF5";
        ram_buffer(5744) := X"2442FFFF";
        ram_buffer(5745) := X"8F848098";
        ram_buffer(5746) := X"0C028350";
        ram_buffer(5747) := X"02002821";
        ram_buffer(5748) := X"1051FFF9";
        ram_buffer(5749) := X"00401821";
        ram_buffer(5750) := X"1454FFB1";
        ram_buffer(5751) := X"24620001";
        ram_buffer(5752) := X"2402FFFF";
        ram_buffer(5753) := X"AE420000";
        ram_buffer(5754) := X"00001021";
        ram_buffer(5755) := X"8FBF002C";
        ram_buffer(5756) := X"8FB60028";
        ram_buffer(5757) := X"8FB50024";
        ram_buffer(5758) := X"8FB40020";
        ram_buffer(5759) := X"8FB3001C";
        ram_buffer(5760) := X"8FB20018";
        ram_buffer(5761) := X"8FB10014";
        ram_buffer(5762) := X"8FB00010";
        ram_buffer(5763) := X"03E00008";
        ram_buffer(5764) := X"27BD0030";
        ram_buffer(5765) := X"2402000B";
        ram_buffer(5766) := X"1000FFA1";
        ram_buffer(5767) := X"2403000A";
        ram_buffer(5768) := X"8E030000";
        ram_buffer(5769) := X"00000000";
        ram_buffer(5770) := X"24640001";
        ram_buffer(5771) := X"AE040000";
        ram_buffer(5772) := X"90630000";
        ram_buffer(5773) := X"00000000";
        ram_buffer(5774) := X"10760013";
        ram_buffer(5775) := X"00000000";
        ram_buffer(5776) := X"2442FFFF";
        ram_buffer(5777) := X"0441FFF6";
        ram_buffer(5778) := X"AE020004";
        ram_buffer(5779) := X"8F848098";
        ram_buffer(5780) := X"0C028350";
        ram_buffer(5781) := X"02002821";
        ram_buffer(5782) := X"1056000B";
        ram_buffer(5783) := X"00000000";
        ram_buffer(5784) := X"10550004";
        ram_buffer(5785) := X"00000000";
        ram_buffer(5786) := X"8E020004";
        ram_buffer(5787) := X"1000FFF5";
        ram_buffer(5788) := X"2442FFFF";
        ram_buffer(5789) := X"2405FFFF";
        ram_buffer(5790) := X"AE710000";
        ram_buffer(5791) := X"24020001";
        ram_buffer(5792) := X"1000FFDA";
        ram_buffer(5793) := X"AE450000";
        ram_buffer(5794) := X"2402000B";
        ram_buffer(5795) := X"8F848090";
        ram_buffer(5796) := X"1000FF9E";
        ram_buffer(5797) := X"2405000A";
        ram_buffer(5798) := X"1000FFD4";
        ram_buffer(5799) := X"AE430000";
        ram_buffer(5800) := X"27BDFFD8";
        ram_buffer(5801) := X"8CA20000";
        ram_buffer(5802) := X"AFB40020";
        ram_buffer(5803) := X"AFB3001C";
        ram_buffer(5804) := X"AFB20018";
        ram_buffer(5805) := X"AFB10014";
        ram_buffer(5806) := X"AFB00010";
        ram_buffer(5807) := X"AFBF0024";
        ram_buffer(5808) := X"00A09821";
        ram_buffer(5809) := X"00808021";
        ram_buffer(5810) := X"2411FFFF";
        ram_buffer(5811) := X"24120023";
        ram_buffer(5812) := X"2414000A";
        ram_buffer(5813) := X"10510030";
        ram_buffer(5814) := X"00000000";
        ram_buffer(5815) := X"8F858090";
        ram_buffer(5816) := X"00000000";
        ram_buffer(5817) := X"00A21821";
        ram_buffer(5818) := X"90630001";
        ram_buffer(5819) := X"00000000";
        ram_buffer(5820) := X"30640008";
        ram_buffer(5821) := X"10800048";
        ram_buffer(5822) := X"30630004";
        ram_buffer(5823) := X"8E030004";
        ram_buffer(5824) := X"00000000";
        ram_buffer(5825) := X"2463FFFF";
        ram_buffer(5826) := X"0460003B";
        ram_buffer(5827) := X"AE030004";
        ram_buffer(5828) := X"8E020000";
        ram_buffer(5829) := X"00000000";
        ram_buffer(5830) := X"24440001";
        ram_buffer(5831) := X"AE040000";
        ram_buffer(5832) := X"90420000";
        ram_buffer(5833) := X"00000000";
        ram_buffer(5834) := X"1452FFEE";
        ram_buffer(5835) := X"00000000";
        ram_buffer(5836) := X"10000009";
        ram_buffer(5837) := X"00601021";
        ram_buffer(5838) := X"8E030000";
        ram_buffer(5839) := X"00000000";
        ram_buffer(5840) := X"24640001";
        ram_buffer(5841) := X"AE040000";
        ram_buffer(5842) := X"90630000";
        ram_buffer(5843) := X"00000000";
        ram_buffer(5844) := X"1074000E";
        ram_buffer(5845) := X"00000000";
        ram_buffer(5846) := X"2442FFFF";
        ram_buffer(5847) := X"0441FFF6";
        ram_buffer(5848) := X"AE020004";
        ram_buffer(5849) := X"8F848098";
        ram_buffer(5850) := X"0C028350";
        ram_buffer(5851) := X"02002821";
        ram_buffer(5852) := X"10540006";
        ram_buffer(5853) := X"00000000";
        ram_buffer(5854) := X"1051FFD6";
        ram_buffer(5855) := X"00000000";
        ram_buffer(5856) := X"8E020004";
        ram_buffer(5857) := X"1000FFF5";
        ram_buffer(5858) := X"2442FFFF";
        ram_buffer(5859) := X"2402000A";
        ram_buffer(5860) := X"1451FFD2";
        ram_buffer(5861) := X"00000000";
        ram_buffer(5862) := X"8F828090";
        ram_buffer(5863) := X"00000000";
        ram_buffer(5864) := X"90420000";
        ram_buffer(5865) := X"00000000";
        ram_buffer(5866) := X"30420004";
        ram_buffer(5867) := X"10400008";
        ram_buffer(5868) := X"2402FFFF";
        ram_buffer(5869) := X"02002821";
        ram_buffer(5870) := X"0C029D83";
        ram_buffer(5871) := X"00402021";
        ram_buffer(5872) := X"2403FFFF";
        ram_buffer(5873) := X"10430004";
        ram_buffer(5874) := X"00001021";
        ram_buffer(5875) := X"24020020";
        ram_buffer(5876) := X"AE620000";
        ram_buffer(5877) := X"24020001";
        ram_buffer(5878) := X"8FBF0024";
        ram_buffer(5879) := X"8FB40020";
        ram_buffer(5880) := X"8FB3001C";
        ram_buffer(5881) := X"8FB20018";
        ram_buffer(5882) := X"8FB10014";
        ram_buffer(5883) := X"8FB00010";
        ram_buffer(5884) := X"03E00008";
        ram_buffer(5885) := X"27BD0028";
        ram_buffer(5886) := X"8F848098";
        ram_buffer(5887) := X"0C028350";
        ram_buffer(5888) := X"02002821";
        ram_buffer(5889) := X"1452FFB3";
        ram_buffer(5890) := X"00000000";
        ram_buffer(5891) := X"8E030004";
        ram_buffer(5892) := X"1000FFD1";
        ram_buffer(5893) := X"00601021";
        ram_buffer(5894) := X"1460FFE6";
        ram_buffer(5895) := X"2403003B";
        ram_buffer(5896) := X"1043FFEB";
        ram_buffer(5897) := X"2403003A";
        ram_buffer(5898) := X"1043FFE9";
        ram_buffer(5899) := X"00000000";
        ram_buffer(5900) := X"1000FFE7";
        ram_buffer(5901) := X"24020020";
        ram_buffer(5902) := X"27BDFEB8";
        ram_buffer(5903) := X"AFB3012C";
        ram_buffer(5904) := X"00A09821";
        ram_buffer(5905) := X"3C05100D";
        ram_buffer(5906) := X"AFA40148";
        ram_buffer(5907) := X"24A58F90";
        ram_buffer(5908) := X"02602021";
        ram_buffer(5909) := X"AFBE0140";
        ram_buffer(5910) := X"AFB7013C";
        ram_buffer(5911) := X"AFBF0144";
        ram_buffer(5912) := X"AFB60138";
        ram_buffer(5913) := X"AFB50134";
        ram_buffer(5914) := X"AFB40130";
        ram_buffer(5915) := X"AFB20128";
        ram_buffer(5916) := X"AFB10124";
        ram_buffer(5917) := X"AFB00120";
        ram_buffer(5918) := X"00C0B821";
        ram_buffer(5919) := X"0C02716A";
        ram_buffer(5920) := X"00E0F021";
        ram_buffer(5921) := X"10400040";
        ram_buffer(5922) := X"00409021";
        ram_buffer(5923) := X"0000A021";
        ram_buffer(5924) := X"27B60118";
        ram_buffer(5925) := X"24150004";
        ram_buffer(5926) := X"27A6011C";
        ram_buffer(5927) := X"02C02821";
        ram_buffer(5928) := X"0C02160B";
        ram_buffer(5929) := X"02402021";
        ram_buffer(5930) := X"1040003F";
        ram_buffer(5931) := X"00408821";
        ram_buffer(5932) := X"1295002B";
        ram_buffer(5933) := X"27B0001C";
        ram_buffer(5934) := X"8FA20118";
        ram_buffer(5935) := X"10000005";
        ram_buffer(5936) := X"AFA20018";
        ram_buffer(5937) := X"8FA20118";
        ram_buffer(5938) := X"26100004";
        ram_buffer(5939) := X"12D0001C";
        ram_buffer(5940) := X"AE02FFFC";
        ram_buffer(5941) := X"27A6011C";
        ram_buffer(5942) := X"02C02821";
        ram_buffer(5943) := X"0C02160B";
        ram_buffer(5944) := X"02402021";
        ram_buffer(5945) := X"1440FFF7";
        ram_buffer(5946) := X"00408821";
        ram_buffer(5947) := X"8F828098";
        ram_buffer(5948) := X"3C05100D";
        ram_buffer(5949) := X"8C44000C";
        ram_buffer(5950) := X"02603021";
        ram_buffer(5951) := X"0C027196";
        ram_buffer(5952) := X"24A58340";
        ram_buffer(5953) := X"0C026DBB";
        ram_buffer(5954) := X"02402021";
        ram_buffer(5955) := X"8FBF0144";
        ram_buffer(5956) := X"02201021";
        ram_buffer(5957) := X"8FBE0140";
        ram_buffer(5958) := X"8FB7013C";
        ram_buffer(5959) := X"8FB60138";
        ram_buffer(5960) := X"8FB50134";
        ram_buffer(5961) := X"8FB40130";
        ram_buffer(5962) := X"8FB3012C";
        ram_buffer(5963) := X"8FB20128";
        ram_buffer(5964) := X"8FB10124";
        ram_buffer(5965) := X"8FB00120";
        ram_buffer(5966) := X"03E00008";
        ram_buffer(5967) := X"27BD0148";
        ram_buffer(5968) := X"8FA40148";
        ram_buffer(5969) := X"02802821";
        ram_buffer(5970) := X"AFBE0010";
        ram_buffer(5971) := X"02E03821";
        ram_buffer(5972) := X"0C021B8E";
        ram_buffer(5973) := X"27A60018";
        ram_buffer(5974) := X"1000FFCF";
        ram_buffer(5975) := X"26940001";
        ram_buffer(5976) := X"8F828098";
        ram_buffer(5977) := X"3C05100D";
        ram_buffer(5978) := X"8C44000C";
        ram_buffer(5979) := X"02603021";
        ram_buffer(5980) := X"0C027196";
        ram_buffer(5981) := X"24A58324";
        ram_buffer(5982) := X"0C026DBB";
        ram_buffer(5983) := X"02402021";
        ram_buffer(5984) := X"1000FFE2";
        ram_buffer(5985) := X"00008821";
        ram_buffer(5986) := X"8F828098";
        ram_buffer(5987) := X"3C05100D";
        ram_buffer(5988) := X"8C44000C";
        ram_buffer(5989) := X"02603021";
        ram_buffer(5990) := X"0C027196";
        ram_buffer(5991) := X"24A58308";
        ram_buffer(5992) := X"1000FFDA";
        ram_buffer(5993) := X"00008821";
        ram_buffer(5994) := X"8FA3011C";
        ram_buffer(5995) := X"2402FFFF";
        ram_buffer(5996) := X"1062000B";
        ram_buffer(5997) := X"3C05100D";
        ram_buffer(5998) := X"8F828098";
        ram_buffer(5999) := X"00000000";
        ram_buffer(6000) := X"8C44000C";
        ram_buffer(6001) := X"02603021";
        ram_buffer(6002) := X"0C027196";
        ram_buffer(6003) := X"24A58360";
        ram_buffer(6004) := X"0C026DBB";
        ram_buffer(6005) := X"02402021";
        ram_buffer(6006) := X"1000FFCC";
        ram_buffer(6007) := X"00000000";
        ram_buffer(6008) := X"0C026DBB";
        ram_buffer(6009) := X"02402021";
        ram_buffer(6010) := X"1000FFC8";
        ram_buffer(6011) := X"24110001";
        ram_buffer(6012) := X"27BDF1B0";
        ram_buffer(6013) := X"AFB20E30";
        ram_buffer(6014) := X"00A09021";
        ram_buffer(6015) := X"3C05100D";
        ram_buffer(6016) := X"AFA40E50";
        ram_buffer(6017) := X"24A58F90";
        ram_buffer(6018) := X"02402021";
        ram_buffer(6019) := X"AFBF0E4C";
        ram_buffer(6020) := X"AFBE0E48";
        ram_buffer(6021) := X"AFB70E44";
        ram_buffer(6022) := X"AFB60E40";
        ram_buffer(6023) := X"AFB50E3C";
        ram_buffer(6024) := X"AFB40E38";
        ram_buffer(6025) := X"AFB30E34";
        ram_buffer(6026) := X"AFB10E2C";
        ram_buffer(6027) := X"0C02716A";
        ram_buffer(6028) := X"AFB00E28";
        ram_buffer(6029) := X"10400077";
        ram_buffer(6030) := X"00408021";
        ram_buffer(6031) := X"27B30018";
        ram_buffer(6032) := X"0000A821";
        ram_buffer(6033) := X"24160064";
        ram_buffer(6034) := X"24110020";
        ram_buffer(6035) := X"24140004";
        ram_buffer(6036) := X"27A60E24";
        ram_buffer(6037) := X"27A50E20";
        ram_buffer(6038) := X"0C02160B";
        ram_buffer(6039) := X"02002021";
        ram_buffer(6040) := X"1040004C";
        ram_buffer(6041) := X"27A50E24";
        ram_buffer(6042) := X"0C0216A8";
        ram_buffer(6043) := X"02002021";
        ram_buffer(6044) := X"10400048";
        ram_buffer(6045) := X"00000000";
        ram_buffer(6046) := X"12B600AD";
        ram_buffer(6047) := X"3C05100D";
        ram_buffer(6048) := X"8FA30E20";
        ram_buffer(6049) := X"8FA20E24";
        ram_buffer(6050) := X"AE63FFFC";
        ram_buffer(6051) := X"1451002A";
        ram_buffer(6052) := X"241E0001";
        ram_buffer(6053) := X"0260B821";
        ram_buffer(6054) := X"241E0001";
        ram_buffer(6055) := X"27A50E20";
        ram_buffer(6056) := X"02002021";
        ram_buffer(6057) := X"0C02160B";
        ram_buffer(6058) := X"27A60E24";
        ram_buffer(6059) := X"27A50E24";
        ram_buffer(6060) := X"1040002E";
        ram_buffer(6061) := X"02002021";
        ram_buffer(6062) := X"0C0216A8";
        ram_buffer(6063) := X"00000000";
        ram_buffer(6064) := X"1040002A";
        ram_buffer(6065) := X"00000000";
        ram_buffer(6066) := X"8FA40E20";
        ram_buffer(6067) := X"8FA20E24";
        ram_buffer(6068) := X"AEE40000";
        ram_buffer(6069) := X"14510018";
        ram_buffer(6070) := X"27DE0001";
        ram_buffer(6071) := X"17D4FFEF";
        ram_buffer(6072) := X"26F70004";
        ram_buffer(6073) := X"8F828098";
        ram_buffer(6074) := X"3C05100D";
        ram_buffer(6075) := X"8C44000C";
        ram_buffer(6076) := X"02403021";
        ram_buffer(6077) := X"0C027196";
        ram_buffer(6078) := X"24A583C8";
        ram_buffer(6079) := X"0C026DBB";
        ram_buffer(6080) := X"02002021";
        ram_buffer(6081) := X"00001021";
        ram_buffer(6082) := X"8FBF0E4C";
        ram_buffer(6083) := X"8FBE0E48";
        ram_buffer(6084) := X"8FB70E44";
        ram_buffer(6085) := X"8FB60E40";
        ram_buffer(6086) := X"8FB50E3C";
        ram_buffer(6087) := X"8FB40E38";
        ram_buffer(6088) := X"8FB30E34";
        ram_buffer(6089) := X"8FB20E30";
        ram_buffer(6090) := X"8FB10E2C";
        ram_buffer(6091) := X"8FB00E28";
        ram_buffer(6092) := X"03E00008";
        ram_buffer(6093) := X"27BD0E50";
        ram_buffer(6094) := X"2403003A";
        ram_buffer(6095) := X"1043003D";
        ram_buffer(6096) := X"AE7EFFF8";
        ram_buffer(6097) := X"2403003F";
        ram_buffer(6098) := X"AE60000C";
        ram_buffer(6099) := X"AE630010";
        ram_buffer(6100) := X"AE600014";
        ram_buffer(6101) := X"AE600018";
        ram_buffer(6102) := X"2403003B";
        ram_buffer(6103) := X"1043002A";
        ram_buffer(6104) := X"2403FFFF";
        ram_buffer(6105) := X"10430029";
        ram_buffer(6106) := X"26B50001";
        ram_buffer(6107) := X"8F828098";
        ram_buffer(6108) := X"3C05100D";
        ram_buffer(6109) := X"8C44000C";
        ram_buffer(6110) := X"02403021";
        ram_buffer(6111) := X"0C027196";
        ram_buffer(6112) := X"24A583F4";
        ram_buffer(6113) := X"0C026DBB";
        ram_buffer(6114) := X"02002021";
        ram_buffer(6115) := X"1000FFDE";
        ram_buffer(6116) := X"00001021";
        ram_buffer(6117) := X"8FA30E24";
        ram_buffer(6118) := X"2402FFFF";
        ram_buffer(6119) := X"1462006E";
        ram_buffer(6120) := X"3C05100D";
        ram_buffer(6121) := X"12A00014";
        ram_buffer(6122) := X"00158940";
        ram_buffer(6123) := X"8FA20E50";
        ram_buffer(6124) := X"00000000";
        ram_buffer(6125) := X"8C430004";
        ram_buffer(6126) := X"00151080";
        ram_buffer(6127) := X"00518821";
        ram_buffer(6128) := X"8FA40E50";
        ram_buffer(6129) := X"8C620000";
        ram_buffer(6130) := X"02203021";
        ram_buffer(6131) := X"0040F809";
        ram_buffer(6132) := X"24050001";
        ram_buffer(6133) := X"00402021";
        ram_buffer(6134) := X"02203021";
        ram_buffer(6135) := X"0C027F93";
        ram_buffer(6136) := X"27A50010";
        ram_buffer(6137) := X"00401821";
        ram_buffer(6138) := X"8FA20E50";
        ram_buffer(6139) := X"00000000";
        ram_buffer(6140) := X"AC4300A4";
        ram_buffer(6141) := X"AC5500A0";
        ram_buffer(6142) := X"0C026DBB";
        ram_buffer(6143) := X"02002021";
        ram_buffer(6144) := X"1000FFC1";
        ram_buffer(6145) := X"24020001";
        ram_buffer(6146) := X"26B50001";
        ram_buffer(6147) := X"1000FF90";
        ram_buffer(6148) := X"26730024";
        ram_buffer(6149) := X"8F828098";
        ram_buffer(6150) := X"3C05100D";
        ram_buffer(6151) := X"8C44000C";
        ram_buffer(6152) := X"02403021";
        ram_buffer(6153) := X"0C027196";
        ram_buffer(6154) := X"24A58380";
        ram_buffer(6155) := X"1000FFB6";
        ram_buffer(6156) := X"00001021";
        ram_buffer(6157) := X"27A60E24";
        ram_buffer(6158) := X"27A50E20";
        ram_buffer(6159) := X"0C02160B";
        ram_buffer(6160) := X"02002021";
        ram_buffer(6161) := X"1040FFC9";
        ram_buffer(6162) := X"00000000";
        ram_buffer(6163) := X"27A50E24";
        ram_buffer(6164) := X"0C0216A8";
        ram_buffer(6165) := X"02002021";
        ram_buffer(6166) := X"1040FFC4";
        ram_buffer(6167) := X"00000000";
        ram_buffer(6168) := X"8FA20E24";
        ram_buffer(6169) := X"00000000";
        ram_buffer(6170) := X"1451FFC0";
        ram_buffer(6171) := X"27A60E24";
        ram_buffer(6172) := X"8FA20E20";
        ram_buffer(6173) := X"27A50E20";
        ram_buffer(6174) := X"02002021";
        ram_buffer(6175) := X"0C02160B";
        ram_buffer(6176) := X"AE62000C";
        ram_buffer(6177) := X"1040FFB9";
        ram_buffer(6178) := X"00000000";
        ram_buffer(6179) := X"27A50E24";
        ram_buffer(6180) := X"0C0216A8";
        ram_buffer(6181) := X"02002021";
        ram_buffer(6182) := X"1040FFB4";
        ram_buffer(6183) := X"00000000";
        ram_buffer(6184) := X"8FA20E24";
        ram_buffer(6185) := X"00000000";
        ram_buffer(6186) := X"1451FFB0";
        ram_buffer(6187) := X"27A60E24";
        ram_buffer(6188) := X"8FA20E20";
        ram_buffer(6189) := X"27A50E20";
        ram_buffer(6190) := X"02002021";
        ram_buffer(6191) := X"0C02160B";
        ram_buffer(6192) := X"AE620010";
        ram_buffer(6193) := X"1040FFA9";
        ram_buffer(6194) := X"00000000";
        ram_buffer(6195) := X"27A50E24";
        ram_buffer(6196) := X"0C0216A8";
        ram_buffer(6197) := X"02002021";
        ram_buffer(6198) := X"1040FFA4";
        ram_buffer(6199) := X"00000000";
        ram_buffer(6200) := X"8FA20E24";
        ram_buffer(6201) := X"00000000";
        ram_buffer(6202) := X"1451FFA0";
        ram_buffer(6203) := X"27A60E24";
        ram_buffer(6204) := X"8FA20E20";
        ram_buffer(6205) := X"27A50E20";
        ram_buffer(6206) := X"02002021";
        ram_buffer(6207) := X"0C02160B";
        ram_buffer(6208) := X"AE620014";
        ram_buffer(6209) := X"1040FF99";
        ram_buffer(6210) := X"00000000";
        ram_buffer(6211) := X"27A50E24";
        ram_buffer(6212) := X"0C0216A8";
        ram_buffer(6213) := X"02002021";
        ram_buffer(6214) := X"1040FF94";
        ram_buffer(6215) := X"00000000";
        ram_buffer(6216) := X"8FA30E20";
        ram_buffer(6217) := X"8FA20E24";
        ram_buffer(6218) := X"1000FF8B";
        ram_buffer(6219) := X"AE630018";
        ram_buffer(6220) := X"8F828098";
        ram_buffer(6221) := X"00000000";
        ram_buffer(6222) := X"8C44000C";
        ram_buffer(6223) := X"02403021";
        ram_buffer(6224) := X"0C027196";
        ram_buffer(6225) := X"24A583A4";
        ram_buffer(6226) := X"0C026DBB";
        ram_buffer(6227) := X"02002021";
        ram_buffer(6228) := X"1000FF6D";
        ram_buffer(6229) := X"00001021";
        ram_buffer(6230) := X"8F828098";
        ram_buffer(6231) := X"00000000";
        ram_buffer(6232) := X"8C44000C";
        ram_buffer(6233) := X"02403021";
        ram_buffer(6234) := X"0C027196";
        ram_buffer(6235) := X"24A58360";
        ram_buffer(6236) := X"0C026DBB";
        ram_buffer(6237) := X"02002021";
        ram_buffer(6238) := X"1000FF63";
        ram_buffer(6239) := X"00001021";
        ram_buffer(6240) := X"27BDFFD0";
        ram_buffer(6241) := X"AFB20020";
        ram_buffer(6242) := X"3C12100D";
        ram_buffer(6243) := X"AFB40028";
        ram_buffer(6244) := X"AFB30024";
        ram_buffer(6245) := X"AFB1001C";
        ram_buffer(6246) := X"AFB00018";
        ram_buffer(6247) := X"AFBF002C";
        ram_buffer(6248) := X"0080A021";
        ram_buffer(6249) := X"00A08021";
        ram_buffer(6250) := X"AFA00010";
        ram_buffer(6251) := X"00008821";
        ram_buffer(6252) := X"2413002C";
        ram_buffer(6253) := X"10000009";
        ram_buffer(6254) := X"26528450";
        ram_buffer(6255) := X"8E82003C";
        ram_buffer(6256) := X"8FA30010";
        ram_buffer(6257) := X"00511021";
        ram_buffer(6258) := X"AC430010";
        ram_buffer(6259) := X"26310054";
        ram_buffer(6260) := X"24020348";
        ram_buffer(6261) := X"12220024";
        ram_buffer(6262) := X"24020001";
        ram_buffer(6263) := X"82020000";
        ram_buffer(6264) := X"00000000";
        ram_buffer(6265) := X"1040FFF5";
        ram_buffer(6266) := X"27A70014";
        ram_buffer(6267) := X"27A60010";
        ram_buffer(6268) := X"02402821";
        ram_buffer(6269) := X"02002021";
        ram_buffer(6270) := X"0C028409";
        ram_buffer(6271) := X"A3B30014";
        ram_buffer(6272) := X"18400021";
        ram_buffer(6273) := X"2402002C";
        ram_buffer(6274) := X"83A30014";
        ram_buffer(6275) := X"00000000";
        ram_buffer(6276) := X"1462001D";
        ram_buffer(6277) := X"00000000";
        ram_buffer(6278) := X"8FA40010";
        ram_buffer(6279) := X"00000000";
        ram_buffer(6280) := X"2C820004";
        ram_buffer(6281) := X"10400021";
        ram_buffer(6282) := X"3C05100D";
        ram_buffer(6283) := X"8E82003C";
        ram_buffer(6284) := X"2403002C";
        ram_buffer(6285) := X"00511021";
        ram_buffer(6286) := X"10000003";
        ram_buffer(6287) := X"AC440010";
        ram_buffer(6288) := X"1043FFE2";
        ram_buffer(6289) := X"26100001";
        ram_buffer(6290) := X"82020000";
        ram_buffer(6291) := X"00000000";
        ram_buffer(6292) := X"1440FFFB";
        ram_buffer(6293) := X"00000000";
        ram_buffer(6294) := X"26310054";
        ram_buffer(6295) := X"24020348";
        ram_buffer(6296) := X"1622FFDE";
        ram_buffer(6297) := X"24020001";
        ram_buffer(6298) := X"8FBF002C";
        ram_buffer(6299) := X"8FB40028";
        ram_buffer(6300) := X"8FB30024";
        ram_buffer(6301) := X"8FB20020";
        ram_buffer(6302) := X"8FB1001C";
        ram_buffer(6303) := X"8FB00018";
        ram_buffer(6304) := X"03E00008";
        ram_buffer(6305) := X"27BD0030";
        ram_buffer(6306) := X"8FBF002C";
        ram_buffer(6307) := X"8FB40028";
        ram_buffer(6308) := X"8FB30024";
        ram_buffer(6309) := X"8FB20020";
        ram_buffer(6310) := X"8FB1001C";
        ram_buffer(6311) := X"8FB00018";
        ram_buffer(6312) := X"00001021";
        ram_buffer(6313) := X"03E00008";
        ram_buffer(6314) := X"27BD0030";
        ram_buffer(6315) := X"8F828098";
        ram_buffer(6316) := X"00000000";
        ram_buffer(6317) := X"8C44000C";
        ram_buffer(6318) := X"24060003";
        ram_buffer(6319) := X"0C027196";
        ram_buffer(6320) := X"24A5841C";
        ram_buffer(6321) := X"1000FFE8";
        ram_buffer(6322) := X"00001021";
        ram_buffer(6323) := X"27BDFFC0";
        ram_buffer(6324) := X"AFB20034";
        ram_buffer(6325) := X"3C12100D";
        ram_buffer(6326) := X"AFB30038";
        ram_buffer(6327) := X"AFB10030";
        ram_buffer(6328) := X"AFB0002C";
        ram_buffer(6329) := X"AFBF003C";
        ram_buffer(6330) := X"00809821";
        ram_buffer(6331) := X"00A08021";
        ram_buffer(6332) := X"00008821";
        ram_buffer(6333) := X"1000000A";
        ram_buffer(6334) := X"2652844C";
        ram_buffer(6335) := X"8E62003C";
        ram_buffer(6336) := X"00000000";
        ram_buffer(6337) := X"00511021";
        ram_buffer(6338) := X"AC430008";
        ram_buffer(6339) := X"AC43000C";
        ram_buffer(6340) := X"26310054";
        ram_buffer(6341) := X"24020348";
        ram_buffer(6342) := X"1222003A";
        ram_buffer(6343) := X"00000000";
        ram_buffer(6344) := X"82020000";
        ram_buffer(6345) := X"00000000";
        ram_buffer(6346) := X"1040FFF4";
        ram_buffer(6347) := X"24030001";
        ram_buffer(6348) := X"27A20020";
        ram_buffer(6349) := X"AFA20014";
        ram_buffer(6350) := X"27A20018";
        ram_buffer(6351) := X"AFA20010";
        ram_buffer(6352) := X"27A70021";
        ram_buffer(6353) := X"2402002C";
        ram_buffer(6354) := X"27A6001C";
        ram_buffer(6355) := X"02402821";
        ram_buffer(6356) := X"02002021";
        ram_buffer(6357) := X"0C028409";
        ram_buffer(6358) := X"A3A20020";
        ram_buffer(6359) := X"28420003";
        ram_buffer(6360) := X"14400030";
        ram_buffer(6361) := X"24030058";
        ram_buffer(6362) := X"93A20021";
        ram_buffer(6363) := X"00000000";
        ram_buffer(6364) := X"304200DF";
        ram_buffer(6365) := X"00021600";
        ram_buffer(6366) := X"00021603";
        ram_buffer(6367) := X"14430029";
        ram_buffer(6368) := X"2402002C";
        ram_buffer(6369) := X"83A30020";
        ram_buffer(6370) := X"00000000";
        ram_buffer(6371) := X"14620025";
        ram_buffer(6372) := X"00000000";
        ram_buffer(6373) := X"8FA4001C";
        ram_buffer(6374) := X"00000000";
        ram_buffer(6375) := X"2482FFFF";
        ram_buffer(6376) := X"2C420004";
        ram_buffer(6377) := X"10400027";
        ram_buffer(6378) := X"00000000";
        ram_buffer(6379) := X"8FA50018";
        ram_buffer(6380) := X"00000000";
        ram_buffer(6381) := X"24A2FFFF";
        ram_buffer(6382) := X"2C420004";
        ram_buffer(6383) := X"10400021";
        ram_buffer(6384) := X"2403002C";
        ram_buffer(6385) := X"8E62003C";
        ram_buffer(6386) := X"00000000";
        ram_buffer(6387) := X"00511021";
        ram_buffer(6388) := X"AC440008";
        ram_buffer(6389) := X"10000003";
        ram_buffer(6390) := X"AC45000C";
        ram_buffer(6391) := X"1043FFCC";
        ram_buffer(6392) := X"26100001";
        ram_buffer(6393) := X"82020000";
        ram_buffer(6394) := X"00000000";
        ram_buffer(6395) := X"1440FFFB";
        ram_buffer(6396) := X"00000000";
        ram_buffer(6397) := X"26310054";
        ram_buffer(6398) := X"24020348";
        ram_buffer(6399) := X"1622FFC8";
        ram_buffer(6400) := X"00000000";
        ram_buffer(6401) := X"8FBF003C";
        ram_buffer(6402) := X"8FB30038";
        ram_buffer(6403) := X"8FB20034";
        ram_buffer(6404) := X"8FB10030";
        ram_buffer(6405) := X"8FB0002C";
        ram_buffer(6406) := X"24020001";
        ram_buffer(6407) := X"03E00008";
        ram_buffer(6408) := X"27BD0040";
        ram_buffer(6409) := X"8FBF003C";
        ram_buffer(6410) := X"8FB30038";
        ram_buffer(6411) := X"8FB20034";
        ram_buffer(6412) := X"8FB10030";
        ram_buffer(6413) := X"8FB0002C";
        ram_buffer(6414) := X"00001021";
        ram_buffer(6415) := X"03E00008";
        ram_buffer(6416) := X"27BD0040";
        ram_buffer(6417) := X"8F828098";
        ram_buffer(6418) := X"3C04100D";
        ram_buffer(6419) := X"8C47000C";
        ram_buffer(6420) := X"24060023";
        ram_buffer(6421) := X"24050001";
        ram_buffer(6422) := X"0C0278D7";
        ram_buffer(6423) := X"24848458";
        ram_buffer(6424) := X"8FBF003C";
        ram_buffer(6425) := X"8FB30038";
        ram_buffer(6426) := X"8FB20034";
        ram_buffer(6427) := X"8FB10030";
        ram_buffer(6428) := X"8FB0002C";
        ram_buffer(6429) := X"00001021";
        ram_buffer(6430) := X"03E00008";
        ram_buffer(6431) := X"27BD0040";
        ram_buffer(6432) := X"80820000";
        ram_buffer(6433) := X"24870001";
        ram_buffer(6434) := X"1040001C";
        ram_buffer(6435) := X"00401821";
        ram_buffer(6436) := X"80A80000";
        ram_buffer(6437) := X"00000000";
        ram_buffer(6438) := X"11000014";
        ram_buffer(6439) := X"24A50001";
        ram_buffer(6440) := X"8F8A8090";
        ram_buffer(6441) := X"24090001";
        ram_buffer(6442) := X"01421021";
        ram_buffer(6443) := X"90420001";
        ram_buffer(6444) := X"00E45823";
        ram_buffer(6445) := X"30420003";
        ram_buffer(6446) := X"24E70001";
        ram_buffer(6447) := X"1049000D";
        ram_buffer(6448) := X"24A50001";
        ram_buffer(6449) := X"14680009";
        ram_buffer(6450) := X"00000000";
        ram_buffer(6451) := X"80E3FFFF";
        ram_buffer(6452) := X"00000000";
        ram_buffer(6453) := X"1060000A";
        ram_buffer(6454) := X"00601021";
        ram_buffer(6455) := X"80A8FFFF";
        ram_buffer(6456) := X"00000000";
        ram_buffer(6457) := X"1500FFF0";
        ram_buffer(6458) := X"00000000";
        ram_buffer(6459) := X"03E00008";
        ram_buffer(6460) := X"00001021";
        ram_buffer(6461) := X"1000FFF3";
        ram_buffer(6462) := X"24630020";
        ram_buffer(6463) := X"00005821";
        ram_buffer(6464) := X"0166102A";
        ram_buffer(6465) := X"03E00008";
        ram_buffer(6466) := X"38420001";
        ram_buffer(6467) := X"8F828098";
        ram_buffer(6468) := X"00000000";
        ram_buffer(6469) := X"8C420004";
        ram_buffer(6470) := X"03E00008";
        ram_buffer(6471) := X"00000000";
        ram_buffer(6472) := X"8F828098";
        ram_buffer(6473) := X"00000000";
        ram_buffer(6474) := X"8C420008";
        ram_buffer(6475) := X"03E00008";
        ram_buffer(6476) := X"00000000";
        ram_buffer(6477) := X"27BDFFE0";
        ram_buffer(6478) := X"2402003D";
        ram_buffer(6479) := X"AFB10018";
        ram_buffer(6480) := X"AFB00014";
        ram_buffer(6481) := X"AFBF001C";
        ram_buffer(6482) := X"00808021";
        ram_buffer(6483) := X"00C08821";
        ram_buffer(6484) := X"10A2000D";
        ram_buffer(6485) := X"AC800004";
        ram_buffer(6486) := X"8C830000";
        ram_buffer(6487) := X"2406000A";
        ram_buffer(6488) := X"AC620018";
        ram_buffer(6489) := X"8C820000";
        ram_buffer(6490) := X"AC660014";
        ram_buffer(6491) := X"AC45001C";
        ram_buffer(6492) := X"8C820000";
        ram_buffer(6493) := X"00000000";
        ram_buffer(6494) := X"8C420000";
        ram_buffer(6495) := X"00000000";
        ram_buffer(6496) := X"0040F809";
        ram_buffer(6497) := X"00000000";
        ram_buffer(6498) := X"24020168";
        ram_buffer(6499) := X"1222000D";
        ram_buffer(6500) := X"24040013";
        ram_buffer(6501) := X"8E030000";
        ram_buffer(6502) := X"00000000";
        ram_buffer(6503) := X"AC620018";
        ram_buffer(6504) := X"8E020000";
        ram_buffer(6505) := X"AC640014";
        ram_buffer(6506) := X"AC51001C";
        ram_buffer(6507) := X"8E020000";
        ram_buffer(6508) := X"00000000";
        ram_buffer(6509) := X"8C420000";
        ram_buffer(6510) := X"00000000";
        ram_buffer(6511) := X"0040F809";
        ram_buffer(6512) := X"02002021";
        ram_buffer(6513) := X"8E110000";
        ram_buffer(6514) := X"24060168";
        ram_buffer(6515) := X"00002821";
        ram_buffer(6516) := X"0C02801D";
        ram_buffer(6517) := X"02002021";
        ram_buffer(6518) := X"02002021";
        ram_buffer(6519) := X"0C026CB7";
        ram_buffer(6520) := X"AE110000";
        ram_buffer(6521) := X"26040050";
        ram_buffer(6522) := X"24060010";
        ram_buffer(6523) := X"00002821";
        ram_buffer(6524) := X"AE000008";
        ram_buffer(6525) := X"AE000014";
        ram_buffer(6526) := X"AE00003C";
        ram_buffer(6527) := X"AE000040";
        ram_buffer(6528) := X"AE000044";
        ram_buffer(6529) := X"AE000048";
        ram_buffer(6530) := X"0C02801D";
        ram_buffer(6531) := X"AE00004C";
        ram_buffer(6532) := X"26040060";
        ram_buffer(6533) := X"24060010";
        ram_buffer(6534) := X"0C02801D";
        ram_buffer(6535) := X"00002821";
        ram_buffer(6536) := X"8F828020";
        ram_buffer(6537) := X"8FBF001C";
        ram_buffer(6538) := X"8F838024";
        ram_buffer(6539) := X"AE020028";
        ram_buffer(6540) := X"24020064";
        ram_buffer(6541) := X"AE03002C";
        ram_buffer(6542) := X"AE020010";
        ram_buffer(6543) := X"8FB10018";
        ram_buffer(6544) := X"8FB00014";
        ram_buffer(6545) := X"03E00008";
        ram_buffer(6546) := X"27BD0020";
        ram_buffer(6547) := X"08026485";
        ram_buffer(6548) := X"00000000";
        ram_buffer(6549) := X"0802646E";
        ram_buffer(6550) := X"00000000";
        ram_buffer(6551) := X"8C820040";
        ram_buffer(6552) := X"00000000";
        ram_buffer(6553) := X"10400002";
        ram_buffer(6554) := X"00000000";
        ram_buffer(6555) := X"AC450080";
        ram_buffer(6556) := X"8C820044";
        ram_buffer(6557) := X"00000000";
        ram_buffer(6558) := X"10400002";
        ram_buffer(6559) := X"00000000";
        ram_buffer(6560) := X"AC450080";
        ram_buffer(6561) := X"8C820048";
        ram_buffer(6562) := X"00000000";
        ram_buffer(6563) := X"10400002";
        ram_buffer(6564) := X"00000000";
        ram_buffer(6565) := X"AC450080";
        ram_buffer(6566) := X"8C82004C";
        ram_buffer(6567) := X"00000000";
        ram_buffer(6568) := X"10400002";
        ram_buffer(6569) := X"00000000";
        ram_buffer(6570) := X"AC450080";
        ram_buffer(6571) := X"8C820050";
        ram_buffer(6572) := X"00000000";
        ram_buffer(6573) := X"10400002";
        ram_buffer(6574) := X"00000000";
        ram_buffer(6575) := X"AC450114";
        ram_buffer(6576) := X"8C820060";
        ram_buffer(6577) := X"00000000";
        ram_buffer(6578) := X"10400002";
        ram_buffer(6579) := X"00000000";
        ram_buffer(6580) := X"AC450114";
        ram_buffer(6581) := X"8C820054";
        ram_buffer(6582) := X"00000000";
        ram_buffer(6583) := X"10400002";
        ram_buffer(6584) := X"00000000";
        ram_buffer(6585) := X"AC450114";
        ram_buffer(6586) := X"8C820064";
        ram_buffer(6587) := X"00000000";
        ram_buffer(6588) := X"10400002";
        ram_buffer(6589) := X"00000000";
        ram_buffer(6590) := X"AC450114";
        ram_buffer(6591) := X"8C820058";
        ram_buffer(6592) := X"00000000";
        ram_buffer(6593) := X"10400002";
        ram_buffer(6594) := X"00000000";
        ram_buffer(6595) := X"AC450114";
        ram_buffer(6596) := X"8C820068";
        ram_buffer(6597) := X"00000000";
        ram_buffer(6598) := X"10400002";
        ram_buffer(6599) := X"00000000";
        ram_buffer(6600) := X"AC450114";
        ram_buffer(6601) := X"8C82005C";
        ram_buffer(6602) := X"00000000";
        ram_buffer(6603) := X"10400002";
        ram_buffer(6604) := X"00000000";
        ram_buffer(6605) := X"AC450114";
        ram_buffer(6606) := X"8C82006C";
        ram_buffer(6607) := X"00000000";
        ram_buffer(6608) := X"10400002";
        ram_buffer(6609) := X"00000000";
        ram_buffer(6610) := X"AC450114";
        ram_buffer(6611) := X"03E00008";
        ram_buffer(6612) := X"00000000";
        ram_buffer(6613) := X"8C830010";
        ram_buffer(6614) := X"27BDFFE0";
        ram_buffer(6615) := X"2462FF9B";
        ram_buffer(6616) := X"2C420002";
        ram_buffer(6617) := X"AFB00010";
        ram_buffer(6618) := X"AFBF001C";
        ram_buffer(6619) := X"AFB20018";
        ram_buffer(6620) := X"AFB10014";
        ram_buffer(6621) := X"1440005C";
        ram_buffer(6622) := X"00808021";
        ram_buffer(6623) := X"24020067";
        ram_buffer(6624) := X"1062000A";
        ram_buffer(6625) := X"24050012";
        ram_buffer(6626) := X"8C820000";
        ram_buffer(6627) := X"00000000";
        ram_buffer(6628) := X"AC430018";
        ram_buffer(6629) := X"8C830000";
        ram_buffer(6630) := X"AC450014";
        ram_buffer(6631) := X"8C620000";
        ram_buffer(6632) := X"00000000";
        ram_buffer(6633) := X"0040F809";
        ram_buffer(6634) := X"00000000";
        ram_buffer(6635) := X"8E020144";
        ram_buffer(6636) := X"00000000";
        ram_buffer(6637) := X"8C430010";
        ram_buffer(6638) := X"00000000";
        ram_buffer(6639) := X"14600037";
        ram_buffer(6640) := X"24120016";
        ram_buffer(6641) := X"8C420000";
        ram_buffer(6642) := X"00000000";
        ram_buffer(6643) := X"0040F809";
        ram_buffer(6644) := X"02002021";
        ram_buffer(6645) := X"8E0300E8";
        ram_buffer(6646) := X"00000000";
        ram_buffer(6647) := X"14600008";
        ram_buffer(6648) := X"00008821";
        ram_buffer(6649) := X"10000021";
        ram_buffer(6650) := X"00000000";
        ram_buffer(6651) := X"8E0300E8";
        ram_buffer(6652) := X"00000000";
        ram_buffer(6653) := X"0223102B";
        ram_buffer(6654) := X"1040001C";
        ram_buffer(6655) := X"00000000";
        ram_buffer(6656) := X"8E020008";
        ram_buffer(6657) := X"00000000";
        ram_buffer(6658) := X"10400005";
        ram_buffer(6659) := X"02002021";
        ram_buffer(6660) := X"8C450000";
        ram_buffer(6661) := X"AC510004";
        ram_buffer(6662) := X"00A0F809";
        ram_buffer(6663) := X"AC430008";
        ram_buffer(6664) := X"8E020150";
        ram_buffer(6665) := X"02002021";
        ram_buffer(6666) := X"8C420004";
        ram_buffer(6667) := X"00002821";
        ram_buffer(6668) := X"0040F809";
        ram_buffer(6669) := X"26310001";
        ram_buffer(6670) := X"1440FFEC";
        ram_buffer(6671) := X"02002021";
        ram_buffer(6672) := X"8E020000";
        ram_buffer(6673) := X"00000000";
        ram_buffer(6674) := X"8C430000";
        ram_buffer(6675) := X"00000000";
        ram_buffer(6676) := X"0060F809";
        ram_buffer(6677) := X"AC520014";
        ram_buffer(6678) := X"8E0300E8";
        ram_buffer(6679) := X"00000000";
        ram_buffer(6680) := X"0223102B";
        ram_buffer(6681) := X"1440FFE6";
        ram_buffer(6682) := X"00000000";
        ram_buffer(6683) := X"8E020144";
        ram_buffer(6684) := X"00000000";
        ram_buffer(6685) := X"8C420008";
        ram_buffer(6686) := X"00000000";
        ram_buffer(6687) := X"0040F809";
        ram_buffer(6688) := X"02002021";
        ram_buffer(6689) := X"8E020144";
        ram_buffer(6690) := X"00000000";
        ram_buffer(6691) := X"8C430010";
        ram_buffer(6692) := X"00000000";
        ram_buffer(6693) := X"1060FFCB";
        ram_buffer(6694) := X"00000000";
        ram_buffer(6695) := X"8E020154";
        ram_buffer(6696) := X"00000000";
        ram_buffer(6697) := X"8C420010";
        ram_buffer(6698) := X"00000000";
        ram_buffer(6699) := X"0040F809";
        ram_buffer(6700) := X"02002021";
        ram_buffer(6701) := X"8E020014";
        ram_buffer(6702) := X"00000000";
        ram_buffer(6703) := X"8C420010";
        ram_buffer(6704) := X"00000000";
        ram_buffer(6705) := X"0040F809";
        ram_buffer(6706) := X"02002021";
        ram_buffer(6707) := X"8FBF001C";
        ram_buffer(6708) := X"8FB20018";
        ram_buffer(6709) := X"8FB10014";
        ram_buffer(6710) := X"02002021";
        ram_buffer(6711) := X"8FB00010";
        ram_buffer(6712) := X"0802646E";
        ram_buffer(6713) := X"27BD0020";
        ram_buffer(6714) := X"8C8200D8";
        ram_buffer(6715) := X"8C83001C";
        ram_buffer(6716) := X"00000000";
        ram_buffer(6717) := X"0043102B";
        ram_buffer(6718) := X"14400009";
        ram_buffer(6719) := X"24050042";
        ram_buffer(6720) := X"8E020144";
        ram_buffer(6721) := X"00000000";
        ram_buffer(6722) := X"8C420008";
        ram_buffer(6723) := X"00000000";
        ram_buffer(6724) := X"0040F809";
        ram_buffer(6725) := X"02002021";
        ram_buffer(6726) := X"1000FFA4";
        ram_buffer(6727) := X"00000000";
        ram_buffer(6728) := X"8C820000";
        ram_buffer(6729) := X"00000000";
        ram_buffer(6730) := X"8C430000";
        ram_buffer(6731) := X"00000000";
        ram_buffer(6732) := X"0060F809";
        ram_buffer(6733) := X"AC450014";
        ram_buffer(6734) := X"1000FFF1";
        ram_buffer(6735) := X"00000000";
        ram_buffer(6736) := X"8C8200D8";
        ram_buffer(6737) := X"27BDFFD8";
        ram_buffer(6738) := X"8C830010";
        ram_buffer(6739) := X"AFB00020";
        ram_buffer(6740) := X"AFBF0024";
        ram_buffer(6741) := X"14400005";
        ram_buffer(6742) := X"00808021";
        ram_buffer(6743) := X"2462FF9B";
        ram_buffer(6744) := X"2C420003";
        ram_buffer(6745) := X"1440000F";
        ram_buffer(6746) := X"00000000";
        ram_buffer(6747) := X"8E020000";
        ram_buffer(6748) := X"24040012";
        ram_buffer(6749) := X"AC430018";
        ram_buffer(6750) := X"8E030000";
        ram_buffer(6751) := X"AC440014";
        ram_buffer(6752) := X"8C620000";
        ram_buffer(6753) := X"02002021";
        ram_buffer(6754) := X"AFA70018";
        ram_buffer(6755) := X"AFA60014";
        ram_buffer(6756) := X"0040F809";
        ram_buffer(6757) := X"AFA50010";
        ram_buffer(6758) := X"8FA70018";
        ram_buffer(6759) := X"8FA60014";
        ram_buffer(6760) := X"8FA50010";
        ram_buffer(6761) := X"8E020154";
        ram_buffer(6762) := X"8FBF0024";
        ram_buffer(6763) := X"8C590000";
        ram_buffer(6764) := X"02002021";
        ram_buffer(6765) := X"8FB00020";
        ram_buffer(6766) := X"03200008";
        ram_buffer(6767) := X"27BD0028";
        ram_buffer(6768) := X"8C820010";
        ram_buffer(6769) := X"27BDFFE8";
        ram_buffer(6770) := X"24030064";
        ram_buffer(6771) := X"AFB00010";
        ram_buffer(6772) := X"AFBF0014";
        ram_buffer(6773) := X"1043000A";
        ram_buffer(6774) := X"00808021";
        ram_buffer(6775) := X"8C830000";
        ram_buffer(6776) := X"24050012";
        ram_buffer(6777) := X"AC620018";
        ram_buffer(6778) := X"8C820000";
        ram_buffer(6779) := X"AC650014";
        ram_buffer(6780) := X"8C420000";
        ram_buffer(6781) := X"00000000";
        ram_buffer(6782) := X"0040F809";
        ram_buffer(6783) := X"00000000";
        ram_buffer(6784) := X"8E020000";
        ram_buffer(6785) := X"00000000";
        ram_buffer(6786) := X"8C420010";
        ram_buffer(6787) := X"00000000";
        ram_buffer(6788) := X"0040F809";
        ram_buffer(6789) := X"02002021";
        ram_buffer(6790) := X"8E020014";
        ram_buffer(6791) := X"00000000";
        ram_buffer(6792) := X"8C420008";
        ram_buffer(6793) := X"00000000";
        ram_buffer(6794) := X"0040F809";
        ram_buffer(6795) := X"02002021";
        ram_buffer(6796) := X"0C023694";
        ram_buffer(6797) := X"02002021";
        ram_buffer(6798) := X"8E020154";
        ram_buffer(6799) := X"00000000";
        ram_buffer(6800) := X"8C420014";
        ram_buffer(6801) := X"00000000";
        ram_buffer(6802) := X"0040F809";
        ram_buffer(6803) := X"02002021";
        ram_buffer(6804) := X"8E020014";
        ram_buffer(6805) := X"00000000";
        ram_buffer(6806) := X"8C420010";
        ram_buffer(6807) := X"00000000";
        ram_buffer(6808) := X"0040F809";
        ram_buffer(6809) := X"02002021";
        ram_buffer(6810) := X"8FBF0014";
        ram_buffer(6811) := X"02002021";
        ram_buffer(6812) := X"8FB00010";
        ram_buffer(6813) := X"0802646E";
        ram_buffer(6814) := X"27BD0018";
        ram_buffer(6815) := X"8C820010";
        ram_buffer(6816) := X"27BDFFE0";
        ram_buffer(6817) := X"24030064";
        ram_buffer(6818) := X"AFB10018";
        ram_buffer(6819) := X"AFB00014";
        ram_buffer(6820) := X"AFBF001C";
        ram_buffer(6821) := X"00808021";
        ram_buffer(6822) := X"1043000A";
        ram_buffer(6823) := X"00A08821";
        ram_buffer(6824) := X"8C830000";
        ram_buffer(6825) := X"24050012";
        ram_buffer(6826) := X"AC620018";
        ram_buffer(6827) := X"8C820000";
        ram_buffer(6828) := X"AC650014";
        ram_buffer(6829) := X"8C420000";
        ram_buffer(6830) := X"00000000";
        ram_buffer(6831) := X"0040F809";
        ram_buffer(6832) := X"00000000";
        ram_buffer(6833) := X"1620001F";
        ram_buffer(6834) := X"00002821";
        ram_buffer(6835) := X"8E020000";
        ram_buffer(6836) := X"00000000";
        ram_buffer(6837) := X"8C420010";
        ram_buffer(6838) := X"00000000";
        ram_buffer(6839) := X"0040F809";
        ram_buffer(6840) := X"02002021";
        ram_buffer(6841) := X"8E020014";
        ram_buffer(6842) := X"00000000";
        ram_buffer(6843) := X"8C420008";
        ram_buffer(6844) := X"00000000";
        ram_buffer(6845) := X"0040F809";
        ram_buffer(6846) := X"02002021";
        ram_buffer(6847) := X"0C022282";
        ram_buffer(6848) := X"02002021";
        ram_buffer(6849) := X"8E020144";
        ram_buffer(6850) := X"00000000";
        ram_buffer(6851) := X"8C420000";
        ram_buffer(6852) := X"00000000";
        ram_buffer(6853) := X"0040F809";
        ram_buffer(6854) := X"02002021";
        ram_buffer(6855) := X"8E0200A8";
        ram_buffer(6856) := X"8FBF001C";
        ram_buffer(6857) := X"0002102B";
        ram_buffer(6858) := X"24420065";
        ram_buffer(6859) := X"AE0000D8";
        ram_buffer(6860) := X"AE020010";
        ram_buffer(6861) := X"8FB10018";
        ram_buffer(6862) := X"8FB00014";
        ram_buffer(6863) := X"03E00008";
        ram_buffer(6864) := X"27BD0020";
        ram_buffer(6865) := X"0C021997";
        ram_buffer(6866) := X"02002021";
        ram_buffer(6867) := X"1000FFDF";
        ram_buffer(6868) := X"00000000";
        ram_buffer(6869) := X"8C820010";
        ram_buffer(6870) := X"27BDFFD8";
        ram_buffer(6871) := X"24030065";
        ram_buffer(6872) := X"AFB20020";
        ram_buffer(6873) := X"AFB1001C";
        ram_buffer(6874) := X"AFB00018";
        ram_buffer(6875) := X"AFBF0024";
        ram_buffer(6876) := X"00808021";
        ram_buffer(6877) := X"00A09021";
        ram_buffer(6878) := X"1043000A";
        ram_buffer(6879) := X"00C08821";
        ram_buffer(6880) := X"8C830000";
        ram_buffer(6881) := X"24050012";
        ram_buffer(6882) := X"AC620018";
        ram_buffer(6883) := X"8C820000";
        ram_buffer(6884) := X"AC650014";
        ram_buffer(6885) := X"8C420000";
        ram_buffer(6886) := X"00000000";
        ram_buffer(6887) := X"0040F809";
        ram_buffer(6888) := X"00000000";
        ram_buffer(6889) := X"8E0200D8";
        ram_buffer(6890) := X"8E03001C";
        ram_buffer(6891) := X"00000000";
        ram_buffer(6892) := X"0043102B";
        ram_buffer(6893) := X"1040002B";
        ram_buffer(6894) := X"24040077";
        ram_buffer(6895) := X"8E020008";
        ram_buffer(6896) := X"00000000";
        ram_buffer(6897) := X"10400008";
        ram_buffer(6898) := X"00000000";
        ram_buffer(6899) := X"8E04001C";
        ram_buffer(6900) := X"8E0500D8";
        ram_buffer(6901) := X"8C430000";
        ram_buffer(6902) := X"AC440008";
        ram_buffer(6903) := X"AC450004";
        ram_buffer(6904) := X"0060F809";
        ram_buffer(6905) := X"02002021";
        ram_buffer(6906) := X"8E020144";
        ram_buffer(6907) := X"00000000";
        ram_buffer(6908) := X"8C43000C";
        ram_buffer(6909) := X"00000000";
        ram_buffer(6910) := X"14600023";
        ram_buffer(6911) := X"00000000";
        ram_buffer(6912) := X"8E02001C";
        ram_buffer(6913) := X"8E0700D8";
        ram_buffer(6914) := X"AFA00010";
        ram_buffer(6915) := X"00473823";
        ram_buffer(6916) := X"0227182B";
        ram_buffer(6917) := X"8E020148";
        ram_buffer(6918) := X"10600002";
        ram_buffer(6919) := X"00000000";
        ram_buffer(6920) := X"02203821";
        ram_buffer(6921) := X"8C420004";
        ram_buffer(6922) := X"02002021";
        ram_buffer(6923) := X"27A60010";
        ram_buffer(6924) := X"0040F809";
        ram_buffer(6925) := X"02402821";
        ram_buffer(6926) := X"8FA40010";
        ram_buffer(6927) := X"8E0300D8";
        ram_buffer(6928) := X"8FBF0024";
        ram_buffer(6929) := X"00641821";
        ram_buffer(6930) := X"AE0300D8";
        ram_buffer(6931) := X"8FB20020";
        ram_buffer(6932) := X"8FB1001C";
        ram_buffer(6933) := X"8FB00018";
        ram_buffer(6934) := X"00801021";
        ram_buffer(6935) := X"03E00008";
        ram_buffer(6936) := X"27BD0028";
        ram_buffer(6937) := X"8E020000";
        ram_buffer(6938) := X"00000000";
        ram_buffer(6939) := X"8C430004";
        ram_buffer(6940) := X"AC440014";
        ram_buffer(6941) := X"2405FFFF";
        ram_buffer(6942) := X"0060F809";
        ram_buffer(6943) := X"02002021";
        ram_buffer(6944) := X"1000FFCE";
        ram_buffer(6945) := X"00000000";
        ram_buffer(6946) := X"8C420004";
        ram_buffer(6947) := X"00000000";
        ram_buffer(6948) := X"0040F809";
        ram_buffer(6949) := X"02002021";
        ram_buffer(6950) := X"1000FFD9";
        ram_buffer(6951) := X"00000000";
        ram_buffer(6952) := X"8C820010";
        ram_buffer(6953) := X"27BDFFD8";
        ram_buffer(6954) := X"24030066";
        ram_buffer(6955) := X"AFB30020";
        ram_buffer(6956) := X"AFB2001C";
        ram_buffer(6957) := X"AFB00014";
        ram_buffer(6958) := X"AFBF0024";
        ram_buffer(6959) := X"AFB10018";
        ram_buffer(6960) := X"00808021";
        ram_buffer(6961) := X"00A09821";
        ram_buffer(6962) := X"1043000A";
        ram_buffer(6963) := X"00C09021";
        ram_buffer(6964) := X"8C830000";
        ram_buffer(6965) := X"24050012";
        ram_buffer(6966) := X"AC620018";
        ram_buffer(6967) := X"8C820000";
        ram_buffer(6968) := X"AC650014";
        ram_buffer(6969) := X"8C420000";
        ram_buffer(6970) := X"00000000";
        ram_buffer(6971) := X"0040F809";
        ram_buffer(6972) := X"00000000";
        ram_buffer(6973) := X"8E0400D8";
        ram_buffer(6974) := X"8E03001C";
        ram_buffer(6975) := X"00000000";
        ram_buffer(6976) := X"0083102B";
        ram_buffer(6977) := X"1040003E";
        ram_buffer(6978) := X"2405FFFF";
        ram_buffer(6979) := X"8E020008";
        ram_buffer(6980) := X"00000000";
        ram_buffer(6981) := X"10400006";
        ram_buffer(6982) := X"00000000";
        ram_buffer(6983) := X"8C450000";
        ram_buffer(6984) := X"AC440004";
        ram_buffer(6985) := X"AC430008";
        ram_buffer(6986) := X"00A0F809";
        ram_buffer(6987) := X"02002021";
        ram_buffer(6988) := X"8E020144";
        ram_buffer(6989) := X"00000000";
        ram_buffer(6990) := X"8C43000C";
        ram_buffer(6991) := X"00000000";
        ram_buffer(6992) := X"14600029";
        ram_buffer(6993) := X"00000000";
        ram_buffer(6994) := X"8E1100E4";
        ram_buffer(6995) := X"00000000";
        ram_buffer(6996) := X"001188C0";
        ram_buffer(6997) := X"0251902B";
        ram_buffer(6998) := X"1640001B";
        ram_buffer(6999) := X"24040015";
        ram_buffer(7000) := X"8E020150";
        ram_buffer(7001) := X"02602821";
        ram_buffer(7002) := X"8C420004";
        ram_buffer(7003) := X"00000000";
        ram_buffer(7004) := X"0040F809";
        ram_buffer(7005) := X"02002021";
        ram_buffer(7006) := X"1040000B";
        ram_buffer(7007) := X"02201021";
        ram_buffer(7008) := X"8E0300D8";
        ram_buffer(7009) := X"8FBF0024";
        ram_buffer(7010) := X"00718821";
        ram_buffer(7011) := X"AE1100D8";
        ram_buffer(7012) := X"8FB30020";
        ram_buffer(7013) := X"8FB2001C";
        ram_buffer(7014) := X"8FB10018";
        ram_buffer(7015) := X"8FB00014";
        ram_buffer(7016) := X"03E00008";
        ram_buffer(7017) := X"27BD0028";
        ram_buffer(7018) := X"8FBF0024";
        ram_buffer(7019) := X"8FB30020";
        ram_buffer(7020) := X"8FB2001C";
        ram_buffer(7021) := X"8FB10018";
        ram_buffer(7022) := X"8FB00014";
        ram_buffer(7023) := X"00001021";
        ram_buffer(7024) := X"03E00008";
        ram_buffer(7025) := X"27BD0028";
        ram_buffer(7026) := X"8E020000";
        ram_buffer(7027) := X"00000000";
        ram_buffer(7028) := X"8C430000";
        ram_buffer(7029) := X"AC440014";
        ram_buffer(7030) := X"0060F809";
        ram_buffer(7031) := X"02002021";
        ram_buffer(7032) := X"1000FFDF";
        ram_buffer(7033) := X"00000000";
        ram_buffer(7034) := X"8C420004";
        ram_buffer(7035) := X"00000000";
        ram_buffer(7036) := X"0040F809";
        ram_buffer(7037) := X"02002021";
        ram_buffer(7038) := X"1000FFD3";
        ram_buffer(7039) := X"00000000";
        ram_buffer(7040) := X"8E020000";
        ram_buffer(7041) := X"24040077";
        ram_buffer(7042) := X"8C430004";
        ram_buffer(7043) := X"AC440014";
        ram_buffer(7044) := X"0060F809";
        ram_buffer(7045) := X"02002021";
        ram_buffer(7046) := X"8FBF0024";
        ram_buffer(7047) := X"8FB30020";
        ram_buffer(7048) := X"8FB2001C";
        ram_buffer(7049) := X"8FB10018";
        ram_buffer(7050) := X"8FB00014";
        ram_buffer(7051) := X"00001021";
        ram_buffer(7052) := X"03E00008";
        ram_buffer(7053) := X"27BD0028";
        ram_buffer(7054) := X"8C820010";
        ram_buffer(7055) := X"27BDFFD0";
        ram_buffer(7056) := X"24030064";
        ram_buffer(7057) := X"AFB30028";
        ram_buffer(7058) := X"AFB20024";
        ram_buffer(7059) := X"AFB10020";
        ram_buffer(7060) := X"AFBF002C";
        ram_buffer(7061) := X"AFB0001C";
        ram_buffer(7062) := X"00808821";
        ram_buffer(7063) := X"00C09021";
        ram_buffer(7064) := X"1043000C";
        ram_buffer(7065) := X"00E09821";
        ram_buffer(7066) := X"8C830000";
        ram_buffer(7067) := X"24080012";
        ram_buffer(7068) := X"AC620018";
        ram_buffer(7069) := X"8C820000";
        ram_buffer(7070) := X"AC680014";
        ram_buffer(7071) := X"8C420000";
        ram_buffer(7072) := X"00000000";
        ram_buffer(7073) := X"0040F809";
        ram_buffer(7074) := X"AFA50010";
        ram_buffer(7075) := X"8FA50010";
        ram_buffer(7076) := X"00000000";
        ram_buffer(7077) := X"00052880";
        ram_buffer(7078) := X"02258021";
        ram_buffer(7079) := X"8E020040";
        ram_buffer(7080) := X"00000000";
        ram_buffer(7081) := X"10400042";
        ram_buffer(7082) := X"00000000";
        ram_buffer(7083) := X"8FA30040";
        ram_buffer(7084) := X"02403021";
        ram_buffer(7085) := X"14600026";
        ram_buffer(7086) := X"00402021";
        ram_buffer(7087) := X"264B0100";
        ram_buffer(7088) := X"24080064";
        ram_buffer(7089) := X"10000007";
        ram_buffer(7090) := X"340A8000";
        ram_buffer(7091) := X"1520001E";
        ram_buffer(7092) := X"00000000";
        ram_buffer(7093) := X"24C60004";
        ram_buffer(7094) := X"A4850000";
        ram_buffer(7095) := X"11660012";
        ram_buffer(7096) := X"24840002";
        ram_buffer(7097) := X"8CC30000";
        ram_buffer(7098) := X"24057FFF";
        ram_buffer(7099) := X"02630018";
        ram_buffer(7100) := X"00001812";
        ram_buffer(7101) := X"24630032";
        ram_buffer(7102) := X"00000000";
        ram_buffer(7103) := X"15000002";
        ram_buffer(7104) := X"0068001A";
        ram_buffer(7105) := X"0007000D";
        ram_buffer(7106) := X"00001812";
        ram_buffer(7107) := X"1C60FFEF";
        ram_buffer(7108) := X"006A482A";
        ram_buffer(7109) := X"24050001";
        ram_buffer(7110) := X"24C60004";
        ram_buffer(7111) := X"A4850000";
        ram_buffer(7112) := X"1566FFF0";
        ram_buffer(7113) := X"24840002";
        ram_buffer(7114) := X"8FBF002C";
        ram_buffer(7115) := X"8FB30028";
        ram_buffer(7116) := X"8FB20024";
        ram_buffer(7117) := X"8FB10020";
        ram_buffer(7118) := X"8FB0001C";
        ram_buffer(7119) := X"AC400080";
        ram_buffer(7120) := X"03E00008";
        ram_buffer(7121) := X"27BD0030";
        ram_buffer(7122) := X"1000FFE2";
        ram_buffer(7123) := X"3065FFFF";
        ram_buffer(7124) := X"26490100";
        ram_buffer(7125) := X"10000008";
        ram_buffer(7126) := X"24050064";
        ram_buffer(7127) := X"11000018";
        ram_buffer(7128) := X"00000000";
        ram_buffer(7129) := X"3063FFFF";
        ram_buffer(7130) := X"24C60004";
        ram_buffer(7131) := X"A4830000";
        ram_buffer(7132) := X"1126FFED";
        ram_buffer(7133) := X"24840002";
        ram_buffer(7134) := X"8CC30000";
        ram_buffer(7135) := X"00000000";
        ram_buffer(7136) := X"02630018";
        ram_buffer(7137) := X"00001812";
        ram_buffer(7138) := X"24630032";
        ram_buffer(7139) := X"00000000";
        ram_buffer(7140) := X"14A00002";
        ram_buffer(7141) := X"0065001A";
        ram_buffer(7142) := X"0007000D";
        ram_buffer(7143) := X"00001812";
        ram_buffer(7144) := X"1C60FFEE";
        ram_buffer(7145) := X"28680100";
        ram_buffer(7146) := X"1000FFEF";
        ram_buffer(7147) := X"24030001";
        ram_buffer(7148) := X"0C026495";
        ram_buffer(7149) := X"02202021";
        ram_buffer(7150) := X"1000FFBC";
        ram_buffer(7151) := X"AE020040";
        ram_buffer(7152) := X"1000FFE9";
        ram_buffer(7153) := X"240300FF";
        ram_buffer(7154) := X"8C820010";
        ram_buffer(7155) := X"27BDFFE0";
        ram_buffer(7156) := X"24030064";
        ram_buffer(7157) := X"AFB20018";
        ram_buffer(7158) := X"AFB10014";
        ram_buffer(7159) := X"AFB00010";
        ram_buffer(7160) := X"AFBF001C";
        ram_buffer(7161) := X"00808821";
        ram_buffer(7162) := X"00A08021";
        ram_buffer(7163) := X"1043000A";
        ram_buffer(7164) := X"00C09021";
        ram_buffer(7165) := X"8C830000";
        ram_buffer(7166) := X"24050012";
        ram_buffer(7167) := X"AC620018";
        ram_buffer(7168) := X"8C820000";
        ram_buffer(7169) := X"AC650014";
        ram_buffer(7170) := X"8C420000";
        ram_buffer(7171) := X"00000000";
        ram_buffer(7172) := X"0040F809";
        ram_buffer(7173) := X"00000000";
        ram_buffer(7174) := X"8E220040";
        ram_buffer(7175) := X"00000000";
        ram_buffer(7176) := X"1040008E";
        ram_buffer(7177) := X"00000000";
        ram_buffer(7178) := X"3C04100D";
        ram_buffer(7179) := X"3C06100D";
        ram_buffer(7180) := X"24848774";
        ram_buffer(7181) := X"00402821";
        ram_buffer(7182) := X"16400071";
        ram_buffer(7183) := X"24C68874";
        ram_buffer(7184) := X"24080064";
        ram_buffer(7185) := X"10000007";
        ram_buffer(7186) := X"340A8000";
        ram_buffer(7187) := X"1520004F";
        ram_buffer(7188) := X"00000000";
        ram_buffer(7189) := X"24840004";
        ram_buffer(7190) := X"A4A70000";
        ram_buffer(7191) := X"10860012";
        ram_buffer(7192) := X"24A50002";
        ram_buffer(7193) := X"8C830000";
        ram_buffer(7194) := X"24077FFF";
        ram_buffer(7195) := X"02030018";
        ram_buffer(7196) := X"00001812";
        ram_buffer(7197) := X"24630032";
        ram_buffer(7198) := X"00000000";
        ram_buffer(7199) := X"15000002";
        ram_buffer(7200) := X"0068001A";
        ram_buffer(7201) := X"0007000D";
        ram_buffer(7202) := X"00001812";
        ram_buffer(7203) := X"1C60FFEF";
        ram_buffer(7204) := X"006A482A";
        ram_buffer(7205) := X"24070001";
        ram_buffer(7206) := X"24840004";
        ram_buffer(7207) := X"A4A70000";
        ram_buffer(7208) := X"1486FFF0";
        ram_buffer(7209) := X"24A50002";
        ram_buffer(7210) := X"8E230010";
        ram_buffer(7211) := X"AC400080";
        ram_buffer(7212) := X"24020064";
        ram_buffer(7213) := X"1062000A";
        ram_buffer(7214) := X"24040012";
        ram_buffer(7215) := X"8E220000";
        ram_buffer(7216) := X"00000000";
        ram_buffer(7217) := X"AC430018";
        ram_buffer(7218) := X"8E230000";
        ram_buffer(7219) := X"AC440014";
        ram_buffer(7220) := X"8C620000";
        ram_buffer(7221) := X"00000000";
        ram_buffer(7222) := X"0040F809";
        ram_buffer(7223) := X"02202021";
        ram_buffer(7224) := X"8E220044";
        ram_buffer(7225) := X"00000000";
        ram_buffer(7226) := X"10400060";
        ram_buffer(7227) := X"00000000";
        ram_buffer(7228) := X"3C04100D";
        ram_buffer(7229) := X"24848674";
        ram_buffer(7230) := X"16400028";
        ram_buffer(7231) := X"00402821";
        ram_buffer(7232) := X"3C09100D";
        ram_buffer(7233) := X"25298774";
        ram_buffer(7234) := X"24070064";
        ram_buffer(7235) := X"10000007";
        ram_buffer(7236) := X"340A8000";
        ram_buffer(7237) := X"1500001F";
        ram_buffer(7238) := X"00000000";
        ram_buffer(7239) := X"24840004";
        ram_buffer(7240) := X"A4A60000";
        ram_buffer(7241) := X"10890012";
        ram_buffer(7242) := X"24A50002";
        ram_buffer(7243) := X"8C830000";
        ram_buffer(7244) := X"24067FFF";
        ram_buffer(7245) := X"02030018";
        ram_buffer(7246) := X"00001812";
        ram_buffer(7247) := X"24630032";
        ram_buffer(7248) := X"00000000";
        ram_buffer(7249) := X"14E00002";
        ram_buffer(7250) := X"0067001A";
        ram_buffer(7251) := X"0007000D";
        ram_buffer(7252) := X"00001812";
        ram_buffer(7253) := X"1C60FFEF";
        ram_buffer(7254) := X"006A402A";
        ram_buffer(7255) := X"24060001";
        ram_buffer(7256) := X"24840004";
        ram_buffer(7257) := X"A4A60000";
        ram_buffer(7258) := X"1489FFF0";
        ram_buffer(7259) := X"24A50002";
        ram_buffer(7260) := X"8FBF001C";
        ram_buffer(7261) := X"8FB20018";
        ram_buffer(7262) := X"8FB10014";
        ram_buffer(7263) := X"8FB00010";
        ram_buffer(7264) := X"AC400080";
        ram_buffer(7265) := X"03E00008";
        ram_buffer(7266) := X"27BD0020";
        ram_buffer(7267) := X"1000FFB1";
        ram_buffer(7268) := X"3067FFFF";
        ram_buffer(7269) := X"1000FFE1";
        ram_buffer(7270) := X"3066FFFF";
        ram_buffer(7271) := X"3C08100D";
        ram_buffer(7272) := X"25088774";
        ram_buffer(7273) := X"10000008";
        ram_buffer(7274) := X"24060064";
        ram_buffer(7275) := X"10E00033";
        ram_buffer(7276) := X"00000000";
        ram_buffer(7277) := X"3063FFFF";
        ram_buffer(7278) := X"24840004";
        ram_buffer(7279) := X"A4A30000";
        ram_buffer(7280) := X"1088FFEB";
        ram_buffer(7281) := X"24A50002";
        ram_buffer(7282) := X"8C830000";
        ram_buffer(7283) := X"00000000";
        ram_buffer(7284) := X"02030018";
        ram_buffer(7285) := X"00001812";
        ram_buffer(7286) := X"24630032";
        ram_buffer(7287) := X"00000000";
        ram_buffer(7288) := X"14C00002";
        ram_buffer(7289) := X"0066001A";
        ram_buffer(7290) := X"0007000D";
        ram_buffer(7291) := X"00001812";
        ram_buffer(7292) := X"1C60FFEE";
        ram_buffer(7293) := X"28670100";
        ram_buffer(7294) := X"1000FFEF";
        ram_buffer(7295) := X"24030001";
        ram_buffer(7296) := X"10000008";
        ram_buffer(7297) := X"24070064";
        ram_buffer(7298) := X"1100001E";
        ram_buffer(7299) := X"00000000";
        ram_buffer(7300) := X"3063FFFF";
        ram_buffer(7301) := X"24840004";
        ram_buffer(7302) := X"A4A30000";
        ram_buffer(7303) := X"1086FFA2";
        ram_buffer(7304) := X"24A50002";
        ram_buffer(7305) := X"8C830000";
        ram_buffer(7306) := X"00000000";
        ram_buffer(7307) := X"02030018";
        ram_buffer(7308) := X"00001812";
        ram_buffer(7309) := X"24630032";
        ram_buffer(7310) := X"00000000";
        ram_buffer(7311) := X"14E00002";
        ram_buffer(7312) := X"0067001A";
        ram_buffer(7313) := X"0007000D";
        ram_buffer(7314) := X"00001812";
        ram_buffer(7315) := X"1C60FFEE";
        ram_buffer(7316) := X"28680100";
        ram_buffer(7317) := X"1000FFEF";
        ram_buffer(7318) := X"24030001";
        ram_buffer(7319) := X"0C026495";
        ram_buffer(7320) := X"02202021";
        ram_buffer(7321) := X"1000FF70";
        ram_buffer(7322) := X"AE220040";
        ram_buffer(7323) := X"0C026495";
        ram_buffer(7324) := X"02202021";
        ram_buffer(7325) := X"1000FF9E";
        ram_buffer(7326) := X"AE220044";
        ram_buffer(7327) := X"1000FFCE";
        ram_buffer(7328) := X"240300FF";
        ram_buffer(7329) := X"1000FFE3";
        ram_buffer(7330) := X"240300FF";
        ram_buffer(7331) := X"18800006";
        ram_buffer(7332) := X"00000000";
        ram_buffer(7333) := X"28820065";
        ram_buffer(7334) := X"14400005";
        ram_buffer(7335) := X"00001021";
        ram_buffer(7336) := X"03E00008";
        ram_buffer(7337) := X"00000000";
        ram_buffer(7338) := X"03E00008";
        ram_buffer(7339) := X"24021388";
        ram_buffer(7340) := X"28820032";
        ram_buffer(7341) := X"10400008";
        ram_buffer(7342) := X"00000000";
        ram_buffer(7343) := X"24021388";
        ram_buffer(7344) := X"14800002";
        ram_buffer(7345) := X"0044001A";
        ram_buffer(7346) := X"0007000D";
        ram_buffer(7347) := X"00001012";
        ram_buffer(7348) := X"03E00008";
        ram_buffer(7349) := X"00000000";
        ram_buffer(7350) := X"24020064";
        ram_buffer(7351) := X"00442023";
        ram_buffer(7352) := X"03E00008";
        ram_buffer(7353) := X"00041040";
        ram_buffer(7354) := X"27BDFFE0";
        ram_buffer(7355) := X"AFB20018";
        ram_buffer(7356) := X"AFB10014";
        ram_buffer(7357) := X"AFBF001C";
        ram_buffer(7358) := X"AFB00010";
        ram_buffer(7359) := X"00808821";
        ram_buffer(7360) := X"18A000A2";
        ram_buffer(7361) := X"00C09021";
        ram_buffer(7362) := X"28A20065";
        ram_buffer(7363) := X"144000A1";
        ram_buffer(7364) := X"00008021";
        ram_buffer(7365) := X"8E220010";
        ram_buffer(7366) := X"24030064";
        ram_buffer(7367) := X"1043000A";
        ram_buffer(7368) := X"24040012";
        ram_buffer(7369) := X"8E230000";
        ram_buffer(7370) := X"00000000";
        ram_buffer(7371) := X"AC620018";
        ram_buffer(7372) := X"8E220000";
        ram_buffer(7373) := X"AC640014";
        ram_buffer(7374) := X"8C420000";
        ram_buffer(7375) := X"00000000";
        ram_buffer(7376) := X"0040F809";
        ram_buffer(7377) := X"02202021";
        ram_buffer(7378) := X"8E220040";
        ram_buffer(7379) := X"00000000";
        ram_buffer(7380) := X"1040009E";
        ram_buffer(7381) := X"00000000";
        ram_buffer(7382) := X"3C04100D";
        ram_buffer(7383) := X"3C06100D";
        ram_buffer(7384) := X"24848774";
        ram_buffer(7385) := X"00402821";
        ram_buffer(7386) := X"16400071";
        ram_buffer(7387) := X"24C68874";
        ram_buffer(7388) := X"24080064";
        ram_buffer(7389) := X"10000007";
        ram_buffer(7390) := X"340A8000";
        ram_buffer(7391) := X"1520004F";
        ram_buffer(7392) := X"00000000";
        ram_buffer(7393) := X"24840004";
        ram_buffer(7394) := X"A4A70000";
        ram_buffer(7395) := X"10860012";
        ram_buffer(7396) := X"24A50002";
        ram_buffer(7397) := X"8C830000";
        ram_buffer(7398) := X"24077FFF";
        ram_buffer(7399) := X"02030018";
        ram_buffer(7400) := X"00001812";
        ram_buffer(7401) := X"24630032";
        ram_buffer(7402) := X"00000000";
        ram_buffer(7403) := X"15000002";
        ram_buffer(7404) := X"0068001A";
        ram_buffer(7405) := X"0007000D";
        ram_buffer(7406) := X"00001812";
        ram_buffer(7407) := X"1C60FFEF";
        ram_buffer(7408) := X"006A482A";
        ram_buffer(7409) := X"24070001";
        ram_buffer(7410) := X"24840004";
        ram_buffer(7411) := X"A4A70000";
        ram_buffer(7412) := X"1486FFF0";
        ram_buffer(7413) := X"24A50002";
        ram_buffer(7414) := X"8E230010";
        ram_buffer(7415) := X"AC400080";
        ram_buffer(7416) := X"24020064";
        ram_buffer(7417) := X"1062000A";
        ram_buffer(7418) := X"24040012";
        ram_buffer(7419) := X"8E220000";
        ram_buffer(7420) := X"00000000";
        ram_buffer(7421) := X"AC430018";
        ram_buffer(7422) := X"8E230000";
        ram_buffer(7423) := X"AC440014";
        ram_buffer(7424) := X"8C620000";
        ram_buffer(7425) := X"00000000";
        ram_buffer(7426) := X"0040F809";
        ram_buffer(7427) := X"02202021";
        ram_buffer(7428) := X"8E220044";
        ram_buffer(7429) := X"00000000";
        ram_buffer(7430) := X"10400070";
        ram_buffer(7431) := X"00000000";
        ram_buffer(7432) := X"3C04100D";
        ram_buffer(7433) := X"24848674";
        ram_buffer(7434) := X"16400028";
        ram_buffer(7435) := X"00402821";
        ram_buffer(7436) := X"3C09100D";
        ram_buffer(7437) := X"25298774";
        ram_buffer(7438) := X"24070064";
        ram_buffer(7439) := X"10000007";
        ram_buffer(7440) := X"340A8000";
        ram_buffer(7441) := X"1500001F";
        ram_buffer(7442) := X"00000000";
        ram_buffer(7443) := X"24840004";
        ram_buffer(7444) := X"A4A60000";
        ram_buffer(7445) := X"11240012";
        ram_buffer(7446) := X"24A50002";
        ram_buffer(7447) := X"8C830000";
        ram_buffer(7448) := X"24067FFF";
        ram_buffer(7449) := X"02030018";
        ram_buffer(7450) := X"00001812";
        ram_buffer(7451) := X"24630032";
        ram_buffer(7452) := X"00000000";
        ram_buffer(7453) := X"14E00002";
        ram_buffer(7454) := X"0067001A";
        ram_buffer(7455) := X"0007000D";
        ram_buffer(7456) := X"00001812";
        ram_buffer(7457) := X"1C60FFEF";
        ram_buffer(7458) := X"006A402A";
        ram_buffer(7459) := X"24060001";
        ram_buffer(7460) := X"24840004";
        ram_buffer(7461) := X"A4A60000";
        ram_buffer(7462) := X"1524FFF0";
        ram_buffer(7463) := X"24A50002";
        ram_buffer(7464) := X"8FBF001C";
        ram_buffer(7465) := X"8FB20018";
        ram_buffer(7466) := X"8FB10014";
        ram_buffer(7467) := X"8FB00010";
        ram_buffer(7468) := X"AC400080";
        ram_buffer(7469) := X"03E00008";
        ram_buffer(7470) := X"27BD0020";
        ram_buffer(7471) := X"1000FFB1";
        ram_buffer(7472) := X"3067FFFF";
        ram_buffer(7473) := X"1000FFE1";
        ram_buffer(7474) := X"3066FFFF";
        ram_buffer(7475) := X"3C08100D";
        ram_buffer(7476) := X"25088774";
        ram_buffer(7477) := X"10000008";
        ram_buffer(7478) := X"24060064";
        ram_buffer(7479) := X"10E00043";
        ram_buffer(7480) := X"00000000";
        ram_buffer(7481) := X"3063FFFF";
        ram_buffer(7482) := X"24840004";
        ram_buffer(7483) := X"A4A30000";
        ram_buffer(7484) := X"1088FFEB";
        ram_buffer(7485) := X"24A50002";
        ram_buffer(7486) := X"8C830000";
        ram_buffer(7487) := X"00000000";
        ram_buffer(7488) := X"02030018";
        ram_buffer(7489) := X"00001812";
        ram_buffer(7490) := X"24630032";
        ram_buffer(7491) := X"00000000";
        ram_buffer(7492) := X"14C00002";
        ram_buffer(7493) := X"0066001A";
        ram_buffer(7494) := X"0007000D";
        ram_buffer(7495) := X"00001812";
        ram_buffer(7496) := X"1C60FFEE";
        ram_buffer(7497) := X"28670100";
        ram_buffer(7498) := X"1000FFEF";
        ram_buffer(7499) := X"24030001";
        ram_buffer(7500) := X"10000008";
        ram_buffer(7501) := X"24070064";
        ram_buffer(7502) := X"1100002E";
        ram_buffer(7503) := X"00000000";
        ram_buffer(7504) := X"3063FFFF";
        ram_buffer(7505) := X"24840004";
        ram_buffer(7506) := X"A4A30000";
        ram_buffer(7507) := X"10C4FFA2";
        ram_buffer(7508) := X"24A50002";
        ram_buffer(7509) := X"8C830000";
        ram_buffer(7510) := X"00000000";
        ram_buffer(7511) := X"02030018";
        ram_buffer(7512) := X"00001812";
        ram_buffer(7513) := X"24630032";
        ram_buffer(7514) := X"00000000";
        ram_buffer(7515) := X"14E00002";
        ram_buffer(7516) := X"0067001A";
        ram_buffer(7517) := X"0007000D";
        ram_buffer(7518) := X"00001812";
        ram_buffer(7519) := X"1C60FFEE";
        ram_buffer(7520) := X"28680100";
        ram_buffer(7521) := X"1000FFEF";
        ram_buffer(7522) := X"24030001";
        ram_buffer(7523) := X"1000FF61";
        ram_buffer(7524) := X"24101388";
        ram_buffer(7525) := X"28A20032";
        ram_buffer(7526) := X"10400008";
        ram_buffer(7527) := X"00000000";
        ram_buffer(7528) := X"24101388";
        ram_buffer(7529) := X"14A00002";
        ram_buffer(7530) := X"0205001A";
        ram_buffer(7531) := X"0007000D";
        ram_buffer(7532) := X"00008012";
        ram_buffer(7533) := X"1000FF57";
        ram_buffer(7534) := X"00000000";
        ram_buffer(7535) := X"24100064";
        ram_buffer(7536) := X"02058023";
        ram_buffer(7537) := X"1000FF53";
        ram_buffer(7538) := X"00108040";
        ram_buffer(7539) := X"0C026495";
        ram_buffer(7540) := X"02202021";
        ram_buffer(7541) := X"1000FF60";
        ram_buffer(7542) := X"AE220040";
        ram_buffer(7543) := X"0C026495";
        ram_buffer(7544) := X"02202021";
        ram_buffer(7545) := X"1000FF8E";
        ram_buffer(7546) := X"AE220044";
        ram_buffer(7547) := X"1000FFBE";
        ram_buffer(7548) := X"240300FF";
        ram_buffer(7549) := X"1000FFD3";
        ram_buffer(7550) := X"240300FF";
        ram_buffer(7551) := X"8C820024";
        ram_buffer(7552) := X"27BDFFE8";
        ram_buffer(7553) := X"2C430006";
        ram_buffer(7554) := X"AFB00010";
        ram_buffer(7555) := X"AFBF0014";
        ram_buffer(7556) := X"106000DD";
        ram_buffer(7557) := X"00808021";
        ram_buffer(7558) := X"00021880";
        ram_buffer(7559) := X"3C02100D";
        ram_buffer(7560) := X"2442847C";
        ram_buffer(7561) := X"00431021";
        ram_buffer(7562) := X"8C420000";
        ram_buffer(7563) := X"00000000";
        ram_buffer(7564) := X"00400008";
        ram_buffer(7565) := X"00000000";
        ram_buffer(7566) := X"8C820010";
        ram_buffer(7567) := X"24030064";
        ram_buffer(7568) := X"1043000A";
        ram_buffer(7569) := X"00000000";
        ram_buffer(7570) := X"8C830000";
        ram_buffer(7571) := X"00000000";
        ram_buffer(7572) := X"AC620018";
        ram_buffer(7573) := X"8C820000";
        ram_buffer(7574) := X"24040012";
        ram_buffer(7575) := X"8C420000";
        ram_buffer(7576) := X"AC640014";
        ram_buffer(7577) := X"0040F809";
        ram_buffer(7578) := X"02002021";
        ram_buffer(7579) := X"8E02003C";
        ram_buffer(7580) := X"24030001";
        ram_buffer(7581) := X"24040003";
        ram_buffer(7582) := X"24050002";
        ram_buffer(7583) := X"AE040038";
        ram_buffer(7584) := X"AE0000D4";
        ram_buffer(7585) := X"AE0300C8";
        ram_buffer(7586) := X"AE040034";
        ram_buffer(7587) := X"AC430000";
        ram_buffer(7588) := X"AC450008";
        ram_buffer(7589) := X"AC45000C";
        ram_buffer(7590) := X"AC400010";
        ram_buffer(7591) := X"AC400014";
        ram_buffer(7592) := X"AC400018";
        ram_buffer(7593) := X"AC450054";
        ram_buffer(7594) := X"AC43005C";
        ram_buffer(7595) := X"AC430060";
        ram_buffer(7596) := X"AC430064";
        ram_buffer(7597) := X"AC430068";
        ram_buffer(7598) := X"AC43006C";
        ram_buffer(7599) := X"AC4400A8";
        ram_buffer(7600) := X"AC4300B0";
        ram_buffer(7601) := X"AC4300B4";
        ram_buffer(7602) := X"AC4300B8";
        ram_buffer(7603) := X"AC4300BC";
        ram_buffer(7604) := X"AC4300C0";
        ram_buffer(7605) := X"8FBF0014";
        ram_buffer(7606) := X"8FB00010";
        ram_buffer(7607) := X"03E00008";
        ram_buffer(7608) := X"27BD0018";
        ram_buffer(7609) := X"8C820010";
        ram_buffer(7610) := X"24030064";
        ram_buffer(7611) := X"1043000A";
        ram_buffer(7612) := X"00000000";
        ram_buffer(7613) := X"8C830000";
        ram_buffer(7614) := X"00000000";
        ram_buffer(7615) := X"AC620018";
        ram_buffer(7616) := X"8C820000";
        ram_buffer(7617) := X"24040012";
        ram_buffer(7618) := X"8C420000";
        ram_buffer(7619) := X"AC640014";
        ram_buffer(7620) := X"0040F809";
        ram_buffer(7621) := X"02002021";
        ram_buffer(7622) := X"8E02003C";
        ram_buffer(7623) := X"24060005";
        ram_buffer(7624) := X"8FBF0014";
        ram_buffer(7625) := X"AE060038";
        ram_buffer(7626) := X"24030001";
        ram_buffer(7627) := X"24040002";
        ram_buffer(7628) := X"24050004";
        ram_buffer(7629) := X"24060003";
        ram_buffer(7630) := X"AE0000C8";
        ram_buffer(7631) := X"AE0300D4";
        ram_buffer(7632) := X"AE050034";
        ram_buffer(7633) := X"8FB00010";
        ram_buffer(7634) := X"AC430000";
        ram_buffer(7635) := X"AC440008";
        ram_buffer(7636) := X"AC44000C";
        ram_buffer(7637) := X"AC400010";
        ram_buffer(7638) := X"AC400014";
        ram_buffer(7639) := X"AC400018";
        ram_buffer(7640) := X"AC440054";
        ram_buffer(7641) := X"AC43005C";
        ram_buffer(7642) := X"AC430060";
        ram_buffer(7643) := X"AC430064";
        ram_buffer(7644) := X"AC430068";
        ram_buffer(7645) := X"AC43006C";
        ram_buffer(7646) := X"AC4600A8";
        ram_buffer(7647) := X"AC4300B0";
        ram_buffer(7648) := X"AC4300B4";
        ram_buffer(7649) := X"AC4300B8";
        ram_buffer(7650) := X"AC4300BC";
        ram_buffer(7651) := X"AC4300C0";
        ram_buffer(7652) := X"AC4500FC";
        ram_buffer(7653) := X"AC440104";
        ram_buffer(7654) := X"AC440108";
        ram_buffer(7655) := X"AC40010C";
        ram_buffer(7656) := X"AC400110";
        ram_buffer(7657) := X"AC400114";
        ram_buffer(7658) := X"03E00008";
        ram_buffer(7659) := X"27BD0018";
        ram_buffer(7660) := X"8C820010";
        ram_buffer(7661) := X"24030064";
        ram_buffer(7662) := X"1043000A";
        ram_buffer(7663) := X"00000000";
        ram_buffer(7664) := X"8C830000";
        ram_buffer(7665) := X"00000000";
        ram_buffer(7666) := X"AC620018";
        ram_buffer(7667) := X"8C820000";
        ram_buffer(7668) := X"24040012";
        ram_buffer(7669) := X"8C420000";
        ram_buffer(7670) := X"AC640014";
        ram_buffer(7671) := X"0040F809";
        ram_buffer(7672) := X"02002021";
        ram_buffer(7673) := X"8E050020";
        ram_buffer(7674) := X"AE000038";
        ram_buffer(7675) := X"24A2FFFF";
        ram_buffer(7676) := X"2C42000A";
        ram_buffer(7677) := X"AE0000C8";
        ram_buffer(7678) := X"AE0000D4";
        ram_buffer(7679) := X"1040006A";
        ram_buffer(7680) := X"AE050034";
        ram_buffer(7681) := X"8E02003C";
        ram_buffer(7682) := X"00001821";
        ram_buffer(7683) := X"24040001";
        ram_buffer(7684) := X"AC430000";
        ram_buffer(7685) := X"24630001";
        ram_buffer(7686) := X"AC440008";
        ram_buffer(7687) := X"AC44000C";
        ram_buffer(7688) := X"AC400010";
        ram_buffer(7689) := X"AC400014";
        ram_buffer(7690) := X"AC400018";
        ram_buffer(7691) := X"1465FFF8";
        ram_buffer(7692) := X"24420054";
        ram_buffer(7693) := X"8FBF0014";
        ram_buffer(7694) := X"8FB00010";
        ram_buffer(7695) := X"03E00008";
        ram_buffer(7696) := X"27BD0018";
        ram_buffer(7697) := X"8C820010";
        ram_buffer(7698) := X"24030064";
        ram_buffer(7699) := X"1043000A";
        ram_buffer(7700) := X"00000000";
        ram_buffer(7701) := X"8C830000";
        ram_buffer(7702) := X"00000000";
        ram_buffer(7703) := X"AC620018";
        ram_buffer(7704) := X"8C820000";
        ram_buffer(7705) := X"24040012";
        ram_buffer(7706) := X"8C420000";
        ram_buffer(7707) := X"AC640014";
        ram_buffer(7708) := X"0040F809";
        ram_buffer(7709) := X"02002021";
        ram_buffer(7710) := X"8E02003C";
        ram_buffer(7711) := X"8FBF0014";
        ram_buffer(7712) := X"24030001";
        ram_buffer(7713) := X"AE030038";
        ram_buffer(7714) := X"AE0000D4";
        ram_buffer(7715) := X"AE0300C8";
        ram_buffer(7716) := X"AE030034";
        ram_buffer(7717) := X"8FB00010";
        ram_buffer(7718) := X"AC430000";
        ram_buffer(7719) := X"AC430008";
        ram_buffer(7720) := X"AC43000C";
        ram_buffer(7721) := X"AC400010";
        ram_buffer(7722) := X"AC400014";
        ram_buffer(7723) := X"AC400018";
        ram_buffer(7724) := X"03E00008";
        ram_buffer(7725) := X"27BD0018";
        ram_buffer(7726) := X"8C820010";
        ram_buffer(7727) := X"24030064";
        ram_buffer(7728) := X"1043000A";
        ram_buffer(7729) := X"00000000";
        ram_buffer(7730) := X"8C830000";
        ram_buffer(7731) := X"00000000";
        ram_buffer(7732) := X"AC620018";
        ram_buffer(7733) := X"8C820000";
        ram_buffer(7734) := X"24040012";
        ram_buffer(7735) := X"8C420000";
        ram_buffer(7736) := X"AC640014";
        ram_buffer(7737) := X"0040F809";
        ram_buffer(7738) := X"02002021";
        ram_buffer(7739) := X"8E02003C";
        ram_buffer(7740) := X"24040004";
        ram_buffer(7741) := X"AE040038";
        ram_buffer(7742) := X"AE040034";
        ram_buffer(7743) := X"24030001";
        ram_buffer(7744) := X"24040043";
        ram_buffer(7745) := X"AE0000C8";
        ram_buffer(7746) := X"AE0300D4";
        ram_buffer(7747) := X"AC440000";
        ram_buffer(7748) := X"2404004D";
        ram_buffer(7749) := X"AC440054";
        ram_buffer(7750) := X"8FBF0014";
        ram_buffer(7751) := X"24040059";
        ram_buffer(7752) := X"AC4400A8";
        ram_buffer(7753) := X"2404004B";
        ram_buffer(7754) := X"8FB00010";
        ram_buffer(7755) := X"AC430008";
        ram_buffer(7756) := X"AC43000C";
        ram_buffer(7757) := X"AC400010";
        ram_buffer(7758) := X"AC400014";
        ram_buffer(7759) := X"AC400018";
        ram_buffer(7760) := X"AC43005C";
        ram_buffer(7761) := X"AC430060";
        ram_buffer(7762) := X"AC400064";
        ram_buffer(7763) := X"AC400068";
        ram_buffer(7764) := X"AC40006C";
        ram_buffer(7765) := X"AC4300B0";
        ram_buffer(7766) := X"AC4300B4";
        ram_buffer(7767) := X"AC4000B8";
        ram_buffer(7768) := X"AC4000BC";
        ram_buffer(7769) := X"AC4000C0";
        ram_buffer(7770) := X"AC4400FC";
        ram_buffer(7771) := X"AC430104";
        ram_buffer(7772) := X"AC430108";
        ram_buffer(7773) := X"AC40010C";
        ram_buffer(7774) := X"AC400110";
        ram_buffer(7775) := X"AC400114";
        ram_buffer(7776) := X"03E00008";
        ram_buffer(7777) := X"27BD0018";
        ram_buffer(7778) := X"8C820000";
        ram_buffer(7779) := X"8FBF0014";
        ram_buffer(7780) := X"8FB00010";
        ram_buffer(7781) := X"8C590000";
        ram_buffer(7782) := X"24030007";
        ram_buffer(7783) := X"AC430014";
        ram_buffer(7784) := X"03200008";
        ram_buffer(7785) := X"27BD0018";
        ram_buffer(7786) := X"8E020000";
        ram_buffer(7787) := X"24040018";
        ram_buffer(7788) := X"AC450018";
        ram_buffer(7789) := X"8E030000";
        ram_buffer(7790) := X"AC440014";
        ram_buffer(7791) := X"2402000A";
        ram_buffer(7792) := X"AC62001C";
        ram_buffer(7793) := X"8E020000";
        ram_buffer(7794) := X"00000000";
        ram_buffer(7795) := X"8C420000";
        ram_buffer(7796) := X"00000000";
        ram_buffer(7797) := X"0040F809";
        ram_buffer(7798) := X"02002021";
        ram_buffer(7799) := X"8E050034";
        ram_buffer(7800) := X"00000000";
        ram_buffer(7801) := X"1CA0FF87";
        ram_buffer(7802) := X"00000000";
        ram_buffer(7803) := X"1000FF39";
        ram_buffer(7804) := X"00000000";
        ram_buffer(7805) := X"8C820010";
        ram_buffer(7806) := X"27BDFFE0";
        ram_buffer(7807) := X"24030064";
        ram_buffer(7808) := X"AFB10018";
        ram_buffer(7809) := X"AFB00014";
        ram_buffer(7810) := X"AFBF001C";
        ram_buffer(7811) := X"00808021";
        ram_buffer(7812) := X"1043000A";
        ram_buffer(7813) := X"00A08821";
        ram_buffer(7814) := X"8C830000";
        ram_buffer(7815) := X"24050012";
        ram_buffer(7816) := X"AC620018";
        ram_buffer(7817) := X"8C820000";
        ram_buffer(7818) := X"AC650014";
        ram_buffer(7819) := X"8C420000";
        ram_buffer(7820) := X"00000000";
        ram_buffer(7821) := X"0040F809";
        ram_buffer(7822) := X"00000000";
        ram_buffer(7823) := X"2E220006";
        ram_buffer(7824) := X"AE110038";
        ram_buffer(7825) := X"AE0000C8";
        ram_buffer(7826) := X"104000B5";
        ram_buffer(7827) := X"AE0000D4";
        ram_buffer(7828) := X"3C05100D";
        ram_buffer(7829) := X"00118880";
        ram_buffer(7830) := X"24A58494";
        ram_buffer(7831) := X"00B18821";
        ram_buffer(7832) := X"8E220000";
        ram_buffer(7833) := X"00000000";
        ram_buffer(7834) := X"00400008";
        ram_buffer(7835) := X"00000000";
        ram_buffer(7836) := X"8E02003C";
        ram_buffer(7837) := X"24040004";
        ram_buffer(7838) := X"AE040034";
        ram_buffer(7839) := X"24030001";
        ram_buffer(7840) := X"24040043";
        ram_buffer(7841) := X"AE0300D4";
        ram_buffer(7842) := X"AC440000";
        ram_buffer(7843) := X"2404004D";
        ram_buffer(7844) := X"AC440054";
        ram_buffer(7845) := X"24040059";
        ram_buffer(7846) := X"AC4400A8";
        ram_buffer(7847) := X"2404004B";
        ram_buffer(7848) := X"AC430008";
        ram_buffer(7849) := X"AC43000C";
        ram_buffer(7850) := X"AC400010";
        ram_buffer(7851) := X"AC400014";
        ram_buffer(7852) := X"AC400018";
        ram_buffer(7853) := X"AC43005C";
        ram_buffer(7854) := X"AC430060";
        ram_buffer(7855) := X"AC400064";
        ram_buffer(7856) := X"AC400068";
        ram_buffer(7857) := X"AC40006C";
        ram_buffer(7858) := X"AC4300B0";
        ram_buffer(7859) := X"AC4300B4";
        ram_buffer(7860) := X"AC4000B8";
        ram_buffer(7861) := X"AC4000BC";
        ram_buffer(7862) := X"AC4000C0";
        ram_buffer(7863) := X"AC4400FC";
        ram_buffer(7864) := X"AC430104";
        ram_buffer(7865) := X"AC430108";
        ram_buffer(7866) := X"AC40010C";
        ram_buffer(7867) := X"AC400110";
        ram_buffer(7868) := X"AC400114";
        ram_buffer(7869) := X"8FBF001C";
        ram_buffer(7870) := X"8FB10018";
        ram_buffer(7871) := X"8FB00014";
        ram_buffer(7872) := X"03E00008";
        ram_buffer(7873) := X"27BD0020";
        ram_buffer(7874) := X"8E02003C";
        ram_buffer(7875) := X"8FBF001C";
        ram_buffer(7876) := X"24030001";
        ram_buffer(7877) := X"24040002";
        ram_buffer(7878) := X"24050004";
        ram_buffer(7879) := X"24060003";
        ram_buffer(7880) := X"AE0300D4";
        ram_buffer(7881) := X"AE050034";
        ram_buffer(7882) := X"8FB10018";
        ram_buffer(7883) := X"8FB00014";
        ram_buffer(7884) := X"AC430000";
        ram_buffer(7885) := X"AC440008";
        ram_buffer(7886) := X"AC44000C";
        ram_buffer(7887) := X"AC400010";
        ram_buffer(7888) := X"AC400014";
        ram_buffer(7889) := X"AC400018";
        ram_buffer(7890) := X"AC440054";
        ram_buffer(7891) := X"AC43005C";
        ram_buffer(7892) := X"AC430060";
        ram_buffer(7893) := X"AC430064";
        ram_buffer(7894) := X"AC430068";
        ram_buffer(7895) := X"AC43006C";
        ram_buffer(7896) := X"AC4600A8";
        ram_buffer(7897) := X"AC4300B0";
        ram_buffer(7898) := X"AC4300B4";
        ram_buffer(7899) := X"AC4300B8";
        ram_buffer(7900) := X"AC4300BC";
        ram_buffer(7901) := X"AC4300C0";
        ram_buffer(7902) := X"AC4500FC";
        ram_buffer(7903) := X"AC440104";
        ram_buffer(7904) := X"AC440108";
        ram_buffer(7905) := X"AC40010C";
        ram_buffer(7906) := X"AC400110";
        ram_buffer(7907) := X"AC400114";
        ram_buffer(7908) := X"03E00008";
        ram_buffer(7909) := X"27BD0020";
        ram_buffer(7910) := X"8E050020";
        ram_buffer(7911) := X"00000000";
        ram_buffer(7912) := X"24A2FFFF";
        ram_buffer(7913) := X"2C42000A";
        ram_buffer(7914) := X"10400067";
        ram_buffer(7915) := X"AE050034";
        ram_buffer(7916) := X"8E02003C";
        ram_buffer(7917) := X"00001821";
        ram_buffer(7918) := X"24040001";
        ram_buffer(7919) := X"AC430000";
        ram_buffer(7920) := X"24630001";
        ram_buffer(7921) := X"AC440008";
        ram_buffer(7922) := X"AC44000C";
        ram_buffer(7923) := X"AC400010";
        ram_buffer(7924) := X"AC400014";
        ram_buffer(7925) := X"AC400018";
        ram_buffer(7926) := X"1465FFF8";
        ram_buffer(7927) := X"24420054";
        ram_buffer(7928) := X"8FBF001C";
        ram_buffer(7929) := X"8FB10018";
        ram_buffer(7930) := X"8FB00014";
        ram_buffer(7931) := X"03E00008";
        ram_buffer(7932) := X"27BD0020";
        ram_buffer(7933) := X"8E02003C";
        ram_buffer(7934) := X"8FBF001C";
        ram_buffer(7935) := X"24030001";
        ram_buffer(7936) := X"AE0300C8";
        ram_buffer(7937) := X"AE030034";
        ram_buffer(7938) := X"8FB10018";
        ram_buffer(7939) := X"8FB00014";
        ram_buffer(7940) := X"AC430000";
        ram_buffer(7941) := X"AC430008";
        ram_buffer(7942) := X"AC43000C";
        ram_buffer(7943) := X"AC400010";
        ram_buffer(7944) := X"AC400014";
        ram_buffer(7945) := X"AC400018";
        ram_buffer(7946) := X"03E00008";
        ram_buffer(7947) := X"27BD0020";
        ram_buffer(7948) := X"8E02003C";
        ram_buffer(7949) := X"24040003";
        ram_buffer(7950) := X"AE040034";
        ram_buffer(7951) := X"24030001";
        ram_buffer(7952) := X"24040052";
        ram_buffer(7953) := X"AE0300D4";
        ram_buffer(7954) := X"8FBF001C";
        ram_buffer(7955) := X"AC440000";
        ram_buffer(7956) := X"24040047";
        ram_buffer(7957) := X"AC440054";
        ram_buffer(7958) := X"24040042";
        ram_buffer(7959) := X"8FB10018";
        ram_buffer(7960) := X"8FB00014";
        ram_buffer(7961) := X"AC430008";
        ram_buffer(7962) := X"AC43000C";
        ram_buffer(7963) := X"AC400010";
        ram_buffer(7964) := X"AC400014";
        ram_buffer(7965) := X"AC400018";
        ram_buffer(7966) := X"AC43005C";
        ram_buffer(7967) := X"AC430060";
        ram_buffer(7968) := X"AC400064";
        ram_buffer(7969) := X"AC400068";
        ram_buffer(7970) := X"AC40006C";
        ram_buffer(7971) := X"AC4400A8";
        ram_buffer(7972) := X"AC4300B0";
        ram_buffer(7973) := X"AC4300B4";
        ram_buffer(7974) := X"AC4000B8";
        ram_buffer(7975) := X"AC4000BC";
        ram_buffer(7976) := X"AC4000C0";
        ram_buffer(7977) := X"03E00008";
        ram_buffer(7978) := X"27BD0020";
        ram_buffer(7979) := X"8E02003C";
        ram_buffer(7980) := X"8FBF001C";
        ram_buffer(7981) := X"24030001";
        ram_buffer(7982) := X"24040002";
        ram_buffer(7983) := X"24050003";
        ram_buffer(7984) := X"AE0300C8";
        ram_buffer(7985) := X"AE050034";
        ram_buffer(7986) := X"8FB10018";
        ram_buffer(7987) := X"8FB00014";
        ram_buffer(7988) := X"AC430000";
        ram_buffer(7989) := X"AC440008";
        ram_buffer(7990) := X"AC44000C";
        ram_buffer(7991) := X"AC400010";
        ram_buffer(7992) := X"AC400014";
        ram_buffer(7993) := X"AC400018";
        ram_buffer(7994) := X"AC440054";
        ram_buffer(7995) := X"AC43005C";
        ram_buffer(7996) := X"AC430060";
        ram_buffer(7997) := X"AC430064";
        ram_buffer(7998) := X"AC430068";
        ram_buffer(7999) := X"AC43006C";
        ram_buffer(8000) := X"AC4500A8";
        ram_buffer(8001) := X"AC4300B0";
        ram_buffer(8002) := X"AC4300B4";
        ram_buffer(8003) := X"AC4300B8";
        ram_buffer(8004) := X"AC4300BC";
        ram_buffer(8005) := X"AC4300C0";
        ram_buffer(8006) := X"03E00008";
        ram_buffer(8007) := X"27BD0020";
        ram_buffer(8008) := X"8E020000";
        ram_buffer(8009) := X"8FBF001C";
        ram_buffer(8010) := X"8FB10018";
        ram_buffer(8011) := X"8C590000";
        ram_buffer(8012) := X"24030008";
        ram_buffer(8013) := X"02002021";
        ram_buffer(8014) := X"8FB00014";
        ram_buffer(8015) := X"AC430014";
        ram_buffer(8016) := X"03200008";
        ram_buffer(8017) := X"27BD0020";
        ram_buffer(8018) := X"8E020000";
        ram_buffer(8019) := X"24040018";
        ram_buffer(8020) := X"AC450018";
        ram_buffer(8021) := X"8E030000";
        ram_buffer(8022) := X"AC440014";
        ram_buffer(8023) := X"2402000A";
        ram_buffer(8024) := X"AC62001C";
        ram_buffer(8025) := X"8E020000";
        ram_buffer(8026) := X"00000000";
        ram_buffer(8027) := X"8C420000";
        ram_buffer(8028) := X"00000000";
        ram_buffer(8029) := X"0040F809";
        ram_buffer(8030) := X"02002021";
        ram_buffer(8031) := X"8E050034";
        ram_buffer(8032) := X"00000000";
        ram_buffer(8033) := X"1CA0FF8A";
        ram_buffer(8034) := X"00000000";
        ram_buffer(8035) := X"1000FF59";
        ram_buffer(8036) := X"00000000";
        ram_buffer(8037) := X"8C820010";
        ram_buffer(8038) := X"27BDFFE8";
        ram_buffer(8039) := X"24030064";
        ram_buffer(8040) := X"AFB00010";
        ram_buffer(8041) := X"AFBF0014";
        ram_buffer(8042) := X"1043000A";
        ram_buffer(8043) := X"00808021";
        ram_buffer(8044) := X"8C830000";
        ram_buffer(8045) := X"24050012";
        ram_buffer(8046) := X"AC620018";
        ram_buffer(8047) := X"8C820000";
        ram_buffer(8048) := X"AC650014";
        ram_buffer(8049) := X"8C420000";
        ram_buffer(8050) := X"00000000";
        ram_buffer(8051) := X"0040F809";
        ram_buffer(8052) := X"00000000";
        ram_buffer(8053) := X"8E02003C";
        ram_buffer(8054) := X"00000000";
        ram_buffer(8055) := X"10400159";
        ram_buffer(8056) := X"24060348";
        ram_buffer(8057) := X"24030008";
        ram_buffer(8058) := X"8E020010";
        ram_buffer(8059) := X"AE030030";
        ram_buffer(8060) := X"24030064";
        ram_buffer(8061) := X"1043000A";
        ram_buffer(8062) := X"24040012";
        ram_buffer(8063) := X"8E030000";
        ram_buffer(8064) := X"00000000";
        ram_buffer(8065) := X"AC620018";
        ram_buffer(8066) := X"8E020000";
        ram_buffer(8067) := X"AC640014";
        ram_buffer(8068) := X"8C420000";
        ram_buffer(8069) := X"00000000";
        ram_buffer(8070) := X"0040F809";
        ram_buffer(8071) := X"02002021";
        ram_buffer(8072) := X"8E020040";
        ram_buffer(8073) := X"00000000";
        ram_buffer(8074) := X"1040014E";
        ram_buffer(8075) := X"00000000";
        ram_buffer(8076) := X"3C05100D";
        ram_buffer(8077) := X"3C08100D";
        ram_buffer(8078) := X"24A58774";
        ram_buffer(8079) := X"00403021";
        ram_buffer(8080) := X"25088874";
        ram_buffer(8081) := X"24070064";
        ram_buffer(8082) := X"1000000C";
        ram_buffer(8083) := X"34098000";
        ram_buffer(8084) := X"2464FFFF";
        ram_buffer(8085) := X"2C847FFF";
        ram_buffer(8086) := X"108000BB";
        ram_buffer(8087) := X"28640100";
        ram_buffer(8088) := X"14800002";
        ram_buffer(8089) := X"00000000";
        ram_buffer(8090) := X"240300FF";
        ram_buffer(8091) := X"24A50004";
        ram_buffer(8092) := X"A4C30000";
        ram_buffer(8093) := X"10A80015";
        ram_buffer(8094) := X"24C60002";
        ram_buffer(8095) := X"8CA30000";
        ram_buffer(8096) := X"00000000";
        ram_buffer(8097) := X"00032040";
        ram_buffer(8098) := X"000318C0";
        ram_buffer(8099) := X"00831821";
        ram_buffer(8100) := X"00032080";
        ram_buffer(8101) := X"00641821";
        ram_buffer(8102) := X"24630032";
        ram_buffer(8103) := X"14E00002";
        ram_buffer(8104) := X"0067001A";
        ram_buffer(8105) := X"0007000D";
        ram_buffer(8106) := X"00001812";
        ram_buffer(8107) := X"0069202A";
        ram_buffer(8108) := X"1480FFE7";
        ram_buffer(8109) := X"00000000";
        ram_buffer(8110) := X"240300FF";
        ram_buffer(8111) := X"24A50004";
        ram_buffer(8112) := X"A4C30000";
        ram_buffer(8113) := X"14A8FFED";
        ram_buffer(8114) := X"24C60002";
        ram_buffer(8115) := X"8E030010";
        ram_buffer(8116) := X"AC400080";
        ram_buffer(8117) := X"24020064";
        ram_buffer(8118) := X"1062000A";
        ram_buffer(8119) := X"24040012";
        ram_buffer(8120) := X"8E020000";
        ram_buffer(8121) := X"00000000";
        ram_buffer(8122) := X"AC430018";
        ram_buffer(8123) := X"8E030000";
        ram_buffer(8124) := X"AC440014";
        ram_buffer(8125) := X"8C620000";
        ram_buffer(8126) := X"00000000";
        ram_buffer(8127) := X"0040F809";
        ram_buffer(8128) := X"02002021";
        ram_buffer(8129) := X"8E020044";
        ram_buffer(8130) := X"00000000";
        ram_buffer(8131) := X"10400109";
        ram_buffer(8132) := X"00000000";
        ram_buffer(8133) := X"3C05100D";
        ram_buffer(8134) := X"3C08100D";
        ram_buffer(8135) := X"24A58674";
        ram_buffer(8136) := X"00403021";
        ram_buffer(8137) := X"25088774";
        ram_buffer(8138) := X"24070064";
        ram_buffer(8139) := X"1000000B";
        ram_buffer(8140) := X"34098000";
        ram_buffer(8141) := X"2C847FFF";
        ram_buffer(8142) := X"10800085";
        ram_buffer(8143) := X"28640100";
        ram_buffer(8144) := X"14800002";
        ram_buffer(8145) := X"00000000";
        ram_buffer(8146) := X"240300FF";
        ram_buffer(8147) := X"24A50004";
        ram_buffer(8148) := X"A4C30000";
        ram_buffer(8149) := X"11050015";
        ram_buffer(8150) := X"24C60002";
        ram_buffer(8151) := X"8CA30000";
        ram_buffer(8152) := X"00000000";
        ram_buffer(8153) := X"00032040";
        ram_buffer(8154) := X"000318C0";
        ram_buffer(8155) := X"00831821";
        ram_buffer(8156) := X"00032080";
        ram_buffer(8157) := X"00641821";
        ram_buffer(8158) := X"24630032";
        ram_buffer(8159) := X"14E00002";
        ram_buffer(8160) := X"0067001A";
        ram_buffer(8161) := X"0007000D";
        ram_buffer(8162) := X"00001812";
        ram_buffer(8163) := X"0069202A";
        ram_buffer(8164) := X"1480FFE8";
        ram_buffer(8165) := X"2464FFFF";
        ram_buffer(8166) := X"240300FF";
        ram_buffer(8167) := X"24A50004";
        ram_buffer(8168) := X"A4C30000";
        ram_buffer(8169) := X"1505FFED";
        ram_buffer(8170) := X"24C60002";
        ram_buffer(8171) := X"8E040050";
        ram_buffer(8172) := X"00000000";
        ram_buffer(8173) := X"108000DA";
        ram_buffer(8174) := X"AC400080";
        ram_buffer(8175) := X"3C05100D";
        ram_buffer(8176) := X"24060011";
        ram_buffer(8177) := X"0C027F93";
        ram_buffer(8178) := X"24A58660";
        ram_buffer(8179) := X"8E040050";
        ram_buffer(8180) := X"3C05100D";
        ram_buffer(8181) := X"24840011";
        ram_buffer(8182) := X"24060100";
        ram_buffer(8183) := X"0C027F93";
        ram_buffer(8184) := X"24A58654";
        ram_buffer(8185) := X"8E020050";
        ram_buffer(8186) := X"8E040060";
        ram_buffer(8187) := X"00000000";
        ram_buffer(8188) := X"108000C1";
        ram_buffer(8189) := X"AC400114";
        ram_buffer(8190) := X"3C05100D";
        ram_buffer(8191) := X"24060011";
        ram_buffer(8192) := X"0C027F93";
        ram_buffer(8193) := X"24A58640";
        ram_buffer(8194) := X"8E040060";
        ram_buffer(8195) := X"3C05100D";
        ram_buffer(8196) := X"24840011";
        ram_buffer(8197) := X"24060100";
        ram_buffer(8198) := X"0C027F93";
        ram_buffer(8199) := X"24A5859C";
        ram_buffer(8200) := X"8E020060";
        ram_buffer(8201) := X"8E040054";
        ram_buffer(8202) := X"00000000";
        ram_buffer(8203) := X"108000B7";
        ram_buffer(8204) := X"AC400114";
        ram_buffer(8205) := X"3C05100D";
        ram_buffer(8206) := X"24060011";
        ram_buffer(8207) := X"0C027F93";
        ram_buffer(8208) := X"24A58588";
        ram_buffer(8209) := X"8E040054";
        ram_buffer(8210) := X"3C05100D";
        ram_buffer(8211) := X"24840011";
        ram_buffer(8212) := X"24060100";
        ram_buffer(8213) := X"0C027F93";
        ram_buffer(8214) := X"24A5857C";
        ram_buffer(8215) := X"8E020054";
        ram_buffer(8216) := X"8E040064";
        ram_buffer(8217) := X"00000000";
        ram_buffer(8218) := X"1080009E";
        ram_buffer(8219) := X"AC400114";
        ram_buffer(8220) := X"3C05100D";
        ram_buffer(8221) := X"24060011";
        ram_buffer(8222) := X"0C027F93";
        ram_buffer(8223) := X"24A58568";
        ram_buffer(8224) := X"8E040064";
        ram_buffer(8225) := X"3C05100D";
        ram_buffer(8226) := X"24060100";
        ram_buffer(8227) := X"24A584C4";
        ram_buffer(8228) := X"0C027F93";
        ram_buffer(8229) := X"24840011";
        ram_buffer(8230) := X"8E020064";
        ram_buffer(8231) := X"24060010";
        ram_buffer(8232) := X"00002821";
        ram_buffer(8233) := X"26040070";
        ram_buffer(8234) := X"0C02801D";
        ram_buffer(8235) := X"AC400114";
        ram_buffer(8236) := X"24060010";
        ram_buffer(8237) := X"24050001";
        ram_buffer(8238) := X"0C02801D";
        ram_buffer(8239) := X"26040080";
        ram_buffer(8240) := X"24060010";
        ram_buffer(8241) := X"24050005";
        ram_buffer(8242) := X"0C02801D";
        ram_buffer(8243) := X"26040090";
        ram_buffer(8244) := X"8E020030";
        ram_buffer(8245) := X"AE0000A4";
        ram_buffer(8246) := X"28420009";
        ram_buffer(8247) := X"AE0000A0";
        ram_buffer(8248) := X"AE0000A8";
        ram_buffer(8249) := X"AE0000AC";
        ram_buffer(8250) := X"14400003";
        ram_buffer(8251) := X"AE0000B0";
        ram_buffer(8252) := X"24020001";
        ram_buffer(8253) := X"AE0200B0";
        ram_buffer(8254) := X"8E020024";
        ram_buffer(8255) := X"24030001";
        ram_buffer(8256) := X"2C440006";
        ram_buffer(8257) := X"AE0000B4";
        ram_buffer(8258) := X"AE0000B8";
        ram_buffer(8259) := X"AE0000BC";
        ram_buffer(8260) := X"AE0000C0";
        ram_buffer(8261) := X"AE0000C4";
        ram_buffer(8262) := X"A20000CC";
        ram_buffer(8263) := X"A60300CE";
        ram_buffer(8264) := X"10800067";
        ram_buffer(8265) := X"A60300D0";
        ram_buffer(8266) := X"00021880";
        ram_buffer(8267) := X"3C02100D";
        ram_buffer(8268) := X"244284AC";
        ram_buffer(8269) := X"00431021";
        ram_buffer(8270) := X"8C420000";
        ram_buffer(8271) := X"00000000";
        ram_buffer(8272) := X"00400008";
        ram_buffer(8273) := X"00000000";
        ram_buffer(8274) := X"1000FF48";
        ram_buffer(8275) := X"24030001";
        ram_buffer(8276) := X"1000FF7E";
        ram_buffer(8277) := X"24030001";
        ram_buffer(8278) := X"8E020010";
        ram_buffer(8279) := X"24030064";
        ram_buffer(8280) := X"1043000A";
        ram_buffer(8281) := X"24040012";
        ram_buffer(8282) := X"8E030000";
        ram_buffer(8283) := X"00000000";
        ram_buffer(8284) := X"AC620018";
        ram_buffer(8285) := X"8E020000";
        ram_buffer(8286) := X"AC640014";
        ram_buffer(8287) := X"8C420000";
        ram_buffer(8288) := X"00000000";
        ram_buffer(8289) := X"0040F809";
        ram_buffer(8290) := X"02002021";
        ram_buffer(8291) := X"8E02003C";
        ram_buffer(8292) := X"8FBF0014";
        ram_buffer(8293) := X"24030001";
        ram_buffer(8294) := X"24040003";
        ram_buffer(8295) := X"24050002";
        ram_buffer(8296) := X"AE040038";
        ram_buffer(8297) := X"AE0000D4";
        ram_buffer(8298) := X"AE0300C8";
        ram_buffer(8299) := X"AE040034";
        ram_buffer(8300) := X"8FB00010";
        ram_buffer(8301) := X"AC430000";
        ram_buffer(8302) := X"AC450008";
        ram_buffer(8303) := X"AC45000C";
        ram_buffer(8304) := X"AC400010";
        ram_buffer(8305) := X"AC400014";
        ram_buffer(8306) := X"AC400018";
        ram_buffer(8307) := X"AC450054";
        ram_buffer(8308) := X"AC43005C";
        ram_buffer(8309) := X"AC430060";
        ram_buffer(8310) := X"AC430064";
        ram_buffer(8311) := X"AC430068";
        ram_buffer(8312) := X"AC43006C";
        ram_buffer(8313) := X"AC4400A8";
        ram_buffer(8314) := X"AC4300B0";
        ram_buffer(8315) := X"AC4300B4";
        ram_buffer(8316) := X"AC4300B8";
        ram_buffer(8317) := X"AC4300BC";
        ram_buffer(8318) := X"AC4300C0";
        ram_buffer(8319) := X"03E00008";
        ram_buffer(8320) := X"27BD0018";
        ram_buffer(8321) := X"8E020010";
        ram_buffer(8322) := X"24030064";
        ram_buffer(8323) := X"1043000A";
        ram_buffer(8324) := X"00000000";
        ram_buffer(8325) := X"8E030000";
        ram_buffer(8326) := X"24040012";
        ram_buffer(8327) := X"AC620018";
        ram_buffer(8328) := X"8E020000";
        ram_buffer(8329) := X"AC640014";
        ram_buffer(8330) := X"8C420000";
        ram_buffer(8331) := X"00000000";
        ram_buffer(8332) := X"0040F809";
        ram_buffer(8333) := X"02002021";
        ram_buffer(8334) := X"8E02003C";
        ram_buffer(8335) := X"8FBF0014";
        ram_buffer(8336) := X"24030001";
        ram_buffer(8337) := X"AE030038";
        ram_buffer(8338) := X"AE0000D4";
        ram_buffer(8339) := X"AE0300C8";
        ram_buffer(8340) := X"AE030034";
        ram_buffer(8341) := X"8FB00010";
        ram_buffer(8342) := X"AC430000";
        ram_buffer(8343) := X"AC430008";
        ram_buffer(8344) := X"AC43000C";
        ram_buffer(8345) := X"AC400010";
        ram_buffer(8346) := X"AC400014";
        ram_buffer(8347) := X"AC400018";
        ram_buffer(8348) := X"03E00008";
        ram_buffer(8349) := X"27BD0018";
        ram_buffer(8350) := X"8FBF0014";
        ram_buffer(8351) := X"02002021";
        ram_buffer(8352) := X"8FB00010";
        ram_buffer(8353) := X"24050005";
        ram_buffer(8354) := X"08021E7D";
        ram_buffer(8355) := X"27BD0018";
        ram_buffer(8356) := X"8FBF0014";
        ram_buffer(8357) := X"02002021";
        ram_buffer(8358) := X"8FB00010";
        ram_buffer(8359) := X"00002821";
        ram_buffer(8360) := X"08021E7D";
        ram_buffer(8361) := X"27BD0018";
        ram_buffer(8362) := X"8FBF0014";
        ram_buffer(8363) := X"02002021";
        ram_buffer(8364) := X"8FB00010";
        ram_buffer(8365) := X"24050004";
        ram_buffer(8366) := X"08021E7D";
        ram_buffer(8367) := X"27BD0018";
        ram_buffer(8368) := X"8E020000";
        ram_buffer(8369) := X"8FBF0014";
        ram_buffer(8370) := X"8C590000";
        ram_buffer(8371) := X"24030007";
        ram_buffer(8372) := X"02002021";
        ram_buffer(8373) := X"8FB00010";
        ram_buffer(8374) := X"AC430014";
        ram_buffer(8375) := X"03200008";
        ram_buffer(8376) := X"27BD0018";
        ram_buffer(8377) := X"0C0264A0";
        ram_buffer(8378) := X"02002021";
        ram_buffer(8379) := X"00402021";
        ram_buffer(8380) := X"1000FF5F";
        ram_buffer(8381) := X"AE020064";
        ram_buffer(8382) := X"0C0264A0";
        ram_buffer(8383) := X"02002021";
        ram_buffer(8384) := X"00402021";
        ram_buffer(8385) := X"1000FF3C";
        ram_buffer(8386) := X"AE020060";
        ram_buffer(8387) := X"0C0264A0";
        ram_buffer(8388) := X"02002021";
        ram_buffer(8389) := X"00402021";
        ram_buffer(8390) := X"1000FF46";
        ram_buffer(8391) := X"AE020054";
        ram_buffer(8392) := X"0C0264A0";
        ram_buffer(8393) := X"02002021";
        ram_buffer(8394) := X"00402021";
        ram_buffer(8395) := X"1000FF23";
        ram_buffer(8396) := X"AE020050";
        ram_buffer(8397) := X"0C026495";
        ram_buffer(8398) := X"02002021";
        ram_buffer(8399) := X"1000FEF5";
        ram_buffer(8400) := X"AE020044";
        ram_buffer(8401) := X"8E020004";
        ram_buffer(8402) := X"00000000";
        ram_buffer(8403) := X"8C420000";
        ram_buffer(8404) := X"00002821";
        ram_buffer(8405) := X"0040F809";
        ram_buffer(8406) := X"02002021";
        ram_buffer(8407) := X"1000FEA1";
        ram_buffer(8408) := X"AE02003C";
        ram_buffer(8409) := X"0C026495";
        ram_buffer(8410) := X"02002021";
        ram_buffer(8411) := X"1000FEB0";
        ram_buffer(8412) := X"AE020040";
        ram_buffer(8413) := X"8C820010";
        ram_buffer(8414) := X"27BDFFE0";
        ram_buffer(8415) := X"24030064";
        ram_buffer(8416) := X"AFB10014";
        ram_buffer(8417) := X"AFB00010";
        ram_buffer(8418) := X"AFBF001C";
        ram_buffer(8419) := X"AFB20018";
        ram_buffer(8420) := X"8C900034";
        ram_buffer(8421) := X"1043000A";
        ram_buffer(8422) := X"00808821";
        ram_buffer(8423) := X"8C830000";
        ram_buffer(8424) := X"24050012";
        ram_buffer(8425) := X"AC620018";
        ram_buffer(8426) := X"8C820000";
        ram_buffer(8427) := X"AC650014";
        ram_buffer(8428) := X"8C420000";
        ram_buffer(8429) := X"00000000";
        ram_buffer(8430) := X"0040F809";
        ram_buffer(8431) := X"00000000";
        ram_buffer(8432) := X"24020003";
        ram_buffer(8433) := X"12020096";
        ram_buffer(8434) := X"2A020005";
        ram_buffer(8435) := X"1440006C";
        ram_buffer(8436) := X"001010C0";
        ram_buffer(8437) := X"8E240004";
        ram_buffer(8438) := X"00109040";
        ram_buffer(8439) := X"00529023";
        ram_buffer(8440) := X"00121940";
        ram_buffer(8441) := X"8C820000";
        ram_buffer(8442) := X"00123080";
        ram_buffer(8443) := X"00C33021";
        ram_buffer(8444) := X"02202021";
        ram_buffer(8445) := X"0040F809";
        ram_buffer(8446) := X"00002821";
        ram_buffer(8447) := X"AE2200A4";
        ram_buffer(8448) := X"AE3200A0";
        ram_buffer(8449) := X"00001821";
        ram_buffer(8450) := X"24040001";
        ram_buffer(8451) := X"AC430004";
        ram_buffer(8452) := X"24630001";
        ram_buffer(8453) := X"0070282A";
        ram_buffer(8454) := X"AC440000";
        ram_buffer(8455) := X"AC400014";
        ram_buffer(8456) := X"AC400018";
        ram_buffer(8457) := X"AC40001C";
        ram_buffer(8458) := X"AC440020";
        ram_buffer(8459) := X"14A0FFF7";
        ram_buffer(8460) := X"24420024";
        ram_buffer(8461) := X"1A000095";
        ram_buffer(8462) := X"24050001";
        ram_buffer(8463) := X"00401821";
        ram_buffer(8464) := X"00002021";
        ram_buffer(8465) := X"24070005";
        ram_buffer(8466) := X"24060002";
        ram_buffer(8467) := X"AC640004";
        ram_buffer(8468) := X"24840001";
        ram_buffer(8469) := X"AC650000";
        ram_buffer(8470) := X"AC650014";
        ram_buffer(8471) := X"AC670018";
        ram_buffer(8472) := X"AC60001C";
        ram_buffer(8473) := X"AC660020";
        ram_buffer(8474) := X"1604FFF8";
        ram_buffer(8475) := X"24630024";
        ram_buffer(8476) := X"00101940";
        ram_buffer(8477) := X"00104880";
        ram_buffer(8478) := X"01234821";
        ram_buffer(8479) := X"00491021";
        ram_buffer(8480) := X"00401821";
        ram_buffer(8481) := X"00002021";
        ram_buffer(8482) := X"24080001";
        ram_buffer(8483) := X"24070006";
        ram_buffer(8484) := X"2406003F";
        ram_buffer(8485) := X"24050002";
        ram_buffer(8486) := X"AC640004";
        ram_buffer(8487) := X"24840001";
        ram_buffer(8488) := X"AC680000";
        ram_buffer(8489) := X"AC670014";
        ram_buffer(8490) := X"AC660018";
        ram_buffer(8491) := X"AC60001C";
        ram_buffer(8492) := X"AC650020";
        ram_buffer(8493) := X"1604FFF8";
        ram_buffer(8494) := X"24630024";
        ram_buffer(8495) := X"00491021";
        ram_buffer(8496) := X"00001821";
        ram_buffer(8497) := X"24040001";
        ram_buffer(8498) := X"2407003F";
        ram_buffer(8499) := X"24060002";
        ram_buffer(8500) := X"AC430004";
        ram_buffer(8501) := X"24630001";
        ram_buffer(8502) := X"0070282A";
        ram_buffer(8503) := X"AC440000";
        ram_buffer(8504) := X"AC440014";
        ram_buffer(8505) := X"AC470018";
        ram_buffer(8506) := X"AC46001C";
        ram_buffer(8507) := X"AC440020";
        ram_buffer(8508) := X"24080002";
        ram_buffer(8509) := X"14A0FFF6";
        ram_buffer(8510) := X"24420024";
        ram_buffer(8511) := X"2A030005";
        ram_buffer(8512) := X"14600034";
        ram_buffer(8513) := X"00001821";
        ram_buffer(8514) := X"24040001";
        ram_buffer(8515) := X"AC430004";
        ram_buffer(8516) := X"24630001";
        ram_buffer(8517) := X"0070282A";
        ram_buffer(8518) := X"AC440000";
        ram_buffer(8519) := X"AC400014";
        ram_buffer(8520) := X"AC400018";
        ram_buffer(8521) := X"AC44001C";
        ram_buffer(8522) := X"AC400020";
        ram_buffer(8523) := X"14A0FFF7";
        ram_buffer(8524) := X"24420024";
        ram_buffer(8525) := X"1A00000C";
        ram_buffer(8526) := X"00001821";
        ram_buffer(8527) := X"24040001";
        ram_buffer(8528) := X"2405003F";
        ram_buffer(8529) := X"AC430004";
        ram_buffer(8530) := X"24630001";
        ram_buffer(8531) := X"AC440000";
        ram_buffer(8532) := X"AC440014";
        ram_buffer(8533) := X"AC450018";
        ram_buffer(8534) := X"AC44001C";
        ram_buffer(8535) := X"AC400020";
        ram_buffer(8536) := X"1603FFF8";
        ram_buffer(8537) := X"24420024";
        ram_buffer(8538) := X"8FBF001C";
        ram_buffer(8539) := X"8FB20018";
        ram_buffer(8540) := X"8FB10014";
        ram_buffer(8541) := X"8FB00010";
        ram_buffer(8542) := X"03E00008";
        ram_buffer(8543) := X"27BD0020";
        ram_buffer(8544) := X"8E220004";
        ram_buffer(8545) := X"00109080";
        ram_buffer(8546) := X"26520002";
        ram_buffer(8547) := X"00121940";
        ram_buffer(8548) := X"00123080";
        ram_buffer(8549) := X"8C420000";
        ram_buffer(8550) := X"00C33021";
        ram_buffer(8551) := X"00002821";
        ram_buffer(8552) := X"0040F809";
        ram_buffer(8553) := X"02202021";
        ram_buffer(8554) := X"AE2200A4";
        ram_buffer(8555) := X"AE3200A0";
        ram_buffer(8556) := X"1E00008F";
        ram_buffer(8557) := X"AC500000";
        ram_buffer(8558) := X"24030001";
        ram_buffer(8559) := X"AC400018";
        ram_buffer(8560) := X"AC400014";
        ram_buffer(8561) := X"AC40001C";
        ram_buffer(8562) := X"AC430020";
        ram_buffer(8563) := X"1000FF99";
        ram_buffer(8564) := X"24420024";
        ram_buffer(8565) := X"2A030002";
        ram_buffer(8566) := X"AC500000";
        ram_buffer(8567) := X"14600009";
        ram_buffer(8568) := X"AC400004";
        ram_buffer(8569) := X"24030001";
        ram_buffer(8570) := X"12080007";
        ram_buffer(8571) := X"AC430008";
        ram_buffer(8572) := X"24030004";
        ram_buffer(8573) := X"16030003";
        ram_buffer(8574) := X"AC48000C";
        ram_buffer(8575) := X"24030003";
        ram_buffer(8576) := X"AC430010";
        ram_buffer(8577) := X"24030001";
        ram_buffer(8578) := X"AC400018";
        ram_buffer(8579) := X"AC400014";
        ram_buffer(8580) := X"AC43001C";
        ram_buffer(8581) := X"AC400020";
        ram_buffer(8582) := X"1000FFC6";
        ram_buffer(8583) := X"24420024";
        ram_buffer(8584) := X"8E220038";
        ram_buffer(8585) := X"00000000";
        ram_buffer(8586) := X"1050001A";
        ram_buffer(8587) := X"02202021";
        ram_buffer(8588) := X"8E220004";
        ram_buffer(8589) := X"00000000";
        ram_buffer(8590) := X"8C420000";
        ram_buffer(8591) := X"240601F8";
        ram_buffer(8592) := X"0040F809";
        ram_buffer(8593) := X"00002821";
        ram_buffer(8594) := X"8E230038";
        ram_buffer(8595) := X"2404000E";
        ram_buffer(8596) := X"AE2200A4";
        ram_buffer(8597) := X"1070001F";
        ram_buffer(8598) := X"AE2400A0";
        ram_buffer(8599) := X"AC500000";
        ram_buffer(8600) := X"AC400004";
        ram_buffer(8601) := X"24040001";
        ram_buffer(8602) := X"2A030003";
        ram_buffer(8603) := X"1460FFD2";
        ram_buffer(8604) := X"AC440008";
        ram_buffer(8605) := X"24040002";
        ram_buffer(8606) := X"24030003";
        ram_buffer(8607) := X"1203FFCE";
        ram_buffer(8608) := X"AC44000C";
        ram_buffer(8609) := X"1000FFCC";
        ram_buffer(8610) := X"AC430010";
        ram_buffer(8611) := X"1000FFDD";
        ram_buffer(8612) := X"AC500000";
        ram_buffer(8613) := X"8E220004";
        ram_buffer(8614) := X"00000000";
        ram_buffer(8615) := X"8C420000";
        ram_buffer(8616) := X"24060168";
        ram_buffer(8617) := X"0040F809";
        ram_buffer(8618) := X"00002821";
        ram_buffer(8619) := X"8E230038";
        ram_buffer(8620) := X"2404000A";
        ram_buffer(8621) := X"AE2200A4";
        ram_buffer(8622) := X"10700006";
        ram_buffer(8623) := X"AE2400A0";
        ram_buffer(8624) := X"24030001";
        ram_buffer(8625) := X"AC500000";
        ram_buffer(8626) := X"AC400004";
        ram_buffer(8627) := X"1000FFE9";
        ram_buffer(8628) := X"AC430008";
        ram_buffer(8629) := X"24070005";
        ram_buffer(8630) := X"24030001";
        ram_buffer(8631) := X"24050002";
        ram_buffer(8632) := X"2404003F";
        ram_buffer(8633) := X"24060003";
        ram_buffer(8634) := X"AC47003C";
        ram_buffer(8635) := X"24070006";
        ram_buffer(8636) := X"AC460000";
        ram_buffer(8637) := X"AC400004";
        ram_buffer(8638) := X"AC430008";
        ram_buffer(8639) := X"AC45000C";
        ram_buffer(8640) := X"AC400018";
        ram_buffer(8641) := X"AC400014";
        ram_buffer(8642) := X"AC40001C";
        ram_buffer(8643) := X"AC430020";
        ram_buffer(8644) := X"AC430024";
        ram_buffer(8645) := X"AC400028";
        ram_buffer(8646) := X"AC430038";
        ram_buffer(8647) := X"AC400040";
        ram_buffer(8648) := X"AC450044";
        ram_buffer(8649) := X"AC430048";
        ram_buffer(8650) := X"AC45004C";
        ram_buffer(8651) := X"AC43005C";
        ram_buffer(8652) := X"AC440060";
        ram_buffer(8653) := X"AC400064";
        ram_buffer(8654) := X"AC430068";
        ram_buffer(8655) := X"AC43006C";
        ram_buffer(8656) := X"AC430070";
        ram_buffer(8657) := X"AC430080";
        ram_buffer(8658) := X"AC440084";
        ram_buffer(8659) := X"AC400088";
        ram_buffer(8660) := X"AC43008C";
        ram_buffer(8661) := X"AC430090";
        ram_buffer(8662) := X"AC400094";
        ram_buffer(8663) := X"AC4700A4";
        ram_buffer(8664) := X"AC4400A8";
        ram_buffer(8665) := X"AC4000AC";
        ram_buffer(8666) := X"AC4500B0";
        ram_buffer(8667) := X"AC4300B4";
        ram_buffer(8668) := X"AC4000B8";
        ram_buffer(8669) := X"AC4300C8";
        ram_buffer(8670) := X"AC4400CC";
        ram_buffer(8671) := X"AC4500D0";
        ram_buffer(8672) := X"AC4300D4";
        ram_buffer(8673) := X"AC4600D8";
        ram_buffer(8674) := X"AC4000DC";
        ram_buffer(8675) := X"AC4300E0";
        ram_buffer(8676) := X"AC4500E4";
        ram_buffer(8677) := X"AC4000F0";
        ram_buffer(8678) := X"AC4000EC";
        ram_buffer(8679) := X"AC4300F4";
        ram_buffer(8680) := X"AC4000F8";
        ram_buffer(8681) := X"AC4300FC";
        ram_buffer(8682) := X"AC450100";
        ram_buffer(8683) := X"AC430110";
        ram_buffer(8684) := X"AC440114";
        ram_buffer(8685) := X"AC430118";
        ram_buffer(8686) := X"AC40011C";
        ram_buffer(8687) := X"AC430120";
        ram_buffer(8688) := X"AC430124";
        ram_buffer(8689) := X"AC430134";
        ram_buffer(8690) := X"AC440138";
        ram_buffer(8691) := X"AC43013C";
        ram_buffer(8692) := X"AC400140";
        ram_buffer(8693) := X"AC430144";
        ram_buffer(8694) := X"AC400148";
        ram_buffer(8695) := X"AC430158";
        ram_buffer(8696) := X"AC44015C";
        ram_buffer(8697) := X"AC430160";
        ram_buffer(8698) := X"1000FF5F";
        ram_buffer(8699) := X"AC400164";
        ram_buffer(8700) := X"2A030002";
        ram_buffer(8701) := X"1460FF70";
        ram_buffer(8702) := X"AC400004";
        ram_buffer(8703) := X"1000FF9A";
        ram_buffer(8704) := X"24040001";
        ram_buffer(8705) := X"8C830004";
        ram_buffer(8706) := X"27BDFFE8";
        ram_buffer(8707) := X"8C620000";
        ram_buffer(8708) := X"24061000";
        ram_buffer(8709) := X"AFBF0014";
        ram_buffer(8710) := X"AFB00010";
        ram_buffer(8711) := X"8C900014";
        ram_buffer(8712) := X"0040F809";
        ram_buffer(8713) := X"24050001";
        ram_buffer(8714) := X"8FBF0014";
        ram_buffer(8715) := X"AE020018";
        ram_buffer(8716) := X"AE020000";
        ram_buffer(8717) := X"24021000";
        ram_buffer(8718) := X"AE020004";
        ram_buffer(8719) := X"8FB00010";
        ram_buffer(8720) := X"03E00008";
        ram_buffer(8721) := X"27BD0018";
        ram_buffer(8722) := X"27BDFFE0";
        ram_buffer(8723) := X"AFB00014";
        ram_buffer(8724) := X"8C900014";
        ram_buffer(8725) := X"AFB10018";
        ram_buffer(8726) := X"8E070014";
        ram_buffer(8727) := X"00808821";
        ram_buffer(8728) := X"8E040018";
        ram_buffer(8729) := X"24061000";
        ram_buffer(8730) := X"AFBF001C";
        ram_buffer(8731) := X"0C0278D7";
        ram_buffer(8732) := X"24050001";
        ram_buffer(8733) := X"24031000";
        ram_buffer(8734) := X"10430007";
        ram_buffer(8735) := X"00000000";
        ram_buffer(8736) := X"8E220000";
        ram_buffer(8737) := X"24040024";
        ram_buffer(8738) := X"8C430000";
        ram_buffer(8739) := X"AC440014";
        ram_buffer(8740) := X"0060F809";
        ram_buffer(8741) := X"02202021";
        ram_buffer(8742) := X"8E020018";
        ram_buffer(8743) := X"8FBF001C";
        ram_buffer(8744) := X"AE020000";
        ram_buffer(8745) := X"24021000";
        ram_buffer(8746) := X"AE020004";
        ram_buffer(8747) := X"8FB10018";
        ram_buffer(8748) := X"8FB00014";
        ram_buffer(8749) := X"24020001";
        ram_buffer(8750) := X"03E00008";
        ram_buffer(8751) := X"27BD0020";
        ram_buffer(8752) := X"27BDFFE0";
        ram_buffer(8753) := X"AFB00010";
        ram_buffer(8754) := X"8C900014";
        ram_buffer(8755) := X"AFB10014";
        ram_buffer(8756) := X"8E110004";
        ram_buffer(8757) := X"24021000";
        ram_buffer(8758) := X"00518823";
        ram_buffer(8759) := X"AFB20018";
        ram_buffer(8760) := X"AFBF001C";
        ram_buffer(8761) := X"1620001B";
        ram_buffer(8762) := X"00809021";
        ram_buffer(8763) := X"8E040014";
        ram_buffer(8764) := X"0C026F0C";
        ram_buffer(8765) := X"00000000";
        ram_buffer(8766) := X"8E020014";
        ram_buffer(8767) := X"00000000";
        ram_buffer(8768) := X"9442000C";
        ram_buffer(8769) := X"00000000";
        ram_buffer(8770) := X"30420040";
        ram_buffer(8771) := X"14400007";
        ram_buffer(8772) := X"24030024";
        ram_buffer(8773) := X"8FBF001C";
        ram_buffer(8774) := X"8FB20018";
        ram_buffer(8775) := X"8FB10014";
        ram_buffer(8776) := X"8FB00010";
        ram_buffer(8777) := X"03E00008";
        ram_buffer(8778) := X"27BD0020";
        ram_buffer(8779) := X"8E420000";
        ram_buffer(8780) := X"8FBF001C";
        ram_buffer(8781) := X"8FB10014";
        ram_buffer(8782) := X"8FB00010";
        ram_buffer(8783) := X"8C590000";
        ram_buffer(8784) := X"02402021";
        ram_buffer(8785) := X"8FB20018";
        ram_buffer(8786) := X"AC430014";
        ram_buffer(8787) := X"03200008";
        ram_buffer(8788) := X"27BD0020";
        ram_buffer(8789) := X"8E070014";
        ram_buffer(8790) := X"8E040018";
        ram_buffer(8791) := X"02203021";
        ram_buffer(8792) := X"0C0278D7";
        ram_buffer(8793) := X"24050001";
        ram_buffer(8794) := X"1222FFE0";
        ram_buffer(8795) := X"24040024";
        ram_buffer(8796) := X"8E420000";
        ram_buffer(8797) := X"00000000";
        ram_buffer(8798) := X"8C430000";
        ram_buffer(8799) := X"AC440014";
        ram_buffer(8800) := X"0060F809";
        ram_buffer(8801) := X"02402021";
        ram_buffer(8802) := X"1000FFD8";
        ram_buffer(8803) := X"00000000";
        ram_buffer(8804) := X"8C820014";
        ram_buffer(8805) := X"27BDFFE0";
        ram_buffer(8806) := X"AFB10018";
        ram_buffer(8807) := X"AFBF001C";
        ram_buffer(8808) := X"AFB00014";
        ram_buffer(8809) := X"10400010";
        ram_buffer(8810) := X"00A08821";
        ram_buffer(8811) := X"3C031009";
        ram_buffer(8812) := X"24638804";
        ram_buffer(8813) := X"AC430008";
        ram_buffer(8814) := X"3C031009";
        ram_buffer(8815) := X"24638848";
        ram_buffer(8816) := X"AC43000C";
        ram_buffer(8817) := X"8FBF001C";
        ram_buffer(8818) := X"3C031009";
        ram_buffer(8819) := X"246388C0";
        ram_buffer(8820) := X"AC510014";
        ram_buffer(8821) := X"8FB00014";
        ram_buffer(8822) := X"8FB10018";
        ram_buffer(8823) := X"AC430010";
        ram_buffer(8824) := X"03E00008";
        ram_buffer(8825) := X"27BD0020";
        ram_buffer(8826) := X"8C820004";
        ram_buffer(8827) := X"2406001C";
        ram_buffer(8828) := X"8C420000";
        ram_buffer(8829) := X"00002821";
        ram_buffer(8830) := X"0040F809";
        ram_buffer(8831) := X"00808021";
        ram_buffer(8832) := X"1000FFEA";
        ram_buffer(8833) := X"AE020014";
        ram_buffer(8834) := X"27BDFFE8";
        ram_buffer(8835) := X"00002821";
        ram_buffer(8836) := X"AFB00010";
        ram_buffer(8837) := X"AFBF0014";
        ram_buffer(8838) := X"0C02283F";
        ram_buffer(8839) := X"00808021";
        ram_buffer(8840) := X"8E0200A8";
        ram_buffer(8841) := X"00000000";
        ram_buffer(8842) := X"10400039";
        ram_buffer(8843) := X"00000000";
        ram_buffer(8844) := X"0C0260BE";
        ram_buffer(8845) := X"02002021";
        ram_buffer(8846) := X"8E0200AC";
        ram_buffer(8847) := X"00000000";
        ram_buffer(8848) := X"1440002B";
        ram_buffer(8849) := X"00000000";
        ram_buffer(8850) := X"8E0200DC";
        ram_buffer(8851) := X"00000000";
        ram_buffer(8852) := X"1440001D";
        ram_buffer(8853) := X"02002021";
        ram_buffer(8854) := X"0C024A2E";
        ram_buffer(8855) := X"00000000";
        ram_buffer(8856) := X"8E0200A0";
        ram_buffer(8857) := X"00000000";
        ram_buffer(8858) := X"28420002";
        ram_buffer(8859) := X"1440001D";
        ram_buffer(8860) := X"00000000";
        ram_buffer(8861) := X"24050001";
        ram_buffer(8862) := X"0C023E08";
        ram_buffer(8863) := X"02002021";
        ram_buffer(8864) := X"00002821";
        ram_buffer(8865) := X"0C023722";
        ram_buffer(8866) := X"02002021";
        ram_buffer(8867) := X"0C023694";
        ram_buffer(8868) := X"02002021";
        ram_buffer(8869) := X"8E020004";
        ram_buffer(8870) := X"00000000";
        ram_buffer(8871) := X"8C420018";
        ram_buffer(8872) := X"00000000";
        ram_buffer(8873) := X"0040F809";
        ram_buffer(8874) := X"02002021";
        ram_buffer(8875) := X"8E020154";
        ram_buffer(8876) := X"8FBF0014";
        ram_buffer(8877) := X"02002021";
        ram_buffer(8878) := X"8C590004";
        ram_buffer(8879) := X"8FB00010";
        ram_buffer(8880) := X"03200008";
        ram_buffer(8881) := X"27BD0018";
        ram_buffer(8882) := X"0C025C02";
        ram_buffer(8883) := X"00000000";
        ram_buffer(8884) := X"8E0200A0";
        ram_buffer(8885) := X"00000000";
        ram_buffer(8886) := X"28420002";
        ram_buffer(8887) := X"1040FFE5";
        ram_buffer(8888) := X"00000000";
        ram_buffer(8889) := X"8E0500B0";
        ram_buffer(8890) := X"1000FFE3";
        ram_buffer(8891) := X"0005282B";
        ram_buffer(8892) := X"8E020000";
        ram_buffer(8893) := X"24040001";
        ram_buffer(8894) := X"8C430000";
        ram_buffer(8895) := X"AC440014";
        ram_buffer(8896) := X"0060F809";
        ram_buffer(8897) := X"02002021";
        ram_buffer(8898) := X"1000FFD5";
        ram_buffer(8899) := X"00000000";
        ram_buffer(8900) := X"0C023F7A";
        ram_buffer(8901) := X"02002021";
        ram_buffer(8902) := X"0C02432E";
        ram_buffer(8903) := X"02002021";
        ram_buffer(8904) := X"00002821";
        ram_buffer(8905) := X"0C023916";
        ram_buffer(8906) := X"02002021";
        ram_buffer(8907) := X"1000FFC0";
        ram_buffer(8908) := X"00000000";
        ram_buffer(8909) := X"27BDF588";
        ram_buffer(8910) := X"AFB20A58";
        ram_buffer(8911) := X"8C9200A0";
        ram_buffer(8912) := X"AFBE0A70";
        ram_buffer(8913) := X"AFBF0A74";
        ram_buffer(8914) := X"AFB70A6C";
        ram_buffer(8915) := X"AFB60A68";
        ram_buffer(8916) := X"AFB50A64";
        ram_buffer(8917) := X"AFB40A60";
        ram_buffer(8918) := X"AFB30A5C";
        ram_buffer(8919) := X"AFB10A54";
        ram_buffer(8920) := X"AFB00A50";
        ram_buffer(8921) := X"1A4002C8";
        ram_buffer(8922) := X"0080F021";
        ram_buffer(8923) := X"8FD500A4";
        ram_buffer(8924) := X"00000000";
        ram_buffer(8925) := X"8EA20014";
        ram_buffer(8926) := X"00000000";
        ram_buffer(8927) := X"14400005";
        ram_buffer(8928) := X"2402003F";
        ram_buffer(8929) := X"8EA40018";
        ram_buffer(8930) := X"00000000";
        ram_buffer(8931) := X"10820261";
        ram_buffer(8932) := X"00000000";
        ram_buffer(8933) := X"8FD10034";
        ram_buffer(8934) := X"24020001";
        ram_buffer(8935) := X"1A2002CF";
        ram_buffer(8936) := X"AFC200DC";
        ram_buffer(8937) := X"00008021";
        ram_buffer(8938) := X"27A70010";
        ram_buffer(8939) := X"00E02021";
        ram_buffer(8940) := X"24060100";
        ram_buffer(8941) := X"0C02801D";
        ram_buffer(8942) := X"240500FF";
        ram_buffer(8943) := X"26100001";
        ram_buffer(8944) := X"1611FFFA";
        ram_buffer(8945) := X"24470100";
        ram_buffer(8946) := X"1A4001FE";
        ram_buffer(8947) := X"26B50004";
        ram_buffer(8948) := X"24120001";
        ram_buffer(8949) := X"8EB4FFFC";
        ram_buffer(8950) := X"00000000";
        ram_buffer(8951) := X"2682FFFF";
        ram_buffer(8952) := X"2C420004";
        ram_buffer(8953) := X"104000DD";
        ram_buffer(8954) := X"24030018";
        ram_buffer(8955) := X"02A09821";
        ram_buffer(8956) := X"00008821";
        ram_buffer(8957) := X"8E700000";
        ram_buffer(8958) := X"00000000";
        ram_buffer(8959) := X"06000006";
        ram_buffer(8960) := X"03C02021";
        ram_buffer(8961) := X"8FC20034";
        ram_buffer(8962) := X"00000000";
        ram_buffer(8963) := X"0202102A";
        ram_buffer(8964) := X"1440000A";
        ram_buffer(8965) := X"00000000";
        ram_buffer(8966) := X"8FC20000";
        ram_buffer(8967) := X"24030011";
        ram_buffer(8968) := X"AC520018";
        ram_buffer(8969) := X"8FC50000";
        ram_buffer(8970) := X"AC430014";
        ram_buffer(8971) := X"8CA20000";
        ram_buffer(8972) := X"00000000";
        ram_buffer(8973) := X"0040F809";
        ram_buffer(8974) := X"00000000";
        ram_buffer(8975) := X"1A200006";
        ram_buffer(8976) := X"00000000";
        ram_buffer(8977) := X"8E62FFFC";
        ram_buffer(8978) := X"00000000";
        ram_buffer(8979) := X"0050802A";
        ram_buffer(8980) := X"12000137";
        ram_buffer(8981) := X"24030011";
        ram_buffer(8982) := X"26310001";
        ram_buffer(8983) := X"1691FFE5";
        ram_buffer(8984) := X"26730004";
        ram_buffer(8985) := X"8EA30010";
        ram_buffer(8986) := X"8FC200DC";
        ram_buffer(8987) := X"AFA30A3C";
        ram_buffer(8988) := X"8EA30018";
        ram_buffer(8989) := X"8EB00014";
        ram_buffer(8990) := X"AFA30A44";
        ram_buffer(8991) := X"8EB1001C";
        ram_buffer(8992) := X"104000CE";
        ram_buffer(8993) := X"00000000";
        ram_buffer(8994) := X"8FA30A3C";
        ram_buffer(8995) := X"00000000";
        ram_buffer(8996) := X"2C620040";
        ram_buffer(8997) := X"1040000A";
        ram_buffer(8998) := X"0203102A";
        ram_buffer(8999) := X"14400008";
        ram_buffer(9000) := X"2A020040";
        ram_buffer(9001) := X"10400006";
        ram_buffer(9002) := X"00000000";
        ram_buffer(9003) := X"8FA20A44";
        ram_buffer(9004) := X"00000000";
        ram_buffer(9005) := X"2C42000E";
        ram_buffer(9006) := X"144001BA";
        ram_buffer(9007) := X"2E22000E";
        ram_buffer(9008) := X"8FC20000";
        ram_buffer(9009) := X"2405000F";
        ram_buffer(9010) := X"AC520018";
        ram_buffer(9011) := X"8FC40000";
        ram_buffer(9012) := X"AC450014";
        ram_buffer(9013) := X"8C820000";
        ram_buffer(9014) := X"00000000";
        ram_buffer(9015) := X"0040F809";
        ram_buffer(9016) := X"03C02021";
        ram_buffer(9017) := X"8FA20A3C";
        ram_buffer(9018) := X"00000000";
        ram_buffer(9019) := X"14400102";
        ram_buffer(9020) := X"00000000";
        ram_buffer(9021) := X"16000103";
        ram_buffer(9022) := X"00000000";
        ram_buffer(9023) := X"1A80003B";
        ram_buffer(9024) := X"00000000";
        ram_buffer(9025) := X"8FA20A44";
        ram_buffer(9026) := X"AFB50A38";
        ram_buffer(9027) := X"2442FFFF";
        ram_buffer(9028) := X"AFA20A4C";
        ram_buffer(9029) := X"AFA00A48";
        ram_buffer(9030) := X"2413000F";
        ram_buffer(9031) := X"8FA20A38";
        ram_buffer(9032) := X"27A30010";
        ram_buffer(9033) := X"8C420000";
        ram_buffer(9034) := X"00000000";
        ram_buffer(9035) := X"00021200";
        ram_buffer(9036) := X"00621021";
        ram_buffer(9037) := X"8FA30A3C";
        ram_buffer(9038) := X"00000000";
        ram_buffer(9039) := X"10600006";
        ram_buffer(9040) := X"0000B021";
        ram_buffer(9041) := X"8C440000";
        ram_buffer(9042) := X"00000000";
        ram_buffer(9043) := X"04800157";
        ram_buffer(9044) := X"03C02021";
        ram_buffer(9045) := X"0060B021";
        ram_buffer(9046) := X"0216202A";
        ram_buffer(9047) := X"1480001B";
        ram_buffer(9048) := X"00000000";
        ram_buffer(9049) := X"8FA30A4C";
        ram_buffer(9050) := X"00000000";
        ram_buffer(9051) := X"122300FB";
        ram_buffer(9052) := X"00000000";
        ram_buffer(9053) := X"8FA30A44";
        ram_buffer(9054) := X"00000000";
        ram_buffer(9055) := X"14600131";
        ram_buffer(9056) := X"00162080";
        ram_buffer(9057) := X"0044B821";
        ram_buffer(9058) := X"8EE60000";
        ram_buffer(9059) := X"26D60001";
        ram_buffer(9060) := X"04C0000A";
        ram_buffer(9061) := X"03C02021";
        ram_buffer(9062) := X"8FC60000";
        ram_buffer(9063) := X"00000000";
        ram_buffer(9064) := X"ACD20018";
        ram_buffer(9065) := X"8FC70000";
        ram_buffer(9066) := X"ACD30014";
        ram_buffer(9067) := X"8CE60000";
        ram_buffer(9068) := X"00000000";
        ram_buffer(9069) := X"00C0F809";
        ram_buffer(9070) := X"00000000";
        ram_buffer(9071) := X"0216202A";
        ram_buffer(9072) := X"AEF10000";
        ram_buffer(9073) := X"1080FFF0";
        ram_buffer(9074) := X"26F70004";
        ram_buffer(9075) := X"8FA20A48";
        ram_buffer(9076) := X"8FA30A38";
        ram_buffer(9077) := X"24420001";
        ram_buffer(9078) := X"AFA20A48";
        ram_buffer(9079) := X"24630004";
        ram_buffer(9080) := X"0054102A";
        ram_buffer(9081) := X"1440FFCD";
        ram_buffer(9082) := X"AFA30A38";
        ram_buffer(9083) := X"8FC200A0";
        ram_buffer(9084) := X"26520001";
        ram_buffer(9085) := X"0052102A";
        ram_buffer(9086) := X"1040FF76";
        ram_buffer(9087) := X"26B50024";
        ram_buffer(9088) := X"8FC200DC";
        ram_buffer(9089) := X"00000000";
        ram_buffer(9090) := X"1440016A";
        ram_buffer(9091) := X"00000000";
        ram_buffer(9092) := X"8FD00034";
        ram_buffer(9093) := X"00000000";
        ram_buffer(9094) := X"1A000044";
        ram_buffer(9095) := X"00000000";
        ram_buffer(9096) := X"8FA20A10";
        ram_buffer(9097) := X"00000000";
        ram_buffer(9098) := X"1040020E";
        ram_buffer(9099) := X"2404002C";
        ram_buffer(9100) := X"2A020002";
        ram_buffer(9101) := X"1440003D";
        ram_buffer(9102) := X"00000000";
        ram_buffer(9103) := X"8FA20A14";
        ram_buffer(9104) := X"00000000";
        ram_buffer(9105) := X"104001FE";
        ram_buffer(9106) := X"2404002C";
        ram_buffer(9107) := X"2A020003";
        ram_buffer(9108) := X"14400036";
        ram_buffer(9109) := X"00000000";
        ram_buffer(9110) := X"8FA20A18";
        ram_buffer(9111) := X"00000000";
        ram_buffer(9112) := X"104001EE";
        ram_buffer(9113) := X"2404002C";
        ram_buffer(9114) := X"2A020004";
        ram_buffer(9115) := X"1440002F";
        ram_buffer(9116) := X"00000000";
        ram_buffer(9117) := X"8FA20A1C";
        ram_buffer(9118) := X"00000000";
        ram_buffer(9119) := X"104001DE";
        ram_buffer(9120) := X"2404002C";
        ram_buffer(9121) := X"2A020005";
        ram_buffer(9122) := X"14400028";
        ram_buffer(9123) := X"00000000";
        ram_buffer(9124) := X"8FA20A20";
        ram_buffer(9125) := X"00000000";
        ram_buffer(9126) := X"104001CE";
        ram_buffer(9127) := X"2404002C";
        ram_buffer(9128) := X"2A020006";
        ram_buffer(9129) := X"14400021";
        ram_buffer(9130) := X"00000000";
        ram_buffer(9131) := X"8FA20A24";
        ram_buffer(9132) := X"00000000";
        ram_buffer(9133) := X"104001B5";
        ram_buffer(9134) := X"2404002C";
        ram_buffer(9135) := X"2A020007";
        ram_buffer(9136) := X"1440001A";
        ram_buffer(9137) := X"00000000";
        ram_buffer(9138) := X"8FA20A28";
        ram_buffer(9139) := X"00000000";
        ram_buffer(9140) := X"104001A5";
        ram_buffer(9141) := X"2404002C";
        ram_buffer(9142) := X"2A020008";
        ram_buffer(9143) := X"14400013";
        ram_buffer(9144) := X"00000000";
        ram_buffer(9145) := X"8FA20A2C";
        ram_buffer(9146) := X"00000000";
        ram_buffer(9147) := X"104001B0";
        ram_buffer(9148) := X"2404002C";
        ram_buffer(9149) := X"2A020009";
        ram_buffer(9150) := X"1440000C";
        ram_buffer(9151) := X"00000000";
        ram_buffer(9152) := X"8FA20A30";
        ram_buffer(9153) := X"00000000";
        ram_buffer(9154) := X"1040018E";
        ram_buffer(9155) := X"2404002C";
        ram_buffer(9156) := X"2A10000A";
        ram_buffer(9157) := X"16000005";
        ram_buffer(9158) := X"00000000";
        ram_buffer(9159) := X"8FA20A34";
        ram_buffer(9160) := X"00000000";
        ram_buffer(9161) := X"1040016A";
        ram_buffer(9162) := X"00000000";
        ram_buffer(9163) := X"8FBF0A74";
        ram_buffer(9164) := X"8FBE0A70";
        ram_buffer(9165) := X"8FB70A6C";
        ram_buffer(9166) := X"8FB60A68";
        ram_buffer(9167) := X"8FB50A64";
        ram_buffer(9168) := X"8FB40A60";
        ram_buffer(9169) := X"8FB30A5C";
        ram_buffer(9170) := X"8FB20A58";
        ram_buffer(9171) := X"8FB10A54";
        ram_buffer(9172) := X"8FB00A50";
        ram_buffer(9173) := X"03E00008";
        ram_buffer(9174) := X"27BD0A78";
        ram_buffer(9175) := X"8FC20000";
        ram_buffer(9176) := X"00000000";
        ram_buffer(9177) := X"AC540018";
        ram_buffer(9178) := X"8FC50000";
        ram_buffer(9179) := X"AC430014";
        ram_buffer(9180) := X"24020004";
        ram_buffer(9181) := X"ACA2001C";
        ram_buffer(9182) := X"8FC20000";
        ram_buffer(9183) := X"00000000";
        ram_buffer(9184) := X"8C420000";
        ram_buffer(9185) := X"00000000";
        ram_buffer(9186) := X"0040F809";
        ram_buffer(9187) := X"03C02021";
        ram_buffer(9188) := X"1E80FF17";
        ram_buffer(9189) := X"02A09821";
        ram_buffer(9190) := X"8EA30010";
        ram_buffer(9191) := X"8FC200DC";
        ram_buffer(9192) := X"AFA30A3C";
        ram_buffer(9193) := X"8EA30018";
        ram_buffer(9194) := X"8EB00014";
        ram_buffer(9195) := X"AFA30A44";
        ram_buffer(9196) := X"8EB1001C";
        ram_buffer(9197) := X"1440FF34";
        ram_buffer(9198) := X"00000000";
        ram_buffer(9199) := X"8FA20A3C";
        ram_buffer(9200) := X"00000000";
        ram_buffer(9201) := X"14400003";
        ram_buffer(9202) := X"2402003F";
        ram_buffer(9203) := X"120200EF";
        ram_buffer(9204) := X"00000000";
        ram_buffer(9205) := X"8FC20000";
        ram_buffer(9206) := X"2405000F";
        ram_buffer(9207) := X"AC520018";
        ram_buffer(9208) := X"8FC40000";
        ram_buffer(9209) := X"AC450014";
        ram_buffer(9210) := X"8C820000";
        ram_buffer(9211) := X"00000000";
        ram_buffer(9212) := X"0040F809";
        ram_buffer(9213) := X"03C02021";
        ram_buffer(9214) := X"1A80FF7C";
        ram_buffer(9215) := X"27A20010";
        ram_buffer(9216) := X"8EB00000";
        ram_buffer(9217) := X"00000000";
        ram_buffer(9218) := X"00108080";
        ram_buffer(9219) := X"00501021";
        ram_buffer(9220) := X"8C420A00";
        ram_buffer(9221) := X"00000000";
        ram_buffer(9222) := X"144000D1";
        ram_buffer(9223) := X"24030011";
        ram_buffer(9224) := X"27A20010";
        ram_buffer(9225) := X"00508021";
        ram_buffer(9226) := X"24020001";
        ram_buffer(9227) := X"1282FF6F";
        ram_buffer(9228) := X"AE020A00";
        ram_buffer(9229) := X"8EB00004";
        ram_buffer(9230) := X"27A20010";
        ram_buffer(9231) := X"00108080";
        ram_buffer(9232) := X"00501021";
        ram_buffer(9233) := X"8C420A00";
        ram_buffer(9234) := X"00000000";
        ram_buffer(9235) := X"144000B9";
        ram_buffer(9236) := X"24030011";
        ram_buffer(9237) := X"27A20010";
        ram_buffer(9238) := X"00508021";
        ram_buffer(9239) := X"24020001";
        ram_buffer(9240) := X"AE020A00";
        ram_buffer(9241) := X"24020002";
        ram_buffer(9242) := X"1282FF60";
        ram_buffer(9243) := X"27A20010";
        ram_buffer(9244) := X"8EB00008";
        ram_buffer(9245) := X"00000000";
        ram_buffer(9246) := X"00108080";
        ram_buffer(9247) := X"00501021";
        ram_buffer(9248) := X"8C420A00";
        ram_buffer(9249) := X"00000000";
        ram_buffer(9250) := X"1440009F";
        ram_buffer(9251) := X"24030011";
        ram_buffer(9252) := X"27A20010";
        ram_buffer(9253) := X"00508021";
        ram_buffer(9254) := X"24020001";
        ram_buffer(9255) := X"AE020A00";
        ram_buffer(9256) := X"24020003";
        ram_buffer(9257) := X"1282FF51";
        ram_buffer(9258) := X"27A20010";
        ram_buffer(9259) := X"8EB0000C";
        ram_buffer(9260) := X"00000000";
        ram_buffer(9261) := X"00108080";
        ram_buffer(9262) := X"00501021";
        ram_buffer(9263) := X"8C420A00";
        ram_buffer(9264) := X"00000000";
        ram_buffer(9265) := X"14400085";
        ram_buffer(9266) := X"24030011";
        ram_buffer(9267) := X"27A20010";
        ram_buffer(9268) := X"00508021";
        ram_buffer(9269) := X"24020001";
        ram_buffer(9270) := X"AE020A00";
        ram_buffer(9271) := X"8FC200A0";
        ram_buffer(9272) := X"26520001";
        ram_buffer(9273) := X"0052102A";
        ram_buffer(9274) := X"1040FEBA";
        ram_buffer(9275) := X"26B50024";
        ram_buffer(9276) := X"1000FF43";
        ram_buffer(9277) := X"00000000";
        ram_buffer(9278) := X"24020001";
        ram_buffer(9279) := X"1282FF01";
        ram_buffer(9280) := X"00000000";
        ram_buffer(9281) := X"8FC20000";
        ram_buffer(9282) := X"2405000F";
        ram_buffer(9283) := X"AC520018";
        ram_buffer(9284) := X"8FC40000";
        ram_buffer(9285) := X"AC450014";
        ram_buffer(9286) := X"8C820000";
        ram_buffer(9287) := X"00000000";
        ram_buffer(9288) := X"0040F809";
        ram_buffer(9289) := X"03C02021";
        ram_buffer(9290) := X"1000FEF4";
        ram_buffer(9291) := X"00000000";
        ram_buffer(9292) := X"8FC20000";
        ram_buffer(9293) := X"00000000";
        ram_buffer(9294) := X"AC520018";
        ram_buffer(9295) := X"8FC50000";
        ram_buffer(9296) := X"AC430014";
        ram_buffer(9297) := X"8CA20000";
        ram_buffer(9298) := X"00000000";
        ram_buffer(9299) := X"0040F809";
        ram_buffer(9300) := X"03C02021";
        ram_buffer(9301) := X"1000FEC1";
        ram_buffer(9302) := X"26310001";
        ram_buffer(9303) := X"8FA30A44";
        ram_buffer(9304) := X"00162080";
        ram_buffer(9305) := X"14600030";
        ram_buffer(9306) := X"0044B821";
        ram_buffer(9307) := X"8EE60000";
        ram_buffer(9308) := X"00000000";
        ram_buffer(9309) := X"04C0000C";
        ram_buffer(9310) := X"26D60001";
        ram_buffer(9311) := X"10C0000A";
        ram_buffer(9312) := X"03C02021";
        ram_buffer(9313) := X"8FC60000";
        ram_buffer(9314) := X"00000000";
        ram_buffer(9315) := X"ACD20018";
        ram_buffer(9316) := X"8FC70000";
        ram_buffer(9317) := X"ACD30014";
        ram_buffer(9318) := X"8CE60000";
        ram_buffer(9319) := X"00000000";
        ram_buffer(9320) := X"00C0F809";
        ram_buffer(9321) := X"00000000";
        ram_buffer(9322) := X"0216202A";
        ram_buffer(9323) := X"AEF10000";
        ram_buffer(9324) := X"1080FFEE";
        ram_buffer(9325) := X"26F70004";
        ram_buffer(9326) := X"8FA20A48";
        ram_buffer(9327) := X"8FA30A38";
        ram_buffer(9328) := X"24420001";
        ram_buffer(9329) := X"AFA20A48";
        ram_buffer(9330) := X"24630004";
        ram_buffer(9331) := X"0054102A";
        ram_buffer(9332) := X"1440FED2";
        ram_buffer(9333) := X"AFA30A38";
        ram_buffer(9334) := X"1000FF04";
        ram_buffer(9335) := X"00000000";
        ram_buffer(9336) := X"8FA20A44";
        ram_buffer(9337) := X"00000000";
        ram_buffer(9338) := X"1046000A";
        ram_buffer(9339) := X"03C02021";
        ram_buffer(9340) := X"8FC60000";
        ram_buffer(9341) := X"00000000";
        ram_buffer(9342) := X"ACD20018";
        ram_buffer(9343) := X"8FC70000";
        ram_buffer(9344) := X"ACD30014";
        ram_buffer(9345) := X"8CE60000";
        ram_buffer(9346) := X"00000000";
        ram_buffer(9347) := X"00C0F809";
        ram_buffer(9348) := X"00000000";
        ram_buffer(9349) := X"26D60001";
        ram_buffer(9350) := X"0216202A";
        ram_buffer(9351) := X"AEF10000";
        ram_buffer(9352) := X"1480FEEA";
        ram_buffer(9353) := X"26F70004";
        ram_buffer(9354) := X"8EE60000";
        ram_buffer(9355) := X"00000000";
        ram_buffer(9356) := X"04C1FFEB";
        ram_buffer(9357) := X"00000000";
        ram_buffer(9358) := X"8FC60000";
        ram_buffer(9359) := X"1000FFEE";
        ram_buffer(9360) := X"03C02021";
        ram_buffer(9361) := X"00441021";
        ram_buffer(9362) := X"8FC60000";
        ram_buffer(9363) := X"AFA20A40";
        ram_buffer(9364) := X"ACD20018";
        ram_buffer(9365) := X"8FC70000";
        ram_buffer(9366) := X"ACD30014";
        ram_buffer(9367) := X"8CE60000";
        ram_buffer(9368) := X"00000000";
        ram_buffer(9369) := X"00C0F809";
        ram_buffer(9370) := X"03C02021";
        ram_buffer(9371) := X"26D60001";
        ram_buffer(9372) := X"8FA20A40";
        ram_buffer(9373) := X"0216202A";
        ram_buffer(9374) := X"AC510000";
        ram_buffer(9375) := X"1080FFF2";
        ram_buffer(9376) := X"24420004";
        ram_buffer(9377) := X"8FA20A48";
        ram_buffer(9378) := X"8FA30A38";
        ram_buffer(9379) := X"24420001";
        ram_buffer(9380) := X"AFA20A48";
        ram_buffer(9381) := X"24630004";
        ram_buffer(9382) := X"0054102A";
        ram_buffer(9383) := X"1440FE9F";
        ram_buffer(9384) := X"AFA30A38";
        ram_buffer(9385) := X"1000FED1";
        ram_buffer(9386) := X"00000000";
        ram_buffer(9387) := X"8FC50000";
        ram_buffer(9388) := X"00000000";
        ram_buffer(9389) := X"ACB20018";
        ram_buffer(9390) := X"8FC60000";
        ram_buffer(9391) := X"ACB30014";
        ram_buffer(9392) := X"8CC60000";
        ram_buffer(9393) := X"AFA20A40";
        ram_buffer(9394) := X"00C0F809";
        ram_buffer(9395) := X"0060B021";
        ram_buffer(9396) := X"8FA20A40";
        ram_buffer(9397) := X"1000FEA1";
        ram_buffer(9398) := X"0216202A";
        ram_buffer(9399) := X"8FC20000";
        ram_buffer(9400) := X"00000000";
        ram_buffer(9401) := X"AC520018";
        ram_buffer(9402) := X"8FC50000";
        ram_buffer(9403) := X"AC430014";
        ram_buffer(9404) := X"8CA20000";
        ram_buffer(9405) := X"00000000";
        ram_buffer(9406) := X"0040F809";
        ram_buffer(9407) := X"03C02021";
        ram_buffer(9408) := X"1000FF73";
        ram_buffer(9409) := X"27A20010";
        ram_buffer(9410) := X"8FC20000";
        ram_buffer(9411) := X"00000000";
        ram_buffer(9412) := X"AC520018";
        ram_buffer(9413) := X"8FC50000";
        ram_buffer(9414) := X"AC430014";
        ram_buffer(9415) := X"8CA20000";
        ram_buffer(9416) := X"00000000";
        ram_buffer(9417) := X"0040F809";
        ram_buffer(9418) := X"03C02021";
        ram_buffer(9419) := X"1000FF59";
        ram_buffer(9420) := X"27A20010";
        ram_buffer(9421) := X"8FC20000";
        ram_buffer(9422) := X"00000000";
        ram_buffer(9423) := X"AC520018";
        ram_buffer(9424) := X"8FC50000";
        ram_buffer(9425) := X"AC430014";
        ram_buffer(9426) := X"8CA20000";
        ram_buffer(9427) := X"00000000";
        ram_buffer(9428) := X"0040F809";
        ram_buffer(9429) := X"03C02021";
        ram_buffer(9430) := X"1000FF3F";
        ram_buffer(9431) := X"27A20010";
        ram_buffer(9432) := X"8FC20000";
        ram_buffer(9433) := X"00000000";
        ram_buffer(9434) := X"AC520018";
        ram_buffer(9435) := X"8FC50000";
        ram_buffer(9436) := X"AC430014";
        ram_buffer(9437) := X"8CA20000";
        ram_buffer(9438) := X"00000000";
        ram_buffer(9439) := X"0040F809";
        ram_buffer(9440) := X"03C02021";
        ram_buffer(9441) := X"1000FF27";
        ram_buffer(9442) := X"27A20010";
        ram_buffer(9443) := X"1460FF11";
        ram_buffer(9444) := X"00000000";
        ram_buffer(9445) := X"1220FF18";
        ram_buffer(9446) := X"00000000";
        ram_buffer(9447) := X"1000FF0D";
        ram_buffer(9448) := X"00000000";
        ram_buffer(9449) := X"1440FE4F";
        ram_buffer(9450) := X"00000000";
        ram_buffer(9451) := X"1000FE44";
        ram_buffer(9452) := X"00000000";
        ram_buffer(9453) := X"8FD10034";
        ram_buffer(9454) := X"00000000";
        ram_buffer(9455) := X"1A20FEDB";
        ram_buffer(9456) := X"00000000";
        ram_buffer(9457) := X"8FA20010";
        ram_buffer(9458) := X"00000000";
        ram_buffer(9459) := X"04400106";
        ram_buffer(9460) := X"2404002C";
        ram_buffer(9461) := X"2A220002";
        ram_buffer(9462) := X"1440FED4";
        ram_buffer(9463) := X"00000000";
        ram_buffer(9464) := X"8FA20110";
        ram_buffer(9465) := X"00000000";
        ram_buffer(9466) := X"044000F6";
        ram_buffer(9467) := X"2404002C";
        ram_buffer(9468) := X"2A220003";
        ram_buffer(9469) := X"1440FECD";
        ram_buffer(9470) := X"00000000";
        ram_buffer(9471) := X"8FA20210";
        ram_buffer(9472) := X"00000000";
        ram_buffer(9473) := X"044000E6";
        ram_buffer(9474) := X"2404002C";
        ram_buffer(9475) := X"2A220004";
        ram_buffer(9476) := X"1440FEC6";
        ram_buffer(9477) := X"00000000";
        ram_buffer(9478) := X"8FA20310";
        ram_buffer(9479) := X"00000000";
        ram_buffer(9480) := X"044000D6";
        ram_buffer(9481) := X"2404002C";
        ram_buffer(9482) := X"2A220005";
        ram_buffer(9483) := X"1440FEBF";
        ram_buffer(9484) := X"00000000";
        ram_buffer(9485) := X"8FA20410";
        ram_buffer(9486) := X"00000000";
        ram_buffer(9487) := X"044000C6";
        ram_buffer(9488) := X"2404002C";
        ram_buffer(9489) := X"2A220006";
        ram_buffer(9490) := X"1440FEB8";
        ram_buffer(9491) := X"00000000";
        ram_buffer(9492) := X"8FA20510";
        ram_buffer(9493) := X"00000000";
        ram_buffer(9494) := X"044000B6";
        ram_buffer(9495) := X"2404002C";
        ram_buffer(9496) := X"2A220007";
        ram_buffer(9497) := X"1440FEB1";
        ram_buffer(9498) := X"00000000";
        ram_buffer(9499) := X"8FA20610";
        ram_buffer(9500) := X"00000000";
        ram_buffer(9501) := X"044000A6";
        ram_buffer(9502) := X"2404002C";
        ram_buffer(9503) := X"2A220008";
        ram_buffer(9504) := X"1440FEAA";
        ram_buffer(9505) := X"00000000";
        ram_buffer(9506) := X"8FA20710";
        ram_buffer(9507) := X"00000000";
        ram_buffer(9508) := X"04400096";
        ram_buffer(9509) := X"2404002C";
        ram_buffer(9510) := X"2A220009";
        ram_buffer(9511) := X"1440FEA3";
        ram_buffer(9512) := X"00000000";
        ram_buffer(9513) := X"8FA20810";
        ram_buffer(9514) := X"00000000";
        ram_buffer(9515) := X"04400082";
        ram_buffer(9516) := X"2404002C";
        ram_buffer(9517) := X"2A31000A";
        ram_buffer(9518) := X"1620FE9C";
        ram_buffer(9519) := X"00000000";
        ram_buffer(9520) := X"8FA20910";
        ram_buffer(9521) := X"00000000";
        ram_buffer(9522) := X"0441FE98";
        ram_buffer(9523) := X"00000000";
        ram_buffer(9524) := X"8FC20000";
        ram_buffer(9525) := X"2404002C";
        ram_buffer(9526) := X"AC440014";
        ram_buffer(9527) := X"8FBF0A74";
        ram_buffer(9528) := X"8FB70A6C";
        ram_buffer(9529) := X"8FB60A68";
        ram_buffer(9530) := X"8FB50A64";
        ram_buffer(9531) := X"8FB40A60";
        ram_buffer(9532) := X"8FB30A5C";
        ram_buffer(9533) := X"8FB20A58";
        ram_buffer(9534) := X"8FB10A54";
        ram_buffer(9535) := X"8FB00A50";
        ram_buffer(9536) := X"8C590000";
        ram_buffer(9537) := X"03C02021";
        ram_buffer(9538) := X"8FBE0A70";
        ram_buffer(9539) := X"03200008";
        ram_buffer(9540) := X"27BD0A78";
        ram_buffer(9541) := X"8FD00034";
        ram_buffer(9542) := X"00000000";
        ram_buffer(9543) := X"1A0000BB";
        ram_buffer(9544) := X"AFC000DC";
        ram_buffer(9545) := X"00103080";
        ram_buffer(9546) := X"00002821";
        ram_buffer(9547) := X"0C02801D";
        ram_buffer(9548) := X"27A40A10";
        ram_buffer(9549) := X"1E40FDA6";
        ram_buffer(9550) := X"26B50004";
        ram_buffer(9551) := X"1000FE38";
        ram_buffer(9552) := X"26B5FFFC";
        ram_buffer(9553) := X"8FC20000";
        ram_buffer(9554) := X"00000000";
        ram_buffer(9555) := X"8C450000";
        ram_buffer(9556) := X"AC440014";
        ram_buffer(9557) := X"00A0F809";
        ram_buffer(9558) := X"03C02021";
        ram_buffer(9559) := X"8FD00034";
        ram_buffer(9560) := X"1000FE6C";
        ram_buffer(9561) := X"2A10000A";
        ram_buffer(9562) := X"8FC20000";
        ram_buffer(9563) := X"00000000";
        ram_buffer(9564) := X"8C450000";
        ram_buffer(9565) := X"AC440014";
        ram_buffer(9566) := X"00A0F809";
        ram_buffer(9567) := X"03C02021";
        ram_buffer(9568) := X"8FD00034";
        ram_buffer(9569) := X"1000FE55";
        ram_buffer(9570) := X"2A020008";
        ram_buffer(9571) := X"8FC20000";
        ram_buffer(9572) := X"00000000";
        ram_buffer(9573) := X"8C450000";
        ram_buffer(9574) := X"AC440014";
        ram_buffer(9575) := X"00A0F809";
        ram_buffer(9576) := X"03C02021";
        ram_buffer(9577) := X"8FD00034";
        ram_buffer(9578) := X"1000FE45";
        ram_buffer(9579) := X"2A020007";
        ram_buffer(9580) := X"8FC20000";
        ram_buffer(9581) := X"00000000";
        ram_buffer(9582) := X"8C450000";
        ram_buffer(9583) := X"AC440014";
        ram_buffer(9584) := X"00A0F809";
        ram_buffer(9585) := X"03C02021";
        ram_buffer(9586) := X"8FD00034";
        ram_buffer(9587) := X"1000FE4A";
        ram_buffer(9588) := X"2A020009";
        ram_buffer(9589) := X"8FC20000";
        ram_buffer(9590) := X"00000000";
        ram_buffer(9591) := X"8C450000";
        ram_buffer(9592) := X"AC440014";
        ram_buffer(9593) := X"00A0F809";
        ram_buffer(9594) := X"03C02021";
        ram_buffer(9595) := X"8FD00034";
        ram_buffer(9596) := X"1000FE2C";
        ram_buffer(9597) := X"2A020006";
        ram_buffer(9598) := X"8FC20000";
        ram_buffer(9599) := X"00000000";
        ram_buffer(9600) := X"8C450000";
        ram_buffer(9601) := X"AC440014";
        ram_buffer(9602) := X"00A0F809";
        ram_buffer(9603) := X"03C02021";
        ram_buffer(9604) := X"8FD00034";
        ram_buffer(9605) := X"1000FE1C";
        ram_buffer(9606) := X"2A020005";
        ram_buffer(9607) := X"8FC20000";
        ram_buffer(9608) := X"00000000";
        ram_buffer(9609) := X"8C450000";
        ram_buffer(9610) := X"AC440014";
        ram_buffer(9611) := X"00A0F809";
        ram_buffer(9612) := X"03C02021";
        ram_buffer(9613) := X"8FD00034";
        ram_buffer(9614) := X"1000FE0C";
        ram_buffer(9615) := X"2A020004";
        ram_buffer(9616) := X"8FC20000";
        ram_buffer(9617) := X"00000000";
        ram_buffer(9618) := X"8C450000";
        ram_buffer(9619) := X"AC440014";
        ram_buffer(9620) := X"00A0F809";
        ram_buffer(9621) := X"03C02021";
        ram_buffer(9622) := X"8FD00034";
        ram_buffer(9623) := X"1000FDFC";
        ram_buffer(9624) := X"2A020003";
        ram_buffer(9625) := X"8FC20000";
        ram_buffer(9626) := X"00000000";
        ram_buffer(9627) := X"8C450000";
        ram_buffer(9628) := X"AC440014";
        ram_buffer(9629) := X"00A0F809";
        ram_buffer(9630) := X"03C02021";
        ram_buffer(9631) := X"8FD00034";
        ram_buffer(9632) := X"1000FDEC";
        ram_buffer(9633) := X"2A020002";
        ram_buffer(9634) := X"8C820000";
        ram_buffer(9635) := X"24060011";
        ram_buffer(9636) := X"AC400018";
        ram_buffer(9637) := X"8C850000";
        ram_buffer(9638) := X"AC460014";
        ram_buffer(9639) := X"8CA20000";
        ram_buffer(9640) := X"00000000";
        ram_buffer(9641) := X"0040F809";
        ram_buffer(9642) := X"00000000";
        ram_buffer(9643) := X"8FD200A0";
        ram_buffer(9644) := X"1000FD2E";
        ram_buffer(9645) := X"00000000";
        ram_buffer(9646) := X"8FC20000";
        ram_buffer(9647) := X"00000000";
        ram_buffer(9648) := X"8C450000";
        ram_buffer(9649) := X"AC440014";
        ram_buffer(9650) := X"00A0F809";
        ram_buffer(9651) := X"03C02021";
        ram_buffer(9652) := X"8FD10034";
        ram_buffer(9653) := X"1000FF78";
        ram_buffer(9654) := X"2A31000A";
        ram_buffer(9655) := X"1A40FE13";
        ram_buffer(9656) := X"26B50004";
        ram_buffer(9657) := X"1000FD3B";
        ram_buffer(9658) := X"24120001";
        ram_buffer(9659) := X"8FC20000";
        ram_buffer(9660) := X"00000000";
        ram_buffer(9661) := X"8C450000";
        ram_buffer(9662) := X"AC440014";
        ram_buffer(9663) := X"00A0F809";
        ram_buffer(9664) := X"03C02021";
        ram_buffer(9665) := X"8FD10034";
        ram_buffer(9666) := X"1000FF64";
        ram_buffer(9667) := X"2A220009";
        ram_buffer(9668) := X"8FC20000";
        ram_buffer(9669) := X"00000000";
        ram_buffer(9670) := X"8C450000";
        ram_buffer(9671) := X"AC440014";
        ram_buffer(9672) := X"00A0F809";
        ram_buffer(9673) := X"03C02021";
        ram_buffer(9674) := X"8FD10034";
        ram_buffer(9675) := X"1000FF54";
        ram_buffer(9676) := X"2A220008";
        ram_buffer(9677) := X"8FC20000";
        ram_buffer(9678) := X"00000000";
        ram_buffer(9679) := X"8C450000";
        ram_buffer(9680) := X"AC440014";
        ram_buffer(9681) := X"00A0F809";
        ram_buffer(9682) := X"03C02021";
        ram_buffer(9683) := X"8FD10034";
        ram_buffer(9684) := X"1000FF44";
        ram_buffer(9685) := X"2A220007";
        ram_buffer(9686) := X"8FC20000";
        ram_buffer(9687) := X"00000000";
        ram_buffer(9688) := X"8C450000";
        ram_buffer(9689) := X"AC440014";
        ram_buffer(9690) := X"00A0F809";
        ram_buffer(9691) := X"03C02021";
        ram_buffer(9692) := X"8FD10034";
        ram_buffer(9693) := X"1000FF34";
        ram_buffer(9694) := X"2A220006";
        ram_buffer(9695) := X"8FC20000";
        ram_buffer(9696) := X"00000000";
        ram_buffer(9697) := X"8C450000";
        ram_buffer(9698) := X"AC440014";
        ram_buffer(9699) := X"00A0F809";
        ram_buffer(9700) := X"03C02021";
        ram_buffer(9701) := X"8FD10034";
        ram_buffer(9702) := X"1000FF24";
        ram_buffer(9703) := X"2A220005";
        ram_buffer(9704) := X"8FC20000";
        ram_buffer(9705) := X"00000000";
        ram_buffer(9706) := X"8C450000";
        ram_buffer(9707) := X"AC440014";
        ram_buffer(9708) := X"00A0F809";
        ram_buffer(9709) := X"03C02021";
        ram_buffer(9710) := X"8FD10034";
        ram_buffer(9711) := X"1000FF14";
        ram_buffer(9712) := X"2A220004";
        ram_buffer(9713) := X"8FC20000";
        ram_buffer(9714) := X"00000000";
        ram_buffer(9715) := X"8C450000";
        ram_buffer(9716) := X"AC440014";
        ram_buffer(9717) := X"00A0F809";
        ram_buffer(9718) := X"03C02021";
        ram_buffer(9719) := X"8FD10034";
        ram_buffer(9720) := X"1000FF04";
        ram_buffer(9721) := X"2A220003";
        ram_buffer(9722) := X"8FC20000";
        ram_buffer(9723) := X"00000000";
        ram_buffer(9724) := X"8C450000";
        ram_buffer(9725) := X"AC440014";
        ram_buffer(9726) := X"00A0F809";
        ram_buffer(9727) := X"03C02021";
        ram_buffer(9728) := X"8FD10034";
        ram_buffer(9729) := X"1000FEF4";
        ram_buffer(9730) := X"2A220002";
        ram_buffer(9731) := X"1E40FCF0";
        ram_buffer(9732) := X"26B50004";
        ram_buffer(9733) := X"1000FDC5";
        ram_buffer(9734) := X"00000000";
        ram_buffer(9735) := X"8C820154";
        ram_buffer(9736) := X"8C830144";
        ram_buffer(9737) := X"27BDFFE8";
        ram_buffer(9738) := X"8C420008";
        ram_buffer(9739) := X"AFBF0014";
        ram_buffer(9740) := X"AFB00010";
        ram_buffer(9741) := X"00808021";
        ram_buffer(9742) := X"0040F809";
        ram_buffer(9743) := X"AC60000C";
        ram_buffer(9744) := X"8E020154";
        ram_buffer(9745) := X"8FBF0014";
        ram_buffer(9746) := X"02002021";
        ram_buffer(9747) := X"8C59000C";
        ram_buffer(9748) := X"8FB00010";
        ram_buffer(9749) := X"03200008";
        ram_buffer(9750) := X"27BD0018";
        ram_buffer(9751) := X"8C820164";
        ram_buffer(9752) := X"27BDFFE0";
        ram_buffer(9753) := X"8C420008";
        ram_buffer(9754) := X"AFB00014";
        ram_buffer(9755) := X"8C900144";
        ram_buffer(9756) := X"AFB10018";
        ram_buffer(9757) := X"AFBF001C";
        ram_buffer(9758) := X"0040F809";
        ram_buffer(9759) := X"00808821";
        ram_buffer(9760) := X"8E020014";
        ram_buffer(9761) := X"24030001";
        ram_buffer(9762) := X"1043001F";
        ram_buffer(9763) := X"00000000";
        ram_buffer(9764) := X"10400014";
        ram_buffer(9765) := X"24040002";
        ram_buffer(9766) := X"1444000A";
        ram_buffer(9767) := X"00000000";
        ram_buffer(9768) := X"8E2200B0";
        ram_buffer(9769) := X"00000000";
        ram_buffer(9770) := X"10400002";
        ram_buffer(9771) := X"00000000";
        ram_buffer(9772) := X"AE030014";
        ram_buffer(9773) := X"8E020020";
        ram_buffer(9774) := X"00000000";
        ram_buffer(9775) := X"24420001";
        ram_buffer(9776) := X"AE020020";
        ram_buffer(9777) := X"8E020018";
        ram_buffer(9778) := X"8FBF001C";
        ram_buffer(9779) := X"24420001";
        ram_buffer(9780) := X"AE020018";
        ram_buffer(9781) := X"8FB10018";
        ram_buffer(9782) := X"8FB00014";
        ram_buffer(9783) := X"03E00008";
        ram_buffer(9784) := X"27BD0020";
        ram_buffer(9785) := X"8E2200B0";
        ram_buffer(9786) := X"24030002";
        ram_buffer(9787) := X"1440FFF5";
        ram_buffer(9788) := X"AE030014";
        ram_buffer(9789) := X"8E020020";
        ram_buffer(9790) := X"00000000";
        ram_buffer(9791) := X"24420001";
        ram_buffer(9792) := X"1000FFF0";
        ram_buffer(9793) := X"AE020020";
        ram_buffer(9794) := X"24020002";
        ram_buffer(9795) := X"AE020014";
        ram_buffer(9796) := X"8E020018";
        ram_buffer(9797) := X"8FBF001C";
        ram_buffer(9798) := X"24420001";
        ram_buffer(9799) := X"AE020018";
        ram_buffer(9800) := X"8FB10018";
        ram_buffer(9801) := X"8FB00014";
        ram_buffer(9802) := X"03E00008";
        ram_buffer(9803) := X"27BD0020";
        ram_buffer(9804) := X"8C8200EC";
        ram_buffer(9805) := X"27BDFFD8";
        ram_buffer(9806) := X"24030001";
        ram_buffer(9807) := X"AFB00010";
        ram_buffer(9808) := X"AFBF0024";
        ram_buffer(9809) := X"AFB40020";
        ram_buffer(9810) := X"AFB3001C";
        ram_buffer(9811) := X"AFB20018";
        ram_buffer(9812) := X"AFB10014";
        ram_buffer(9813) := X"1043007F";
        ram_buffer(9814) := X"00808021";
        ram_buffer(9815) := X"2443FFFF";
        ram_buffer(9816) := X"2C630004";
        ram_buffer(9817) := X"106000B2";
        ram_buffer(9818) := X"00000000";
        ram_buffer(9819) := X"8E0500E0";
        ram_buffer(9820) := X"8E040018";
        ram_buffer(9821) := X"0C0264AB";
        ram_buffer(9822) := X"000528C0";
        ram_buffer(9823) := X"8E0500E4";
        ram_buffer(9824) := X"8E04001C";
        ram_buffer(9825) := X"AE020100";
        ram_buffer(9826) := X"0C0264AB";
        ram_buffer(9827) := X"000528C0";
        ram_buffer(9828) := X"8E0600EC";
        ram_buffer(9829) := X"AE020104";
        ram_buffer(9830) := X"18C00085";
        ram_buffer(9831) := X"AE000108";
        ram_buffer(9832) := X"261400F0";
        ram_buffer(9833) := X"00002821";
        ram_buffer(9834) := X"00009821";
        ram_buffer(9835) := X"2412000B";
        ram_buffer(9836) := X"8E820000";
        ram_buffer(9837) := X"00000000";
        ram_buffer(9838) := X"8C430008";
        ram_buffer(9839) := X"8C47001C";
        ram_buffer(9840) := X"8C44000C";
        ram_buffer(9841) := X"14600002";
        ram_buffer(9842) := X"00E3001B";
        ram_buffer(9843) := X"0007000D";
        ram_buffer(9844) := X"000340C0";
        ram_buffer(9845) := X"AC430034";
        ram_buffer(9846) := X"AC440038";
        ram_buffer(9847) := X"AC480040";
        ram_buffer(9848) := X"00003810";
        ram_buffer(9849) := X"00000000";
        ram_buffer(9850) := X"00000000";
        ram_buffer(9851) := X"00640018";
        ram_buffer(9852) := X"00008812";
        ram_buffer(9853) := X"10E00002";
        ram_buffer(9854) := X"AC51003C";
        ram_buffer(9855) := X"00E01821";
        ram_buffer(9856) := X"8C470020";
        ram_buffer(9857) := X"00000000";
        ram_buffer(9858) := X"14800002";
        ram_buffer(9859) := X"00E4001B";
        ram_buffer(9860) := X"0007000D";
        ram_buffer(9861) := X"00003810";
        ram_buffer(9862) := X"10E00002";
        ram_buffer(9863) := X"AC430044";
        ram_buffer(9864) := X"00E02021";
        ram_buffer(9865) := X"02252821";
        ram_buffer(9866) := X"28A5000B";
        ram_buffer(9867) := X"10A00075";
        ram_buffer(9868) := X"AC440048";
        ram_buffer(9869) := X"1A200040";
        ram_buffer(9870) := X"2624FFFF";
        ram_buffer(9871) := X"8E020108";
        ram_buffer(9872) := X"00000000";
        ram_buffer(9873) := X"24430042";
        ram_buffer(9874) := X"00031880";
        ram_buffer(9875) := X"02031821";
        ram_buffer(9876) := X"24450001";
        ram_buffer(9877) := X"18800036";
        ram_buffer(9878) := X"AC730004";
        ram_buffer(9879) := X"24430043";
        ram_buffer(9880) := X"00031880";
        ram_buffer(9881) := X"02031821";
        ram_buffer(9882) := X"2A270003";
        ram_buffer(9883) := X"14E00030";
        ram_buffer(9884) := X"AC730004";
        ram_buffer(9885) := X"24430044";
        ram_buffer(9886) := X"00031880";
        ram_buffer(9887) := X"02031821";
        ram_buffer(9888) := X"2A270004";
        ram_buffer(9889) := X"14E0002A";
        ram_buffer(9890) := X"AC730004";
        ram_buffer(9891) := X"24430045";
        ram_buffer(9892) := X"00031880";
        ram_buffer(9893) := X"02031821";
        ram_buffer(9894) := X"2A270005";
        ram_buffer(9895) := X"14E00024";
        ram_buffer(9896) := X"AC730004";
        ram_buffer(9897) := X"24430046";
        ram_buffer(9898) := X"00031880";
        ram_buffer(9899) := X"02031821";
        ram_buffer(9900) := X"2A270006";
        ram_buffer(9901) := X"14E0001E";
        ram_buffer(9902) := X"AC730004";
        ram_buffer(9903) := X"24430047";
        ram_buffer(9904) := X"00031880";
        ram_buffer(9905) := X"02031821";
        ram_buffer(9906) := X"2A270007";
        ram_buffer(9907) := X"14E00018";
        ram_buffer(9908) := X"AC730004";
        ram_buffer(9909) := X"24430048";
        ram_buffer(9910) := X"00031880";
        ram_buffer(9911) := X"02031821";
        ram_buffer(9912) := X"2A270008";
        ram_buffer(9913) := X"14E00012";
        ram_buffer(9914) := X"AC730004";
        ram_buffer(9915) := X"24430049";
        ram_buffer(9916) := X"00031880";
        ram_buffer(9917) := X"02031821";
        ram_buffer(9918) := X"2A270009";
        ram_buffer(9919) := X"14E0000C";
        ram_buffer(9920) := X"AC730004";
        ram_buffer(9921) := X"2443004A";
        ram_buffer(9922) := X"00031880";
        ram_buffer(9923) := X"02031821";
        ram_buffer(9924) := X"2A31000A";
        ram_buffer(9925) := X"24420009";
        ram_buffer(9926) := X"16200005";
        ram_buffer(9927) := X"AC730004";
        ram_buffer(9928) := X"24420042";
        ram_buffer(9929) := X"00021080";
        ram_buffer(9930) := X"02021021";
        ram_buffer(9931) := X"AC530004";
        ram_buffer(9932) := X"00852021";
        ram_buffer(9933) := X"AE040108";
        ram_buffer(9934) := X"26730001";
        ram_buffer(9935) := X"0266102A";
        ram_buffer(9936) := X"1040001B";
        ram_buffer(9937) := X"26940004";
        ram_buffer(9938) := X"8E050108";
        ram_buffer(9939) := X"1000FF98";
        ram_buffer(9940) := X"00000000";
        ram_buffer(9941) := X"8C8300F0";
        ram_buffer(9942) := X"00000000";
        ram_buffer(9943) := X"8C650020";
        ram_buffer(9944) := X"8C64000C";
        ram_buffer(9945) := X"8C67001C";
        ram_buffer(9946) := X"14800002";
        ram_buffer(9947) := X"00A4001B";
        ram_buffer(9948) := X"0007000D";
        ram_buffer(9949) := X"AE050104";
        ram_buffer(9950) := X"24050008";
        ram_buffer(9951) := X"AE070100";
        ram_buffer(9952) := X"AC620034";
        ram_buffer(9953) := X"AC620038";
        ram_buffer(9954) := X"AC62003C";
        ram_buffer(9955) := X"AC650040";
        ram_buffer(9956) := X"00003010";
        ram_buffer(9957) := X"10C00002";
        ram_buffer(9958) := X"AC620044";
        ram_buffer(9959) := X"00C02021";
        ram_buffer(9960) := X"24020001";
        ram_buffer(9961) := X"AC640048";
        ram_buffer(9962) := X"AE020108";
        ram_buffer(9963) := X"AE00010C";
        ram_buffer(9964) := X"8E0300C4";
        ram_buffer(9965) := X"00000000";
        ram_buffer(9966) := X"1860000A";
        ram_buffer(9967) := X"00000000";
        ram_buffer(9968) := X"8E020100";
        ram_buffer(9969) := X"00000000";
        ram_buffer(9970) := X"00430018";
        ram_buffer(9971) := X"3C030001";
        ram_buffer(9972) := X"00001012";
        ram_buffer(9973) := X"0043182A";
        ram_buffer(9974) := X"10600013";
        ram_buffer(9975) := X"00000000";
        ram_buffer(9976) := X"AE0200C0";
        ram_buffer(9977) := X"8FBF0024";
        ram_buffer(9978) := X"8FB40020";
        ram_buffer(9979) := X"8FB3001C";
        ram_buffer(9980) := X"8FB20018";
        ram_buffer(9981) := X"8FB10014";
        ram_buffer(9982) := X"8FB00010";
        ram_buffer(9983) := X"03E00008";
        ram_buffer(9984) := X"27BD0028";
        ram_buffer(9985) := X"8E020000";
        ram_buffer(9986) := X"02002021";
        ram_buffer(9987) := X"8C430000";
        ram_buffer(9988) := X"00000000";
        ram_buffer(9989) := X"0060F809";
        ram_buffer(9990) := X"AC520014";
        ram_buffer(9991) := X"8E0600EC";
        ram_buffer(9992) := X"1000FF84";
        ram_buffer(9993) := X"00000000";
        ram_buffer(9994) := X"1000FFED";
        ram_buffer(9995) := X"3402FFFF";
        ram_buffer(9996) := X"8C830000";
        ram_buffer(9997) := X"24050018";
        ram_buffer(9998) := X"AC620018";
        ram_buffer(9999) := X"8C820000";
        ram_buffer(10000) := X"AC650014";
        ram_buffer(10001) := X"24030004";
        ram_buffer(10002) := X"AC43001C";
        ram_buffer(10003) := X"8C820000";
        ram_buffer(10004) := X"00000000";
        ram_buffer(10005) := X"8C420000";
        ram_buffer(10006) := X"00000000";
        ram_buffer(10007) := X"0040F809";
        ram_buffer(10008) := X"00000000";
        ram_buffer(10009) := X"1000FF41";
        ram_buffer(10010) := X"00000000";
        ram_buffer(10011) := X"8C8500A4";
        ram_buffer(10012) := X"00000000";
        ram_buffer(10013) := X"10A00043";
        ram_buffer(10014) := X"00801021";
        ram_buffer(10015) := X"8C830144";
        ram_buffer(10016) := X"00000000";
        ram_buffer(10017) := X"8C640020";
        ram_buffer(10018) := X"00000000";
        ram_buffer(10019) := X"00041880";
        ram_buffer(10020) := X"00042140";
        ram_buffer(10021) := X"00642021";
        ram_buffer(10022) := X"00A41821";
        ram_buffer(10023) := X"8C640000";
        ram_buffer(10024) := X"00000000";
        ram_buffer(10025) := X"1880002E";
        ram_buffer(10026) := X"AC4400EC";
        ram_buffer(10027) := X"8C660004";
        ram_buffer(10028) := X"8C47003C";
        ram_buffer(10029) := X"00062880";
        ram_buffer(10030) := X"00063100";
        ram_buffer(10031) := X"00C52823";
        ram_buffer(10032) := X"000530C0";
        ram_buffer(10033) := X"00C52823";
        ram_buffer(10034) := X"00E52821";
        ram_buffer(10035) := X"AC4500F0";
        ram_buffer(10036) := X"24050001";
        ram_buffer(10037) := X"10850022";
        ram_buffer(10038) := X"00000000";
        ram_buffer(10039) := X"8C660008";
        ram_buffer(10040) := X"00000000";
        ram_buffer(10041) := X"00062880";
        ram_buffer(10042) := X"00063100";
        ram_buffer(10043) := X"00C52823";
        ram_buffer(10044) := X"000530C0";
        ram_buffer(10045) := X"00C52823";
        ram_buffer(10046) := X"00E52821";
        ram_buffer(10047) := X"AC4500F4";
        ram_buffer(10048) := X"24050002";
        ram_buffer(10049) := X"10850016";
        ram_buffer(10050) := X"00000000";
        ram_buffer(10051) := X"8C66000C";
        ram_buffer(10052) := X"00000000";
        ram_buffer(10053) := X"00062880";
        ram_buffer(10054) := X"00063100";
        ram_buffer(10055) := X"00C52823";
        ram_buffer(10056) := X"000530C0";
        ram_buffer(10057) := X"00C52823";
        ram_buffer(10058) := X"00E52821";
        ram_buffer(10059) := X"AC4500F8";
        ram_buffer(10060) := X"24050003";
        ram_buffer(10061) := X"1085000A";
        ram_buffer(10062) := X"00000000";
        ram_buffer(10063) := X"8C650010";
        ram_buffer(10064) := X"00000000";
        ram_buffer(10065) := X"00052080";
        ram_buffer(10066) := X"00052900";
        ram_buffer(10067) := X"00A42023";
        ram_buffer(10068) := X"000428C0";
        ram_buffer(10069) := X"00A42023";
        ram_buffer(10070) := X"00E43821";
        ram_buffer(10071) := X"AC4700FC";
        ram_buffer(10072) := X"8C660014";
        ram_buffer(10073) := X"8C650018";
        ram_buffer(10074) := X"8C64001C";
        ram_buffer(10075) := X"8C630020";
        ram_buffer(10076) := X"AC460134";
        ram_buffer(10077) := X"AC450138";
        ram_buffer(10078) := X"AC44013C";
        ram_buffer(10079) := X"03E00008";
        ram_buffer(10080) := X"AC430140";
        ram_buffer(10081) := X"8C820034";
        ram_buffer(10082) := X"27BDFFE8";
        ram_buffer(10083) := X"28430005";
        ram_buffer(10084) := X"AFB00010";
        ram_buffer(10085) := X"AFBF0014";
        ram_buffer(10086) := X"1060001A";
        ram_buffer(10087) := X"00808021";
        ram_buffer(10088) := X"1840000F";
        ram_buffer(10089) := X"AE0200EC";
        ram_buffer(10090) := X"8E03003C";
        ram_buffer(10091) := X"24040001";
        ram_buffer(10092) := X"1044000B";
        ram_buffer(10093) := X"AE0300F0";
        ram_buffer(10094) := X"24640054";
        ram_buffer(10095) := X"AE0400F4";
        ram_buffer(10096) := X"24040002";
        ram_buffer(10097) := X"10440006";
        ram_buffer(10098) := X"246400A8";
        ram_buffer(10099) := X"AE0400F8";
        ram_buffer(10100) := X"24040003";
        ram_buffer(10101) := X"10440002";
        ram_buffer(10102) := X"246300FC";
        ram_buffer(10103) := X"AE0300FC";
        ram_buffer(10104) := X"8FBF0014";
        ram_buffer(10105) := X"2402003F";
        ram_buffer(10106) := X"AE000134";
        ram_buffer(10107) := X"AE020138";
        ram_buffer(10108) := X"AE00013C";
        ram_buffer(10109) := X"AE000140";
        ram_buffer(10110) := X"8FB00010";
        ram_buffer(10111) := X"03E00008";
        ram_buffer(10112) := X"27BD0018";
        ram_buffer(10113) := X"8C830000";
        ram_buffer(10114) := X"24050018";
        ram_buffer(10115) := X"AC620018";
        ram_buffer(10116) := X"8C820000";
        ram_buffer(10117) := X"AC650014";
        ram_buffer(10118) := X"24030004";
        ram_buffer(10119) := X"AC43001C";
        ram_buffer(10120) := X"8C820000";
        ram_buffer(10121) := X"00000000";
        ram_buffer(10122) := X"8C420000";
        ram_buffer(10123) := X"00000000";
        ram_buffer(10124) := X"0040F809";
        ram_buffer(10125) := X"00000000";
        ram_buffer(10126) := X"8E020034";
        ram_buffer(10127) := X"1000FFD8";
        ram_buffer(10128) := X"00000000";
        ram_buffer(10129) := X"27BDFFE0";
        ram_buffer(10130) := X"AFB10018";
        ram_buffer(10131) := X"8C910144";
        ram_buffer(10132) := X"24030001";
        ram_buffer(10133) := X"8E220014";
        ram_buffer(10134) := X"AFB00014";
        ram_buffer(10135) := X"AFBF001C";
        ram_buffer(10136) := X"10430060";
        ram_buffer(10137) := X"00808021";
        ram_buffer(10138) := X"10400035";
        ram_buffer(10139) := X"24030002";
        ram_buffer(10140) := X"1443002B";
        ram_buffer(10141) := X"2405002F";
        ram_buffer(10142) := X"8E0200B0";
        ram_buffer(10143) := X"00000000";
        ram_buffer(10144) := X"10400092";
        ram_buffer(10145) := X"00000000";
        ram_buffer(10146) := X"8E020164";
        ram_buffer(10147) := X"02002021";
        ram_buffer(10148) := X"8C420000";
        ram_buffer(10149) := X"00000000";
        ram_buffer(10150) := X"0040F809";
        ram_buffer(10151) := X"00002821";
        ram_buffer(10152) := X"8E020150";
        ram_buffer(10153) := X"24050002";
        ram_buffer(10154) := X"8C420000";
        ram_buffer(10155) := X"00000000";
        ram_buffer(10156) := X"0040F809";
        ram_buffer(10157) := X"02002021";
        ram_buffer(10158) := X"8E220020";
        ram_buffer(10159) := X"00000000";
        ram_buffer(10160) := X"1040007A";
        ram_buffer(10161) := X"00000000";
        ram_buffer(10162) := X"8E020154";
        ram_buffer(10163) := X"00000000";
        ram_buffer(10164) := X"8C42000C";
        ram_buffer(10165) := X"00000000";
        ram_buffer(10166) := X"0040F809";
        ram_buffer(10167) := X"02002021";
        ram_buffer(10168) := X"AE20000C";
        ram_buffer(10169) := X"8E24001C";
        ram_buffer(10170) := X"8E250018";
        ram_buffer(10171) := X"2482FFFF";
        ram_buffer(10172) := X"00451026";
        ram_buffer(10173) := X"8E030008";
        ram_buffer(10174) := X"2C420001";
        ram_buffer(10175) := X"10600003";
        ram_buffer(10176) := X"AE220010";
        ram_buffer(10177) := X"AC65000C";
        ram_buffer(10178) := X"AC640010";
        ram_buffer(10179) := X"8FBF001C";
        ram_buffer(10180) := X"8FB10018";
        ram_buffer(10181) := X"8FB00014";
        ram_buffer(10182) := X"03E00008";
        ram_buffer(10183) := X"27BD0020";
        ram_buffer(10184) := X"8C820000";
        ram_buffer(10185) := X"00000000";
        ram_buffer(10186) := X"8C430000";
        ram_buffer(10187) := X"00000000";
        ram_buffer(10188) := X"0060F809";
        ram_buffer(10189) := X"AC450014";
        ram_buffer(10190) := X"1000FFEA";
        ram_buffer(10191) := X"00000000";
        ram_buffer(10192) := X"0C02271B";
        ram_buffer(10193) := X"00000000";
        ram_buffer(10194) := X"0C02264C";
        ram_buffer(10195) := X"02002021";
        ram_buffer(10196) := X"8E0200A8";
        ram_buffer(10197) := X"00000000";
        ram_buffer(10198) := X"10400040";
        ram_buffer(10199) := X"00000000";
        ram_buffer(10200) := X"8E020160";
        ram_buffer(10201) := X"00000000";
        ram_buffer(10202) := X"8C420000";
        ram_buffer(10203) := X"00000000";
        ram_buffer(10204) := X"0040F809";
        ram_buffer(10205) := X"02002021";
        ram_buffer(10206) := X"8E020164";
        ram_buffer(10207) := X"8E0500B0";
        ram_buffer(10208) := X"8C420000";
        ram_buffer(10209) := X"00000000";
        ram_buffer(10210) := X"0040F809";
        ram_buffer(10211) := X"02002021";
        ram_buffer(10212) := X"8E22001C";
        ram_buffer(10213) := X"8E030150";
        ram_buffer(10214) := X"28420002";
        ram_buffer(10215) := X"8C630000";
        ram_buffer(10216) := X"14400002";
        ram_buffer(10217) := X"00002821";
        ram_buffer(10218) := X"24050003";
        ram_buffer(10219) := X"0060F809";
        ram_buffer(10220) := X"02002021";
        ram_buffer(10221) := X"8E020148";
        ram_buffer(10222) := X"00002821";
        ram_buffer(10223) := X"8C420000";
        ram_buffer(10224) := X"00000000";
        ram_buffer(10225) := X"0040F809";
        ram_buffer(10226) := X"02002021";
        ram_buffer(10227) := X"8E0200B0";
        ram_buffer(10228) := X"00000000";
        ram_buffer(10229) := X"1440001F";
        ram_buffer(10230) := X"24020001";
        ram_buffer(10231) := X"1000FFC1";
        ram_buffer(10232) := X"AE22000C";
        ram_buffer(10233) := X"0C02271B";
        ram_buffer(10234) := X"00000000";
        ram_buffer(10235) := X"0C02264C";
        ram_buffer(10236) := X"02002021";
        ram_buffer(10237) := X"8E020134";
        ram_buffer(10238) := X"00000000";
        ram_buffer(10239) := X"14400009";
        ram_buffer(10240) := X"00000000";
        ram_buffer(10241) := X"8E02013C";
        ram_buffer(10242) := X"00000000";
        ram_buffer(10243) := X"10400005";
        ram_buffer(10244) := X"00000000";
        ram_buffer(10245) := X"8E0200AC";
        ram_buffer(10246) := X"00000000";
        ram_buffer(10247) := X"10400031";
        ram_buffer(10248) := X"24030002";
        ram_buffer(10249) := X"8E020164";
        ram_buffer(10250) := X"02002021";
        ram_buffer(10251) := X"8C420000";
        ram_buffer(10252) := X"00000000";
        ram_buffer(10253) := X"0040F809";
        ram_buffer(10254) := X"24050001";
        ram_buffer(10255) := X"8E020150";
        ram_buffer(10256) := X"24050002";
        ram_buffer(10257) := X"8C420000";
        ram_buffer(10258) := X"00000000";
        ram_buffer(10259) := X"0040F809";
        ram_buffer(10260) := X"02002021";
        ram_buffer(10261) := X"1000FFA3";
        ram_buffer(10262) := X"AE20000C";
        ram_buffer(10263) := X"8E020158";
        ram_buffer(10264) := X"00000000";
        ram_buffer(10265) := X"8C420000";
        ram_buffer(10266) := X"00000000";
        ram_buffer(10267) := X"0040F809";
        ram_buffer(10268) := X"02002021";
        ram_buffer(10269) := X"8E02015C";
        ram_buffer(10270) := X"00000000";
        ram_buffer(10271) := X"8C420000";
        ram_buffer(10272) := X"00000000";
        ram_buffer(10273) := X"0040F809";
        ram_buffer(10274) := X"02002021";
        ram_buffer(10275) := X"8E02014C";
        ram_buffer(10276) := X"00002821";
        ram_buffer(10277) := X"8C420000";
        ram_buffer(10278) := X"00000000";
        ram_buffer(10279) := X"0040F809";
        ram_buffer(10280) := X"02002021";
        ram_buffer(10281) := X"1000FFAE";
        ram_buffer(10282) := X"00000000";
        ram_buffer(10283) := X"8E020154";
        ram_buffer(10284) := X"00000000";
        ram_buffer(10285) := X"8C420008";
        ram_buffer(10286) := X"00000000";
        ram_buffer(10287) := X"0040F809";
        ram_buffer(10288) := X"02002021";
        ram_buffer(10289) := X"1000FF80";
        ram_buffer(10290) := X"00000000";
        ram_buffer(10291) := X"0C02271B";
        ram_buffer(10292) := X"02002021";
        ram_buffer(10293) := X"0C02264C";
        ram_buffer(10294) := X"02002021";
        ram_buffer(10295) := X"1000FF6A";
        ram_buffer(10296) := X"00000000";
        ram_buffer(10297) := X"8E220018";
        ram_buffer(10298) := X"00000000";
        ram_buffer(10299) := X"24420001";
        ram_buffer(10300) := X"AE230014";
        ram_buffer(10301) := X"1000FF60";
        ram_buffer(10302) := X"AE220018";
        ram_buffer(10303) := X"8C820004";
        ram_buffer(10304) := X"27BDFFD0";
        ram_buffer(10305) := X"8C420000";
        ram_buffer(10306) := X"24060024";
        ram_buffer(10307) := X"AFB40020";
        ram_buffer(10308) := X"AFB3001C";
        ram_buffer(10309) := X"AFB00010";
        ram_buffer(10310) := X"AFBF002C";
        ram_buffer(10311) := X"AFB60028";
        ram_buffer(10312) := X"AFB50024";
        ram_buffer(10313) := X"AFB20018";
        ram_buffer(10314) := X"AFB10014";
        ram_buffer(10315) := X"00A0A021";
        ram_buffer(10316) := X"24050001";
        ram_buffer(10317) := X"0040F809";
        ram_buffer(10318) := X"00808021";
        ram_buffer(10319) := X"3C031009";
        ram_buffer(10320) := X"00409821";
        ram_buffer(10321) := X"24639E44";
        ram_buffer(10322) := X"8E02001C";
        ram_buffer(10323) := X"AE130144";
        ram_buffer(10324) := X"AE630000";
        ram_buffer(10325) := X"3C031009";
        ram_buffer(10326) := X"2463981C";
        ram_buffer(10327) := X"AE630004";
        ram_buffer(10328) := X"3C031009";
        ram_buffer(10329) := X"2463985C";
        ram_buffer(10330) := X"AE630008";
        ram_buffer(10331) := X"10400005";
        ram_buffer(10332) := X"AE600010";
        ram_buffer(10333) := X"8E030018";
        ram_buffer(10334) := X"00000000";
        ram_buffer(10335) := X"146000BD";
        ram_buffer(10336) := X"00000000";
        ram_buffer(10337) := X"8E020000";
        ram_buffer(10338) := X"2404001F";
        ram_buffer(10339) := X"8C430000";
        ram_buffer(10340) := X"AC440014";
        ram_buffer(10341) := X"0060F809";
        ram_buffer(10342) := X"02002021";
        ram_buffer(10343) := X"8E02001C";
        ram_buffer(10344) := X"3403FFDD";
        ram_buffer(10345) := X"0043102A";
        ram_buffer(10346) := X"10400046";
        ram_buffer(10347) := X"00000000";
        ram_buffer(10348) := X"8E020018";
        ram_buffer(10349) := X"00000000";
        ram_buffer(10350) := X"0043102A";
        ram_buffer(10351) := X"10400041";
        ram_buffer(10352) := X"00000000";
        ram_buffer(10353) := X"8E020030";
        ram_buffer(10354) := X"24030008";
        ram_buffer(10355) := X"1043000A";
        ram_buffer(10356) := X"00000000";
        ram_buffer(10357) := X"8E030000";
        ram_buffer(10358) := X"2404000D";
        ram_buffer(10359) := X"AC620018";
        ram_buffer(10360) := X"8E020000";
        ram_buffer(10361) := X"AC640014";
        ram_buffer(10362) := X"8C420000";
        ram_buffer(10363) := X"00000000";
        ram_buffer(10364) := X"0040F809";
        ram_buffer(10365) := X"02002021";
        ram_buffer(10366) := X"8E080034";
        ram_buffer(10367) := X"00000000";
        ram_buffer(10368) := X"2902000B";
        ram_buffer(10369) := X"104000AF";
        ram_buffer(10370) := X"00000000";
        ram_buffer(10371) := X"24020001";
        ram_buffer(10372) := X"AE0200E0";
        ram_buffer(10373) := X"AE0200E4";
        ram_buffer(10374) := X"8E11003C";
        ram_buffer(10375) := X"190000B9";
        ram_buffer(10376) := X"24060001";
        ram_buffer(10377) := X"24050001";
        ram_buffer(10378) := X"0000A821";
        ram_buffer(10379) := X"10000012";
        ram_buffer(10380) := X"24120010";
        ram_buffer(10381) := X"8E27000C";
        ram_buffer(10382) := X"00000000";
        ram_buffer(10383) := X"24E3FFFF";
        ram_buffer(10384) := X"2C630004";
        ram_buffer(10385) := X"10600012";
        ram_buffer(10386) := X"00000000";
        ram_buffer(10387) := X"00A2182A";
        ram_buffer(10388) := X"00C7482A";
        ram_buffer(10389) := X"10600002";
        ram_buffer(10390) := X"02A8202A";
        ram_buffer(10391) := X"00402821";
        ram_buffer(10392) := X"11200002";
        ram_buffer(10393) := X"AE0500E0";
        ram_buffer(10394) := X"00E03021";
        ram_buffer(10395) := X"AE0600E4";
        ram_buffer(10396) := X"1080001F";
        ram_buffer(10397) := X"26310054";
        ram_buffer(10398) := X"8E220008";
        ram_buffer(10399) := X"26B50001";
        ram_buffer(10400) := X"2443FFFF";
        ram_buffer(10401) := X"2C630004";
        ram_buffer(10402) := X"1460FFEA";
        ram_buffer(10403) := X"02002021";
        ram_buffer(10404) := X"8E020000";
        ram_buffer(10405) := X"00000000";
        ram_buffer(10406) := X"8C430000";
        ram_buffer(10407) := X"00000000";
        ram_buffer(10408) := X"0060F809";
        ram_buffer(10409) := X"AC520014";
        ram_buffer(10410) := X"8E220008";
        ram_buffer(10411) := X"8E27000C";
        ram_buffer(10412) := X"8E0500E0";
        ram_buffer(10413) := X"8E0600E4";
        ram_buffer(10414) := X"8E080034";
        ram_buffer(10415) := X"1000FFE4";
        ram_buffer(10416) := X"00A2182A";
        ram_buffer(10417) := X"8E020000";
        ram_buffer(10418) := X"3403FFDC";
        ram_buffer(10419) := X"AC430018";
        ram_buffer(10420) := X"8E030000";
        ram_buffer(10421) := X"24040028";
        ram_buffer(10422) := X"8C630000";
        ram_buffer(10423) := X"AC440014";
        ram_buffer(10424) := X"0060F809";
        ram_buffer(10425) := X"02002021";
        ram_buffer(10426) := X"1000FFB6";
        ram_buffer(10427) := X"00000000";
        ram_buffer(10428) := X"8E11003C";
        ram_buffer(10429) := X"19000085";
        ram_buffer(10430) := X"00000000";
        ram_buffer(10431) := X"00009021";
        ram_buffer(10432) := X"24160008";
        ram_buffer(10433) := X"10000002";
        ram_buffer(10434) := X"24150001";
        ram_buffer(10435) := X"8E0500E0";
        ram_buffer(10436) := X"AE320004";
        ram_buffer(10437) := X"AE360024";
        ram_buffer(10438) := X"8E220008";
        ram_buffer(10439) := X"8E040018";
        ram_buffer(10440) := X"000528C0";
        ram_buffer(10441) := X"00820018";
        ram_buffer(10442) := X"26310054";
        ram_buffer(10443) := X"00002012";
        ram_buffer(10444) := X"0C0264AB";
        ram_buffer(10445) := X"26520001";
        ram_buffer(10446) := X"AE22FFC8";
        ram_buffer(10447) := X"8E04001C";
        ram_buffer(10448) := X"8E22FFB8";
        ram_buffer(10449) := X"8E0500E4";
        ram_buffer(10450) := X"00820018";
        ram_buffer(10451) := X"00002012";
        ram_buffer(10452) := X"0C0264AB";
        ram_buffer(10453) := X"000528C0";
        ram_buffer(10454) := X"AE22FFCC";
        ram_buffer(10455) := X"8E040018";
        ram_buffer(10456) := X"8E22FFB4";
        ram_buffer(10457) := X"8E0500E0";
        ram_buffer(10458) := X"00820018";
        ram_buffer(10459) := X"00002012";
        ram_buffer(10460) := X"0C0264AB";
        ram_buffer(10461) := X"00000000";
        ram_buffer(10462) := X"AE22FFD4";
        ram_buffer(10463) := X"8E04001C";
        ram_buffer(10464) := X"8E22FFB8";
        ram_buffer(10465) := X"8E0500E4";
        ram_buffer(10466) := X"00820018";
        ram_buffer(10467) := X"00002012";
        ram_buffer(10468) := X"0C0264AB";
        ram_buffer(10469) := X"00000000";
        ram_buffer(10470) := X"AE22FFD8";
        ram_buffer(10471) := X"AE35FFDC";
        ram_buffer(10472) := X"8E020034";
        ram_buffer(10473) := X"00000000";
        ram_buffer(10474) := X"0242102A";
        ram_buffer(10475) := X"1440FFD7";
        ram_buffer(10476) := X"00000000";
        ram_buffer(10477) := X"8E0500E4";
        ram_buffer(10478) := X"00000000";
        ram_buffer(10479) := X"000528C0";
        ram_buffer(10480) := X"8E04001C";
        ram_buffer(10481) := X"0C0264AB";
        ram_buffer(10482) := X"00000000";
        ram_buffer(10483) := X"8E0300A4";
        ram_buffer(10484) := X"00000000";
        ram_buffer(10485) := X"1060000F";
        ram_buffer(10486) := X"AE0200E8";
        ram_buffer(10487) := X"0C0222CD";
        ram_buffer(10488) := X"02002021";
        ram_buffer(10489) := X"8E0200DC";
        ram_buffer(10490) := X"00000000";
        ram_buffer(10491) := X"1040000C";
        ram_buffer(10492) := X"24020001";
        ram_buffer(10493) := X"1680002F";
        ram_buffer(10494) := X"AE0200B0";
        ram_buffer(10495) := X"AE600014";
        ram_buffer(10496) := X"AE600020";
        ram_buffer(10497) := X"AE600018";
        ram_buffer(10498) := X"8E0200A0";
        ram_buffer(10499) := X"1000000E";
        ram_buffer(10500) := X"00021040";
        ram_buffer(10501) := X"24020001";
        ram_buffer(10502) := X"AE0000DC";
        ram_buffer(10503) := X"AE0200A0";
        ram_buffer(10504) := X"8E0200B0";
        ram_buffer(10505) := X"1280001D";
        ram_buffer(10506) := X"00000000";
        ram_buffer(10507) := X"14400021";
        ram_buffer(10508) := X"24020001";
        ram_buffer(10509) := X"24020002";
        ram_buffer(10510) := X"AE620014";
        ram_buffer(10511) := X"AE600020";
        ram_buffer(10512) := X"AE600018";
        ram_buffer(10513) := X"8E0200A0";
        ram_buffer(10514) := X"8FBF002C";
        ram_buffer(10515) := X"AE62001C";
        ram_buffer(10516) := X"8FB60028";
        ram_buffer(10517) := X"8FB50024";
        ram_buffer(10518) := X"8FB40020";
        ram_buffer(10519) := X"8FB3001C";
        ram_buffer(10520) := X"8FB20018";
        ram_buffer(10521) := X"8FB10014";
        ram_buffer(10522) := X"8FB00010";
        ram_buffer(10523) := X"03E00008";
        ram_buffer(10524) := X"27BD0030";
        ram_buffer(10525) := X"8E030034";
        ram_buffer(10526) := X"00000000";
        ram_buffer(10527) := X"1860FF41";
        ram_buffer(10528) := X"00000000";
        ram_buffer(10529) := X"8E030020";
        ram_buffer(10530) := X"00000000";
        ram_buffer(10531) := X"1C60FF45";
        ram_buffer(10532) := X"3403FFDD";
        ram_buffer(10533) := X"1000FF3B";
        ram_buffer(10534) := X"00000000";
        ram_buffer(10535) := X"AE600014";
        ram_buffer(10536) := X"AE600020";
        ram_buffer(10537) := X"1040FFE7";
        ram_buffer(10538) := X"AE600018";
        ram_buffer(10539) := X"1000FFD6";
        ram_buffer(10540) := X"00000000";
        ram_buffer(10541) := X"AE620014";
        ram_buffer(10542) := X"AE600020";
        ram_buffer(10543) := X"1000FFD2";
        ram_buffer(10544) := X"AE600018";
        ram_buffer(10545) := X"8E020000";
        ram_buffer(10546) := X"24040018";
        ram_buffer(10547) := X"AC480018";
        ram_buffer(10548) := X"8E030000";
        ram_buffer(10549) := X"AC440014";
        ram_buffer(10550) := X"2402000A";
        ram_buffer(10551) := X"AC62001C";
        ram_buffer(10552) := X"8E020000";
        ram_buffer(10553) := X"00000000";
        ram_buffer(10554) := X"8C420000";
        ram_buffer(10555) := X"00000000";
        ram_buffer(10556) := X"0040F809";
        ram_buffer(10557) := X"02002021";
        ram_buffer(10558) := X"8E080034";
        ram_buffer(10559) := X"1000FF44";
        ram_buffer(10560) := X"24020001";
        ram_buffer(10561) := X"1000FFAE";
        ram_buffer(10562) := X"24050008";
        ram_buffer(10563) := X"1000FFAC";
        ram_buffer(10564) := X"000628C0";
        ram_buffer(10565) := X"8C820014";
        ram_buffer(10566) := X"27BDFFE8";
        ram_buffer(10567) := X"8C430000";
        ram_buffer(10568) := X"AFB00010";
        ram_buffer(10569) := X"24650001";
        ram_buffer(10570) := X"AFBF0014";
        ram_buffer(10571) := X"AC450000";
        ram_buffer(10572) := X"2405FFFF";
        ram_buffer(10573) := X"A0650000";
        ram_buffer(10574) := X"8C430004";
        ram_buffer(10575) := X"00808021";
        ram_buffer(10576) := X"2463FFFF";
        ram_buffer(10577) := X"10600012";
        ram_buffer(10578) := X"AC430004";
        ram_buffer(10579) := X"8E020014";
        ram_buffer(10580) := X"00000000";
        ram_buffer(10581) := X"8C430000";
        ram_buffer(10582) := X"00000000";
        ram_buffer(10583) := X"24640001";
        ram_buffer(10584) := X"AC440000";
        ram_buffer(10585) := X"2404FFD9";
        ram_buffer(10586) := X"A0640000";
        ram_buffer(10587) := X"8C430004";
        ram_buffer(10588) := X"00000000";
        ram_buffer(10589) := X"2463FFFF";
        ram_buffer(10590) := X"1060001E";
        ram_buffer(10591) := X"AC430004";
        ram_buffer(10592) := X"8FBF0014";
        ram_buffer(10593) := X"8FB00010";
        ram_buffer(10594) := X"03E00008";
        ram_buffer(10595) := X"27BD0018";
        ram_buffer(10596) := X"8C42000C";
        ram_buffer(10597) := X"00000000";
        ram_buffer(10598) := X"0040F809";
        ram_buffer(10599) := X"00000000";
        ram_buffer(10600) := X"1440FFEA";
        ram_buffer(10601) := X"24040016";
        ram_buffer(10602) := X"8E020000";
        ram_buffer(10603) := X"00000000";
        ram_buffer(10604) := X"8C430000";
        ram_buffer(10605) := X"AC440014";
        ram_buffer(10606) := X"0060F809";
        ram_buffer(10607) := X"02002021";
        ram_buffer(10608) := X"8E020014";
        ram_buffer(10609) := X"00000000";
        ram_buffer(10610) := X"8C430000";
        ram_buffer(10611) := X"00000000";
        ram_buffer(10612) := X"24640001";
        ram_buffer(10613) := X"AC440000";
        ram_buffer(10614) := X"2404FFD9";
        ram_buffer(10615) := X"A0640000";
        ram_buffer(10616) := X"8C430004";
        ram_buffer(10617) := X"00000000";
        ram_buffer(10618) := X"2463FFFF";
        ram_buffer(10619) := X"1460FFE4";
        ram_buffer(10620) := X"AC430004";
        ram_buffer(10621) := X"8C42000C";
        ram_buffer(10622) := X"00000000";
        ram_buffer(10623) := X"0040F809";
        ram_buffer(10624) := X"02002021";
        ram_buffer(10625) := X"1440FFDE";
        ram_buffer(10626) := X"24030016";
        ram_buffer(10627) := X"8E020000";
        ram_buffer(10628) := X"8FBF0014";
        ram_buffer(10629) := X"8C590000";
        ram_buffer(10630) := X"02002021";
        ram_buffer(10631) := X"8FB00010";
        ram_buffer(10632) := X"AC430014";
        ram_buffer(10633) := X"03200008";
        ram_buffer(10634) := X"27BD0018";
        ram_buffer(10635) := X"3402FFFE";
        ram_buffer(10636) := X"00E2102B";
        ram_buffer(10637) := X"14400003";
        ram_buffer(10638) := X"00000000";
        ram_buffer(10639) := X"03E00008";
        ram_buffer(10640) := X"00000000";
        ram_buffer(10641) := X"8C820014";
        ram_buffer(10642) := X"27BDFFD0";
        ram_buffer(10643) := X"8C430000";
        ram_buffer(10644) := X"AFB10020";
        ram_buffer(10645) := X"00C08821";
        ram_buffer(10646) := X"24660001";
        ram_buffer(10647) := X"AFB20024";
        ram_buffer(10648) := X"AFB0001C";
        ram_buffer(10649) := X"AFBF002C";
        ram_buffer(10650) := X"AFB30028";
        ram_buffer(10651) := X"AC460000";
        ram_buffer(10652) := X"2406FFFF";
        ram_buffer(10653) := X"A0660000";
        ram_buffer(10654) := X"8C430004";
        ram_buffer(10655) := X"00E08021";
        ram_buffer(10656) := X"2463FFFF";
        ram_buffer(10657) := X"00809021";
        ram_buffer(10658) := X"10600076";
        ram_buffer(10659) := X"AC430004";
        ram_buffer(10660) := X"8E420014";
        ram_buffer(10661) := X"00000000";
        ram_buffer(10662) := X"8C430000";
        ram_buffer(10663) := X"00000000";
        ram_buffer(10664) := X"24640001";
        ram_buffer(10665) := X"AC440000";
        ram_buffer(10666) := X"A0650000";
        ram_buffer(10667) := X"8C430004";
        ram_buffer(10668) := X"00000000";
        ram_buffer(10669) := X"2463FFFF";
        ram_buffer(10670) := X"1060005C";
        ram_buffer(10671) := X"AC430004";
        ram_buffer(10672) := X"8E420014";
        ram_buffer(10673) := X"26130002";
        ram_buffer(10674) := X"8C430000";
        ram_buffer(10675) := X"00132203";
        ram_buffer(10676) := X"24650001";
        ram_buffer(10677) := X"AC450000";
        ram_buffer(10678) := X"A0640000";
        ram_buffer(10679) := X"8C430004";
        ram_buffer(10680) := X"00000000";
        ram_buffer(10681) := X"2463FFFF";
        ram_buffer(10682) := X"10600042";
        ram_buffer(10683) := X"AC430004";
        ram_buffer(10684) := X"8E420014";
        ram_buffer(10685) := X"00000000";
        ram_buffer(10686) := X"8C430000";
        ram_buffer(10687) := X"00000000";
        ram_buffer(10688) := X"24640001";
        ram_buffer(10689) := X"AC440000";
        ram_buffer(10690) := X"A0730000";
        ram_buffer(10691) := X"8C430004";
        ram_buffer(10692) := X"00000000";
        ram_buffer(10693) := X"2463FFFF";
        ram_buffer(10694) := X"10600028";
        ram_buffer(10695) := X"AC430004";
        ram_buffer(10696) := X"1200000F";
        ram_buffer(10697) := X"24130016";
        ram_buffer(10698) := X"8E420014";
        ram_buffer(10699) := X"92240000";
        ram_buffer(10700) := X"8C430000";
        ram_buffer(10701) := X"2610FFFF";
        ram_buffer(10702) := X"24650001";
        ram_buffer(10703) := X"AC450000";
        ram_buffer(10704) := X"A0640000";
        ram_buffer(10705) := X"8C430004";
        ram_buffer(10706) := X"26310001";
        ram_buffer(10707) := X"2463FFFF";
        ram_buffer(10708) := X"1060000A";
        ram_buffer(10709) := X"AC430004";
        ram_buffer(10710) := X"1600FFF3";
        ram_buffer(10711) := X"00000000";
        ram_buffer(10712) := X"8FBF002C";
        ram_buffer(10713) := X"8FB30028";
        ram_buffer(10714) := X"8FB20024";
        ram_buffer(10715) := X"8FB10020";
        ram_buffer(10716) := X"8FB0001C";
        ram_buffer(10717) := X"03E00008";
        ram_buffer(10718) := X"27BD0030";
        ram_buffer(10719) := X"8C42000C";
        ram_buffer(10720) := X"00000000";
        ram_buffer(10721) := X"0040F809";
        ram_buffer(10722) := X"02402021";
        ram_buffer(10723) := X"1440FFF2";
        ram_buffer(10724) := X"02402021";
        ram_buffer(10725) := X"8E420000";
        ram_buffer(10726) := X"00000000";
        ram_buffer(10727) := X"8C430000";
        ram_buffer(10728) := X"00000000";
        ram_buffer(10729) := X"0060F809";
        ram_buffer(10730) := X"AC530014";
        ram_buffer(10731) := X"1600FFDE";
        ram_buffer(10732) := X"00000000";
        ram_buffer(10733) := X"1000FFEA";
        ram_buffer(10734) := X"00000000";
        ram_buffer(10735) := X"8C42000C";
        ram_buffer(10736) := X"00000000";
        ram_buffer(10737) := X"0040F809";
        ram_buffer(10738) := X"02402021";
        ram_buffer(10739) := X"1440FFD4";
        ram_buffer(10740) := X"24040016";
        ram_buffer(10741) := X"8E420000";
        ram_buffer(10742) := X"00000000";
        ram_buffer(10743) := X"8C430000";
        ram_buffer(10744) := X"AC440014";
        ram_buffer(10745) := X"0060F809";
        ram_buffer(10746) := X"02402021";
        ram_buffer(10747) := X"1000FFCC";
        ram_buffer(10748) := X"00000000";
        ram_buffer(10749) := X"8C42000C";
        ram_buffer(10750) := X"00000000";
        ram_buffer(10751) := X"0040F809";
        ram_buffer(10752) := X"02402021";
        ram_buffer(10753) := X"1440FFBA";
        ram_buffer(10754) := X"24040016";
        ram_buffer(10755) := X"8E420000";
        ram_buffer(10756) := X"00000000";
        ram_buffer(10757) := X"8C430000";
        ram_buffer(10758) := X"AC440014";
        ram_buffer(10759) := X"0060F809";
        ram_buffer(10760) := X"02402021";
        ram_buffer(10761) := X"1000FFB2";
        ram_buffer(10762) := X"00000000";
        ram_buffer(10763) := X"8C42000C";
        ram_buffer(10764) := X"00000000";
        ram_buffer(10765) := X"0040F809";
        ram_buffer(10766) := X"02402021";
        ram_buffer(10767) := X"1440FFA0";
        ram_buffer(10768) := X"24040016";
        ram_buffer(10769) := X"8E420000";
        ram_buffer(10770) := X"00000000";
        ram_buffer(10771) := X"8C430000";
        ram_buffer(10772) := X"AC440014";
        ram_buffer(10773) := X"0060F809";
        ram_buffer(10774) := X"02402021";
        ram_buffer(10775) := X"1000FF98";
        ram_buffer(10776) := X"00000000";
        ram_buffer(10777) := X"8C42000C";
        ram_buffer(10778) := X"00000000";
        ram_buffer(10779) := X"0040F809";
        ram_buffer(10780) := X"AFA50010";
        ram_buffer(10781) := X"8FA50010";
        ram_buffer(10782) := X"1440FF85";
        ram_buffer(10783) := X"24040016";
        ram_buffer(10784) := X"8E420000";
        ram_buffer(10785) := X"00000000";
        ram_buffer(10786) := X"8C430000";
        ram_buffer(10787) := X"AC440014";
        ram_buffer(10788) := X"0060F809";
        ram_buffer(10789) := X"02402021";
        ram_buffer(10790) := X"8FA50010";
        ram_buffer(10791) := X"1000FF7C";
        ram_buffer(10792) := X"00000000";
        ram_buffer(10793) := X"8C820014";
        ram_buffer(10794) := X"27BDFFD8";
        ram_buffer(10795) := X"8C430000";
        ram_buffer(10796) := X"AFB10018";
        ram_buffer(10797) := X"00A08821";
        ram_buffer(10798) := X"24650001";
        ram_buffer(10799) := X"AFB00014";
        ram_buffer(10800) := X"AFBF0024";
        ram_buffer(10801) := X"AFB30020";
        ram_buffer(10802) := X"AFB2001C";
        ram_buffer(10803) := X"AC450000";
        ram_buffer(10804) := X"2405FFFF";
        ram_buffer(10805) := X"A0650000";
        ram_buffer(10806) := X"8C430004";
        ram_buffer(10807) := X"00808021";
        ram_buffer(10808) := X"2463FFFF";
        ram_buffer(10809) := X"1060017B";
        ram_buffer(10810) := X"AC430004";
        ram_buffer(10811) := X"8E020014";
        ram_buffer(10812) := X"00000000";
        ram_buffer(10813) := X"8C430000";
        ram_buffer(10814) := X"00000000";
        ram_buffer(10815) := X"24640001";
        ram_buffer(10816) := X"AC440000";
        ram_buffer(10817) := X"A0710000";
        ram_buffer(10818) := X"8C430004";
        ram_buffer(10819) := X"00000000";
        ram_buffer(10820) := X"2463FFFF";
        ram_buffer(10821) := X"10600187";
        ram_buffer(10822) := X"AC430004";
        ram_buffer(10823) := X"8E110034";
        ram_buffer(10824) := X"8E030014";
        ram_buffer(10825) := X"00111040";
        ram_buffer(10826) := X"8C640000";
        ram_buffer(10827) := X"00518821";
        ram_buffer(10828) := X"26310008";
        ram_buffer(10829) := X"00111203";
        ram_buffer(10830) := X"24850001";
        ram_buffer(10831) := X"AC650000";
        ram_buffer(10832) := X"A0820000";
        ram_buffer(10833) := X"8C620004";
        ram_buffer(10834) := X"00000000";
        ram_buffer(10835) := X"2442FFFF";
        ram_buffer(10836) := X"10400194";
        ram_buffer(10837) := X"AC620004";
        ram_buffer(10838) := X"8E020014";
        ram_buffer(10839) := X"00000000";
        ram_buffer(10840) := X"8C430000";
        ram_buffer(10841) := X"00000000";
        ram_buffer(10842) := X"24640001";
        ram_buffer(10843) := X"AC440000";
        ram_buffer(10844) := X"A0710000";
        ram_buffer(10845) := X"8C430004";
        ram_buffer(10846) := X"00000000";
        ram_buffer(10847) := X"2463FFFF";
        ram_buffer(10848) := X"1060017A";
        ram_buffer(10849) := X"AC430004";
        ram_buffer(10850) := X"8E02001C";
        ram_buffer(10851) := X"3C030001";
        ram_buffer(10852) := X"0043102A";
        ram_buffer(10853) := X"1040008E";
        ram_buffer(10854) := X"00000000";
        ram_buffer(10855) := X"8E020018";
        ram_buffer(10856) := X"00000000";
        ram_buffer(10857) := X"0043102A";
        ram_buffer(10858) := X"10400089";
        ram_buffer(10859) := X"00000000";
        ram_buffer(10860) := X"8E020014";
        ram_buffer(10861) := X"8E040030";
        ram_buffer(10862) := X"8C430000";
        ram_buffer(10863) := X"00000000";
        ram_buffer(10864) := X"24650001";
        ram_buffer(10865) := X"AC450000";
        ram_buffer(10866) := X"A0640000";
        ram_buffer(10867) := X"8C430004";
        ram_buffer(10868) := X"00000000";
        ram_buffer(10869) := X"2463FFFF";
        ram_buffer(10870) := X"10600092";
        ram_buffer(10871) := X"AC430004";
        ram_buffer(10872) := X"8E020014";
        ram_buffer(10873) := X"8E11001C";
        ram_buffer(10874) := X"8C430000";
        ram_buffer(10875) := X"00112203";
        ram_buffer(10876) := X"24650001";
        ram_buffer(10877) := X"AC450000";
        ram_buffer(10878) := X"A0640000";
        ram_buffer(10879) := X"8C430004";
        ram_buffer(10880) := X"00000000";
        ram_buffer(10881) := X"2463FFFF";
        ram_buffer(10882) := X"1060009E";
        ram_buffer(10883) := X"AC430004";
        ram_buffer(10884) := X"8E020014";
        ram_buffer(10885) := X"00000000";
        ram_buffer(10886) := X"8C430000";
        ram_buffer(10887) := X"00000000";
        ram_buffer(10888) := X"24640001";
        ram_buffer(10889) := X"AC440000";
        ram_buffer(10890) := X"A0710000";
        ram_buffer(10891) := X"8C430004";
        ram_buffer(10892) := X"00000000";
        ram_buffer(10893) := X"2463FFFF";
        ram_buffer(10894) := X"106000AA";
        ram_buffer(10895) := X"AC430004";
        ram_buffer(10896) := X"8E020014";
        ram_buffer(10897) := X"8E110018";
        ram_buffer(10898) := X"8C430000";
        ram_buffer(10899) := X"00112203";
        ram_buffer(10900) := X"24650001";
        ram_buffer(10901) := X"AC450000";
        ram_buffer(10902) := X"A0640000";
        ram_buffer(10903) := X"8C430004";
        ram_buffer(10904) := X"00000000";
        ram_buffer(10905) := X"2463FFFF";
        ram_buffer(10906) := X"106000B6";
        ram_buffer(10907) := X"AC430004";
        ram_buffer(10908) := X"8E020014";
        ram_buffer(10909) := X"00000000";
        ram_buffer(10910) := X"8C430000";
        ram_buffer(10911) := X"00000000";
        ram_buffer(10912) := X"24640001";
        ram_buffer(10913) := X"AC440000";
        ram_buffer(10914) := X"A0710000";
        ram_buffer(10915) := X"8C430004";
        ram_buffer(10916) := X"00000000";
        ram_buffer(10917) := X"2463FFFF";
        ram_buffer(10918) := X"106000C2";
        ram_buffer(10919) := X"AC430004";
        ram_buffer(10920) := X"8E020014";
        ram_buffer(10921) := X"8E040034";
        ram_buffer(10922) := X"8C430000";
        ram_buffer(10923) := X"00000000";
        ram_buffer(10924) := X"24650001";
        ram_buffer(10925) := X"AC450000";
        ram_buffer(10926) := X"A0640000";
        ram_buffer(10927) := X"8C430004";
        ram_buffer(10928) := X"00000000";
        ram_buffer(10929) := X"2463FFFF";
        ram_buffer(10930) := X"106000CE";
        ram_buffer(10931) := X"AC430004";
        ram_buffer(10932) := X"8E020034";
        ram_buffer(10933) := X"8E11003C";
        ram_buffer(10934) := X"00009021";
        ram_buffer(10935) := X"1C400022";
        ram_buffer(10936) := X"24130016";
        ram_buffer(10937) := X"100000E6";
        ram_buffer(10938) := X"00000000";
        ram_buffer(10939) := X"8E030014";
        ram_buffer(10940) := X"8E220008";
        ram_buffer(10941) := X"8E25000C";
        ram_buffer(10942) := X"8C640000";
        ram_buffer(10943) := X"00021100";
        ram_buffer(10944) := X"00451021";
        ram_buffer(10945) := X"24850001";
        ram_buffer(10946) := X"AC650000";
        ram_buffer(10947) := X"A0820000";
        ram_buffer(10948) := X"8C620004";
        ram_buffer(10949) := X"00000000";
        ram_buffer(10950) := X"2442FFFF";
        ram_buffer(10951) := X"104000DF";
        ram_buffer(10952) := X"AC620004";
        ram_buffer(10953) := X"8E020014";
        ram_buffer(10954) := X"8E240010";
        ram_buffer(10955) := X"8C430000";
        ram_buffer(10956) := X"26310054";
        ram_buffer(10957) := X"24650001";
        ram_buffer(10958) := X"AC450000";
        ram_buffer(10959) := X"A0640000";
        ram_buffer(10960) := X"8C430004";
        ram_buffer(10961) := X"00000000";
        ram_buffer(10962) := X"2463FFFF";
        ram_buffer(10963) := X"106000BB";
        ram_buffer(10964) := X"AC430004";
        ram_buffer(10965) := X"8E020034";
        ram_buffer(10966) := X"00000000";
        ram_buffer(10967) := X"0242102A";
        ram_buffer(10968) := X"104000C7";
        ram_buffer(10969) := X"00000000";
        ram_buffer(10970) := X"8E020014";
        ram_buffer(10971) := X"8E240000";
        ram_buffer(10972) := X"8C430000";
        ram_buffer(10973) := X"26520001";
        ram_buffer(10974) := X"24650001";
        ram_buffer(10975) := X"AC450000";
        ram_buffer(10976) := X"A0640000";
        ram_buffer(10977) := X"8C430004";
        ram_buffer(10978) := X"00000000";
        ram_buffer(10979) := X"2463FFFF";
        ram_buffer(10980) := X"1460FFD6";
        ram_buffer(10981) := X"AC430004";
        ram_buffer(10982) := X"8C42000C";
        ram_buffer(10983) := X"00000000";
        ram_buffer(10984) := X"0040F809";
        ram_buffer(10985) := X"02002021";
        ram_buffer(10986) := X"1440FFD0";
        ram_buffer(10987) := X"02002021";
        ram_buffer(10988) := X"8E020000";
        ram_buffer(10989) := X"00000000";
        ram_buffer(10990) := X"8C430000";
        ram_buffer(10991) := X"00000000";
        ram_buffer(10992) := X"0060F809";
        ram_buffer(10993) := X"AC530014";
        ram_buffer(10994) := X"1000FFC8";
        ram_buffer(10995) := X"00000000";
        ram_buffer(10996) := X"8E020000";
        ram_buffer(10997) := X"3403FFFF";
        ram_buffer(10998) := X"AC430018";
        ram_buffer(10999) := X"8E030000";
        ram_buffer(11000) := X"24040028";
        ram_buffer(11001) := X"8C630000";
        ram_buffer(11002) := X"AC440014";
        ram_buffer(11003) := X"0060F809";
        ram_buffer(11004) := X"02002021";
        ram_buffer(11005) := X"8E020014";
        ram_buffer(11006) := X"8E040030";
        ram_buffer(11007) := X"8C430000";
        ram_buffer(11008) := X"00000000";
        ram_buffer(11009) := X"24650001";
        ram_buffer(11010) := X"AC450000";
        ram_buffer(11011) := X"A0640000";
        ram_buffer(11012) := X"8C430004";
        ram_buffer(11013) := X"00000000";
        ram_buffer(11014) := X"2463FFFF";
        ram_buffer(11015) := X"1460FF70";
        ram_buffer(11016) := X"AC430004";
        ram_buffer(11017) := X"8C42000C";
        ram_buffer(11018) := X"00000000";
        ram_buffer(11019) := X"0040F809";
        ram_buffer(11020) := X"02002021";
        ram_buffer(11021) := X"1440FF6A";
        ram_buffer(11022) := X"24040016";
        ram_buffer(11023) := X"8E020000";
        ram_buffer(11024) := X"00000000";
        ram_buffer(11025) := X"8C430000";
        ram_buffer(11026) := X"AC440014";
        ram_buffer(11027) := X"0060F809";
        ram_buffer(11028) := X"02002021";
        ram_buffer(11029) := X"8E020014";
        ram_buffer(11030) := X"8E11001C";
        ram_buffer(11031) := X"8C430000";
        ram_buffer(11032) := X"00112203";
        ram_buffer(11033) := X"24650001";
        ram_buffer(11034) := X"AC450000";
        ram_buffer(11035) := X"A0640000";
        ram_buffer(11036) := X"8C430004";
        ram_buffer(11037) := X"00000000";
        ram_buffer(11038) := X"2463FFFF";
        ram_buffer(11039) := X"1460FF64";
        ram_buffer(11040) := X"AC430004";
        ram_buffer(11041) := X"8C42000C";
        ram_buffer(11042) := X"00000000";
        ram_buffer(11043) := X"0040F809";
        ram_buffer(11044) := X"02002021";
        ram_buffer(11045) := X"1440FF5E";
        ram_buffer(11046) := X"24040016";
        ram_buffer(11047) := X"8E020000";
        ram_buffer(11048) := X"00000000";
        ram_buffer(11049) := X"8C430000";
        ram_buffer(11050) := X"AC440014";
        ram_buffer(11051) := X"0060F809";
        ram_buffer(11052) := X"02002021";
        ram_buffer(11053) := X"8E020014";
        ram_buffer(11054) := X"00000000";
        ram_buffer(11055) := X"8C430000";
        ram_buffer(11056) := X"00000000";
        ram_buffer(11057) := X"24640001";
        ram_buffer(11058) := X"AC440000";
        ram_buffer(11059) := X"A0710000";
        ram_buffer(11060) := X"8C430004";
        ram_buffer(11061) := X"00000000";
        ram_buffer(11062) := X"2463FFFF";
        ram_buffer(11063) := X"1460FF58";
        ram_buffer(11064) := X"AC430004";
        ram_buffer(11065) := X"8C42000C";
        ram_buffer(11066) := X"00000000";
        ram_buffer(11067) := X"0040F809";
        ram_buffer(11068) := X"02002021";
        ram_buffer(11069) := X"1440FF52";
        ram_buffer(11070) := X"24040016";
        ram_buffer(11071) := X"8E020000";
        ram_buffer(11072) := X"00000000";
        ram_buffer(11073) := X"8C430000";
        ram_buffer(11074) := X"AC440014";
        ram_buffer(11075) := X"0060F809";
        ram_buffer(11076) := X"02002021";
        ram_buffer(11077) := X"8E020014";
        ram_buffer(11078) := X"8E110018";
        ram_buffer(11079) := X"8C430000";
        ram_buffer(11080) := X"00112203";
        ram_buffer(11081) := X"24650001";
        ram_buffer(11082) := X"AC450000";
        ram_buffer(11083) := X"A0640000";
        ram_buffer(11084) := X"8C430004";
        ram_buffer(11085) := X"00000000";
        ram_buffer(11086) := X"2463FFFF";
        ram_buffer(11087) := X"1460FF4C";
        ram_buffer(11088) := X"AC430004";
        ram_buffer(11089) := X"8C42000C";
        ram_buffer(11090) := X"00000000";
        ram_buffer(11091) := X"0040F809";
        ram_buffer(11092) := X"02002021";
        ram_buffer(11093) := X"1440FF46";
        ram_buffer(11094) := X"24040016";
        ram_buffer(11095) := X"8E020000";
        ram_buffer(11096) := X"00000000";
        ram_buffer(11097) := X"8C430000";
        ram_buffer(11098) := X"AC440014";
        ram_buffer(11099) := X"0060F809";
        ram_buffer(11100) := X"02002021";
        ram_buffer(11101) := X"8E020014";
        ram_buffer(11102) := X"00000000";
        ram_buffer(11103) := X"8C430000";
        ram_buffer(11104) := X"00000000";
        ram_buffer(11105) := X"24640001";
        ram_buffer(11106) := X"AC440000";
        ram_buffer(11107) := X"A0710000";
        ram_buffer(11108) := X"8C430004";
        ram_buffer(11109) := X"00000000";
        ram_buffer(11110) := X"2463FFFF";
        ram_buffer(11111) := X"1460FF40";
        ram_buffer(11112) := X"AC430004";
        ram_buffer(11113) := X"8C42000C";
        ram_buffer(11114) := X"00000000";
        ram_buffer(11115) := X"0040F809";
        ram_buffer(11116) := X"02002021";
        ram_buffer(11117) := X"1440FF3A";
        ram_buffer(11118) := X"24040016";
        ram_buffer(11119) := X"8E020000";
        ram_buffer(11120) := X"00000000";
        ram_buffer(11121) := X"8C430000";
        ram_buffer(11122) := X"AC440014";
        ram_buffer(11123) := X"0060F809";
        ram_buffer(11124) := X"02002021";
        ram_buffer(11125) := X"8E020014";
        ram_buffer(11126) := X"8E040034";
        ram_buffer(11127) := X"8C430000";
        ram_buffer(11128) := X"00000000";
        ram_buffer(11129) := X"24650001";
        ram_buffer(11130) := X"AC450000";
        ram_buffer(11131) := X"A0640000";
        ram_buffer(11132) := X"8C430004";
        ram_buffer(11133) := X"00000000";
        ram_buffer(11134) := X"2463FFFF";
        ram_buffer(11135) := X"1460FF34";
        ram_buffer(11136) := X"AC430004";
        ram_buffer(11137) := X"8C42000C";
        ram_buffer(11138) := X"00000000";
        ram_buffer(11139) := X"0040F809";
        ram_buffer(11140) := X"02002021";
        ram_buffer(11141) := X"1440FF2E";
        ram_buffer(11142) := X"24040016";
        ram_buffer(11143) := X"8E020000";
        ram_buffer(11144) := X"00000000";
        ram_buffer(11145) := X"8C430000";
        ram_buffer(11146) := X"AC440014";
        ram_buffer(11147) := X"0060F809";
        ram_buffer(11148) := X"02002021";
        ram_buffer(11149) := X"1000FF26";
        ram_buffer(11150) := X"00000000";
        ram_buffer(11151) := X"8C42000C";
        ram_buffer(11152) := X"00000000";
        ram_buffer(11153) := X"0040F809";
        ram_buffer(11154) := X"02002021";
        ram_buffer(11155) := X"1440FF41";
        ram_buffer(11156) := X"02002021";
        ram_buffer(11157) := X"8E020000";
        ram_buffer(11158) := X"00000000";
        ram_buffer(11159) := X"8C430000";
        ram_buffer(11160) := X"00000000";
        ram_buffer(11161) := X"0060F809";
        ram_buffer(11162) := X"AC530014";
        ram_buffer(11163) := X"8E020034";
        ram_buffer(11164) := X"00000000";
        ram_buffer(11165) := X"0242102A";
        ram_buffer(11166) := X"1440FF3B";
        ram_buffer(11167) := X"00000000";
        ram_buffer(11168) := X"8FBF0024";
        ram_buffer(11169) := X"8FB30020";
        ram_buffer(11170) := X"8FB2001C";
        ram_buffer(11171) := X"8FB10018";
        ram_buffer(11172) := X"8FB00014";
        ram_buffer(11173) := X"03E00008";
        ram_buffer(11174) := X"27BD0028";
        ram_buffer(11175) := X"8C62000C";
        ram_buffer(11176) := X"00000000";
        ram_buffer(11177) := X"0040F809";
        ram_buffer(11178) := X"02002021";
        ram_buffer(11179) := X"1440FF1D";
        ram_buffer(11180) := X"02002021";
        ram_buffer(11181) := X"8E020000";
        ram_buffer(11182) := X"00000000";
        ram_buffer(11183) := X"8C430000";
        ram_buffer(11184) := X"00000000";
        ram_buffer(11185) := X"0060F809";
        ram_buffer(11186) := X"AC530014";
        ram_buffer(11187) := X"1000FF15";
        ram_buffer(11188) := X"00000000";
        ram_buffer(11189) := X"8C42000C";
        ram_buffer(11190) := X"00000000";
        ram_buffer(11191) := X"0040F809";
        ram_buffer(11192) := X"00000000";
        ram_buffer(11193) := X"1440FE81";
        ram_buffer(11194) := X"24040016";
        ram_buffer(11195) := X"8E020000";
        ram_buffer(11196) := X"00000000";
        ram_buffer(11197) := X"8C430000";
        ram_buffer(11198) := X"AC440014";
        ram_buffer(11199) := X"0060F809";
        ram_buffer(11200) := X"02002021";
        ram_buffer(11201) := X"8E020014";
        ram_buffer(11202) := X"00000000";
        ram_buffer(11203) := X"8C430000";
        ram_buffer(11204) := X"00000000";
        ram_buffer(11205) := X"24640001";
        ram_buffer(11206) := X"AC440000";
        ram_buffer(11207) := X"A0710000";
        ram_buffer(11208) := X"8C430004";
        ram_buffer(11209) := X"00000000";
        ram_buffer(11210) := X"2463FFFF";
        ram_buffer(11211) := X"1460FE7B";
        ram_buffer(11212) := X"AC430004";
        ram_buffer(11213) := X"8C42000C";
        ram_buffer(11214) := X"00000000";
        ram_buffer(11215) := X"0040F809";
        ram_buffer(11216) := X"02002021";
        ram_buffer(11217) := X"1440FE75";
        ram_buffer(11218) := X"24040016";
        ram_buffer(11219) := X"8E020000";
        ram_buffer(11220) := X"00000000";
        ram_buffer(11221) := X"8C430000";
        ram_buffer(11222) := X"AC440014";
        ram_buffer(11223) := X"0060F809";
        ram_buffer(11224) := X"02002021";
        ram_buffer(11225) := X"1000FE6D";
        ram_buffer(11226) := X"00000000";
        ram_buffer(11227) := X"8C42000C";
        ram_buffer(11228) := X"00000000";
        ram_buffer(11229) := X"0040F809";
        ram_buffer(11230) := X"02002021";
        ram_buffer(11231) := X"1440FE82";
        ram_buffer(11232) := X"24040016";
        ram_buffer(11233) := X"8E020000";
        ram_buffer(11234) := X"00000000";
        ram_buffer(11235) := X"8C430000";
        ram_buffer(11236) := X"AC440014";
        ram_buffer(11237) := X"0060F809";
        ram_buffer(11238) := X"02002021";
        ram_buffer(11239) := X"1000FE7A";
        ram_buffer(11240) := X"00000000";
        ram_buffer(11241) := X"8C62000C";
        ram_buffer(11242) := X"00000000";
        ram_buffer(11243) := X"0040F809";
        ram_buffer(11244) := X"02002021";
        ram_buffer(11245) := X"1440FE68";
        ram_buffer(11246) := X"24040016";
        ram_buffer(11247) := X"8E020000";
        ram_buffer(11248) := X"00000000";
        ram_buffer(11249) := X"8C430000";
        ram_buffer(11250) := X"AC440014";
        ram_buffer(11251) := X"0060F809";
        ram_buffer(11252) := X"02002021";
        ram_buffer(11253) := X"1000FE60";
        ram_buffer(11254) := X"00000000";
        ram_buffer(11255) := X"27BDFFD0";
        ram_buffer(11256) := X"AFB10018";
        ram_buffer(11257) := X"AFB00014";
        ram_buffer(11258) := X"AFBF002C";
        ram_buffer(11259) := X"AFB50028";
        ram_buffer(11260) := X"AFB40024";
        ram_buffer(11261) := X"AFB30020";
        ram_buffer(11262) := X"AFB2001C";
        ram_buffer(11263) := X"00808821";
        ram_buffer(11264) := X"10C00015";
        ram_buffer(11265) := X"00A08021";
        ram_buffer(11266) := X"24A20018";
        ram_buffer(11267) := X"00021080";
        ram_buffer(11268) := X"00821021";
        ram_buffer(11269) := X"8C530000";
        ram_buffer(11270) := X"24B00010";
        ram_buffer(11271) := X"126000FD";
        ram_buffer(11272) := X"24040031";
        ram_buffer(11273) := X"8E620114";
        ram_buffer(11274) := X"00000000";
        ram_buffer(11275) := X"10400010";
        ram_buffer(11276) := X"00000000";
        ram_buffer(11277) := X"8FBF002C";
        ram_buffer(11278) := X"8FB50028";
        ram_buffer(11279) := X"8FB40024";
        ram_buffer(11280) := X"8FB30020";
        ram_buffer(11281) := X"8FB2001C";
        ram_buffer(11282) := X"8FB10018";
        ram_buffer(11283) := X"8FB00014";
        ram_buffer(11284) := X"03E00008";
        ram_buffer(11285) := X"27BD0030";
        ram_buffer(11286) := X"24A20014";
        ram_buffer(11287) := X"00021080";
        ram_buffer(11288) := X"00821021";
        ram_buffer(11289) := X"8C530000";
        ram_buffer(11290) := X"1000FFEC";
        ram_buffer(11291) := X"00000000";
        ram_buffer(11292) := X"8E220014";
        ram_buffer(11293) := X"00000000";
        ram_buffer(11294) := X"8C430000";
        ram_buffer(11295) := X"00000000";
        ram_buffer(11296) := X"24640001";
        ram_buffer(11297) := X"AC440000";
        ram_buffer(11298) := X"2404FFFF";
        ram_buffer(11299) := X"A0640000";
        ram_buffer(11300) := X"8C430004";
        ram_buffer(11301) := X"00000000";
        ram_buffer(11302) := X"2463FFFF";
        ram_buffer(11303) := X"10600097";
        ram_buffer(11304) := X"AC430004";
        ram_buffer(11305) := X"8E220014";
        ram_buffer(11306) := X"00000000";
        ram_buffer(11307) := X"8C430000";
        ram_buffer(11308) := X"00000000";
        ram_buffer(11309) := X"24640001";
        ram_buffer(11310) := X"AC440000";
        ram_buffer(11311) := X"2404FFC4";
        ram_buffer(11312) := X"A0640000";
        ram_buffer(11313) := X"8C430004";
        ram_buffer(11314) := X"00000000";
        ram_buffer(11315) := X"2463FFFF";
        ram_buffer(11316) := X"106000C2";
        ram_buffer(11317) := X"AC430004";
        ram_buffer(11318) := X"92640002";
        ram_buffer(11319) := X"92650001";
        ram_buffer(11320) := X"92630003";
        ram_buffer(11321) := X"92620004";
        ram_buffer(11322) := X"00852821";
        ram_buffer(11323) := X"00652821";
        ram_buffer(11324) := X"92640005";
        ram_buffer(11325) := X"92630006";
        ram_buffer(11326) := X"00452821";
        ram_buffer(11327) := X"00852821";
        ram_buffer(11328) := X"92620007";
        ram_buffer(11329) := X"92640008";
        ram_buffer(11330) := X"00652821";
        ram_buffer(11331) := X"00452821";
        ram_buffer(11332) := X"92630009";
        ram_buffer(11333) := X"9262000A";
        ram_buffer(11334) := X"00852821";
        ram_buffer(11335) := X"00652821";
        ram_buffer(11336) := X"9264000B";
        ram_buffer(11337) := X"9263000C";
        ram_buffer(11338) := X"00452821";
        ram_buffer(11339) := X"00852821";
        ram_buffer(11340) := X"9262000D";
        ram_buffer(11341) := X"9264000E";
        ram_buffer(11342) := X"00652821";
        ram_buffer(11343) := X"00452821";
        ram_buffer(11344) := X"9263000F";
        ram_buffer(11345) := X"8E220014";
        ram_buffer(11346) := X"92740010";
        ram_buffer(11347) := X"00852021";
        ram_buffer(11348) := X"00641821";
        ram_buffer(11349) := X"0283A021";
        ram_buffer(11350) := X"8C440000";
        ram_buffer(11351) := X"26920013";
        ram_buffer(11352) := X"00121A03";
        ram_buffer(11353) := X"24850001";
        ram_buffer(11354) := X"AC450000";
        ram_buffer(11355) := X"A0830000";
        ram_buffer(11356) := X"8C430004";
        ram_buffer(11357) := X"00000000";
        ram_buffer(11358) := X"2463FFFF";
        ram_buffer(11359) := X"10600089";
        ram_buffer(11360) := X"AC430004";
        ram_buffer(11361) := X"8E220014";
        ram_buffer(11362) := X"00000000";
        ram_buffer(11363) := X"8C430000";
        ram_buffer(11364) := X"00000000";
        ram_buffer(11365) := X"24640001";
        ram_buffer(11366) := X"AC440000";
        ram_buffer(11367) := X"A0720000";
        ram_buffer(11368) := X"8C430004";
        ram_buffer(11369) := X"00000000";
        ram_buffer(11370) := X"2463FFFF";
        ram_buffer(11371) := X"1060006F";
        ram_buffer(11372) := X"AC430004";
        ram_buffer(11373) := X"8E220014";
        ram_buffer(11374) := X"00000000";
        ram_buffer(11375) := X"8C430000";
        ram_buffer(11376) := X"00000000";
        ram_buffer(11377) := X"24640001";
        ram_buffer(11378) := X"AC440000";
        ram_buffer(11379) := X"A0700000";
        ram_buffer(11380) := X"8C430004";
        ram_buffer(11381) := X"00000000";
        ram_buffer(11382) := X"2463FFFF";
        ram_buffer(11383) := X"10600055";
        ram_buffer(11384) := X"AC430004";
        ram_buffer(11385) := X"26720001";
        ram_buffer(11386) := X"26700011";
        ram_buffer(11387) := X"24150016";
        ram_buffer(11388) := X"8E220014";
        ram_buffer(11389) := X"92440000";
        ram_buffer(11390) := X"8C430000";
        ram_buffer(11391) := X"26520001";
        ram_buffer(11392) := X"24650001";
        ram_buffer(11393) := X"AC450000";
        ram_buffer(11394) := X"A0640000";
        ram_buffer(11395) := X"8C430004";
        ram_buffer(11396) := X"00000000";
        ram_buffer(11397) := X"2463FFFF";
        ram_buffer(11398) := X"10600018";
        ram_buffer(11399) := X"AC430004";
        ram_buffer(11400) := X"1650FFF3";
        ram_buffer(11401) := X"00000000";
        ram_buffer(11402) := X"12800011";
        ram_buffer(11403) := X"26920011";
        ram_buffer(11404) := X"02729021";
        ram_buffer(11405) := X"24140016";
        ram_buffer(11406) := X"8E220014";
        ram_buffer(11407) := X"92040000";
        ram_buffer(11408) := X"8C430000";
        ram_buffer(11409) := X"26100001";
        ram_buffer(11410) := X"24650001";
        ram_buffer(11411) := X"AC450000";
        ram_buffer(11412) := X"A0640000";
        ram_buffer(11413) := X"8C430004";
        ram_buffer(11414) := X"00000000";
        ram_buffer(11415) := X"2463FFFF";
        ram_buffer(11416) := X"10600016";
        ram_buffer(11417) := X"AC430004";
        ram_buffer(11418) := X"1612FFF3";
        ram_buffer(11419) := X"00000000";
        ram_buffer(11420) := X"24020001";
        ram_buffer(11421) := X"1000FF6F";
        ram_buffer(11422) := X"AE620114";
        ram_buffer(11423) := X"8C42000C";
        ram_buffer(11424) := X"00000000";
        ram_buffer(11425) := X"0040F809";
        ram_buffer(11426) := X"02202021";
        ram_buffer(11427) := X"1440FFE4";
        ram_buffer(11428) := X"02202021";
        ram_buffer(11429) := X"8E220000";
        ram_buffer(11430) := X"00000000";
        ram_buffer(11431) := X"8C430000";
        ram_buffer(11432) := X"00000000";
        ram_buffer(11433) := X"0060F809";
        ram_buffer(11434) := X"AC550014";
        ram_buffer(11435) := X"1650FFD0";
        ram_buffer(11436) := X"00000000";
        ram_buffer(11437) := X"1000FFDC";
        ram_buffer(11438) := X"00000000";
        ram_buffer(11439) := X"8C42000C";
        ram_buffer(11440) := X"00000000";
        ram_buffer(11441) := X"0040F809";
        ram_buffer(11442) := X"02202021";
        ram_buffer(11443) := X"1440FFE6";
        ram_buffer(11444) := X"02202021";
        ram_buffer(11445) := X"8E220000";
        ram_buffer(11446) := X"00000000";
        ram_buffer(11447) := X"8C430000";
        ram_buffer(11448) := X"00000000";
        ram_buffer(11449) := X"0060F809";
        ram_buffer(11450) := X"AC540014";
        ram_buffer(11451) := X"1612FFD2";
        ram_buffer(11452) := X"24020001";
        ram_buffer(11453) := X"1000FF4F";
        ram_buffer(11454) := X"AE620114";
        ram_buffer(11455) := X"8C42000C";
        ram_buffer(11456) := X"00000000";
        ram_buffer(11457) := X"0040F809";
        ram_buffer(11458) := X"02202021";
        ram_buffer(11459) := X"1440FF65";
        ram_buffer(11460) := X"24040016";
        ram_buffer(11461) := X"8E220000";
        ram_buffer(11462) := X"00000000";
        ram_buffer(11463) := X"8C430000";
        ram_buffer(11464) := X"AC440014";
        ram_buffer(11465) := X"0060F809";
        ram_buffer(11466) := X"02202021";
        ram_buffer(11467) := X"1000FF5D";
        ram_buffer(11468) := X"00000000";
        ram_buffer(11469) := X"8C42000C";
        ram_buffer(11470) := X"00000000";
        ram_buffer(11471) := X"0040F809";
        ram_buffer(11472) := X"02202021";
        ram_buffer(11473) := X"1440FFA7";
        ram_buffer(11474) := X"24040016";
        ram_buffer(11475) := X"8E220000";
        ram_buffer(11476) := X"00000000";
        ram_buffer(11477) := X"8C430000";
        ram_buffer(11478) := X"AC440014";
        ram_buffer(11479) := X"0060F809";
        ram_buffer(11480) := X"02202021";
        ram_buffer(11481) := X"1000FFA0";
        ram_buffer(11482) := X"26720001";
        ram_buffer(11483) := X"8C42000C";
        ram_buffer(11484) := X"00000000";
        ram_buffer(11485) := X"0040F809";
        ram_buffer(11486) := X"02202021";
        ram_buffer(11487) := X"1440FF8D";
        ram_buffer(11488) := X"24040016";
        ram_buffer(11489) := X"8E220000";
        ram_buffer(11490) := X"00000000";
        ram_buffer(11491) := X"8C430000";
        ram_buffer(11492) := X"AC440014";
        ram_buffer(11493) := X"0060F809";
        ram_buffer(11494) := X"02202021";
        ram_buffer(11495) := X"1000FF85";
        ram_buffer(11496) := X"00000000";
        ram_buffer(11497) := X"8C42000C";
        ram_buffer(11498) := X"00000000";
        ram_buffer(11499) := X"0040F809";
        ram_buffer(11500) := X"02202021";
        ram_buffer(11501) := X"1440FF73";
        ram_buffer(11502) := X"24040016";
        ram_buffer(11503) := X"8E220000";
        ram_buffer(11504) := X"00000000";
        ram_buffer(11505) := X"8C430000";
        ram_buffer(11506) := X"AC440014";
        ram_buffer(11507) := X"0060F809";
        ram_buffer(11508) := X"02202021";
        ram_buffer(11509) := X"1000FF6B";
        ram_buffer(11510) := X"00000000";
        ram_buffer(11511) := X"8C42000C";
        ram_buffer(11512) := X"00000000";
        ram_buffer(11513) := X"0040F809";
        ram_buffer(11514) := X"02202021";
        ram_buffer(11515) := X"1440FF3A";
        ram_buffer(11516) := X"24040016";
        ram_buffer(11517) := X"8E220000";
        ram_buffer(11518) := X"00000000";
        ram_buffer(11519) := X"8C430000";
        ram_buffer(11520) := X"AC440014";
        ram_buffer(11521) := X"0060F809";
        ram_buffer(11522) := X"02202021";
        ram_buffer(11523) := X"1000FF32";
        ram_buffer(11524) := X"00000000";
        ram_buffer(11525) := X"8E220000";
        ram_buffer(11526) := X"00000000";
        ram_buffer(11527) := X"AC500018";
        ram_buffer(11528) := X"8E230000";
        ram_buffer(11529) := X"AC440014";
        ram_buffer(11530) := X"8C620000";
        ram_buffer(11531) := X"00000000";
        ram_buffer(11532) := X"0040F809";
        ram_buffer(11533) := X"02202021";
        ram_buffer(11534) := X"1000FEFA";
        ram_buffer(11535) := X"00000000";
        ram_buffer(11536) := X"8C8200AC";
        ram_buffer(11537) := X"27BDFFE0";
        ram_buffer(11538) := X"AFB00014";
        ram_buffer(11539) := X"AFBF001C";
        ram_buffer(11540) := X"AFB10018";
        ram_buffer(11541) := X"1440002A";
        ram_buffer(11542) := X"00808021";
        ram_buffer(11543) := X"8C8200EC";
        ram_buffer(11544) := X"00000000";
        ram_buffer(11545) := X"18400026";
        ram_buffer(11546) := X"00000000";
        ram_buffer(11547) := X"8C8300DC";
        ram_buffer(11548) := X"8C9100F0";
        ram_buffer(11549) := X"10600337";
        ram_buffer(11550) := X"00000000";
        ram_buffer(11551) := X"8C830134";
        ram_buffer(11552) := X"00000000";
        ram_buffer(11553) := X"1460033D";
        ram_buffer(11554) := X"00000000";
        ram_buffer(11555) := X"8C83013C";
        ram_buffer(11556) := X"00000000";
        ram_buffer(11557) := X"1060029D";
        ram_buffer(11558) := X"24030001";
        ram_buffer(11559) := X"10430018";
        ram_buffer(11560) := X"00000000";
        ram_buffer(11561) := X"8E1100F4";
        ram_buffer(11562) := X"8E03013C";
        ram_buffer(11563) := X"00000000";
        ram_buffer(11564) := X"1060033F";
        ram_buffer(11565) := X"00003021";
        ram_buffer(11566) := X"24030002";
        ram_buffer(11567) := X"10430010";
        ram_buffer(11568) := X"00000000";
        ram_buffer(11569) := X"8E1100F8";
        ram_buffer(11570) := X"8E03013C";
        ram_buffer(11571) := X"00000000";
        ram_buffer(11572) := X"10600330";
        ram_buffer(11573) := X"24030003";
        ram_buffer(11574) := X"10430009";
        ram_buffer(11575) := X"00000000";
        ram_buffer(11576) := X"8E1100FC";
        ram_buffer(11577) := X"8E02013C";
        ram_buffer(11578) := X"00000000";
        ram_buffer(11579) := X"14400004";
        ram_buffer(11580) := X"00003021";
        ram_buffer(11581) := X"8E250014";
        ram_buffer(11582) := X"0C022BF7";
        ram_buffer(11583) := X"02002021";
        ram_buffer(11584) := X"8E0200C0";
        ram_buffer(11585) := X"00000000";
        ram_buffer(11586) := X"144001B8";
        ram_buffer(11587) := X"00000000";
        ram_buffer(11588) := X"8E020014";
        ram_buffer(11589) := X"00000000";
        ram_buffer(11590) := X"8C430000";
        ram_buffer(11591) := X"00000000";
        ram_buffer(11592) := X"24640001";
        ram_buffer(11593) := X"AC440000";
        ram_buffer(11594) := X"2404FFFF";
        ram_buffer(11595) := X"A0640000";
        ram_buffer(11596) := X"8C430004";
        ram_buffer(11597) := X"00000000";
        ram_buffer(11598) := X"2463FFFF";
        ram_buffer(11599) := X"1060019D";
        ram_buffer(11600) := X"AC430004";
        ram_buffer(11601) := X"8E020014";
        ram_buffer(11602) := X"00000000";
        ram_buffer(11603) := X"8C430000";
        ram_buffer(11604) := X"00000000";
        ram_buffer(11605) := X"24640001";
        ram_buffer(11606) := X"AC440000";
        ram_buffer(11607) := X"2404FFDA";
        ram_buffer(11608) := X"A0640000";
        ram_buffer(11609) := X"8C430004";
        ram_buffer(11610) := X"00000000";
        ram_buffer(11611) := X"2463FFFF";
        ram_buffer(11612) := X"10600182";
        ram_buffer(11613) := X"AC430004";
        ram_buffer(11614) := X"8E020014";
        ram_buffer(11615) := X"8E1100EC";
        ram_buffer(11616) := X"8C430000";
        ram_buffer(11617) := X"26310003";
        ram_buffer(11618) := X"00118840";
        ram_buffer(11619) := X"24650001";
        ram_buffer(11620) := X"00112203";
        ram_buffer(11621) := X"AC450000";
        ram_buffer(11622) := X"A0640000";
        ram_buffer(11623) := X"8C430004";
        ram_buffer(11624) := X"00000000";
        ram_buffer(11625) := X"2463FFFF";
        ram_buffer(11626) := X"10600166";
        ram_buffer(11627) := X"AC430004";
        ram_buffer(11628) := X"8E020014";
        ram_buffer(11629) := X"00000000";
        ram_buffer(11630) := X"8C430000";
        ram_buffer(11631) := X"00000000";
        ram_buffer(11632) := X"24640001";
        ram_buffer(11633) := X"AC440000";
        ram_buffer(11634) := X"A0710000";
        ram_buffer(11635) := X"8C430004";
        ram_buffer(11636) := X"00000000";
        ram_buffer(11637) := X"2463FFFF";
        ram_buffer(11638) := X"10600130";
        ram_buffer(11639) := X"AC430004";
        ram_buffer(11640) := X"8E020014";
        ram_buffer(11641) := X"8E0400EC";
        ram_buffer(11642) := X"8C430000";
        ram_buffer(11643) := X"00000000";
        ram_buffer(11644) := X"24650001";
        ram_buffer(11645) := X"AC450000";
        ram_buffer(11646) := X"A0640000";
        ram_buffer(11647) := X"8C430004";
        ram_buffer(11648) := X"00000000";
        ram_buffer(11649) := X"2463FFFF";
        ram_buffer(11650) := X"10600116";
        ram_buffer(11651) := X"AC430004";
        ram_buffer(11652) := X"8E0200EC";
        ram_buffer(11653) := X"00000000";
        ram_buffer(11654) := X"18400060";
        ram_buffer(11655) := X"00000000";
        ram_buffer(11656) := X"8E020014";
        ram_buffer(11657) := X"8E1100F0";
        ram_buffer(11658) := X"8C430000";
        ram_buffer(11659) := X"8E240000";
        ram_buffer(11660) := X"24650001";
        ram_buffer(11661) := X"AC450000";
        ram_buffer(11662) := X"A0640000";
        ram_buffer(11663) := X"8C430004";
        ram_buffer(11664) := X"00000000";
        ram_buffer(11665) := X"2463FFFF";
        ram_buffer(11666) := X"106000B2";
        ram_buffer(11667) := X"AC430004";
        ram_buffer(11668) := X"8E0400DC";
        ram_buffer(11669) := X"8E230014";
        ram_buffer(11670) := X"8E220018";
        ram_buffer(11671) := X"1080007A";
        ram_buffer(11672) := X"00000000";
        ram_buffer(11673) := X"8E040134";
        ram_buffer(11674) := X"00000000";
        ram_buffer(11675) := X"14800079";
        ram_buffer(11676) := X"304200FF";
        ram_buffer(11677) := X"8E02013C";
        ram_buffer(11678) := X"00000000";
        ram_buffer(11679) := X"10400221";
        ram_buffer(11680) := X"00031100";
        ram_buffer(11681) := X"8E0200AC";
        ram_buffer(11682) := X"00000000";
        ram_buffer(11683) := X"1440021C";
        ram_buffer(11684) := X"00000000";
        ram_buffer(11685) := X"1000006F";
        ram_buffer(11686) := X"00001021";
        ram_buffer(11687) := X"00031900";
        ram_buffer(11688) := X"00621021";
        ram_buffer(11689) := X"304200FF";
        ram_buffer(11690) := X"8E030014";
        ram_buffer(11691) := X"00000000";
        ram_buffer(11692) := X"8C640000";
        ram_buffer(11693) := X"00000000";
        ram_buffer(11694) := X"24850001";
        ram_buffer(11695) := X"AC650000";
        ram_buffer(11696) := X"A0820000";
        ram_buffer(11697) := X"8C620004";
        ram_buffer(11698) := X"00000000";
        ram_buffer(11699) := X"2442FFFF";
        ram_buffer(11700) := X"104001DB";
        ram_buffer(11701) := X"AC620004";
        ram_buffer(11702) := X"8E0200EC";
        ram_buffer(11703) := X"00000000";
        ram_buffer(11704) := X"28420004";
        ram_buffer(11705) := X"1440002D";
        ram_buffer(11706) := X"00000000";
        ram_buffer(11707) := X"8E020014";
        ram_buffer(11708) := X"8E1100FC";
        ram_buffer(11709) := X"8C430000";
        ram_buffer(11710) := X"8E240000";
        ram_buffer(11711) := X"24650001";
        ram_buffer(11712) := X"AC450000";
        ram_buffer(11713) := X"A0640000";
        ram_buffer(11714) := X"8C430004";
        ram_buffer(11715) := X"00000000";
        ram_buffer(11716) := X"2463FFFF";
        ram_buffer(11717) := X"106001BC";
        ram_buffer(11718) := X"AC430004";
        ram_buffer(11719) := X"8E0400DC";
        ram_buffer(11720) := X"8E230014";
        ram_buffer(11721) := X"8E220018";
        ram_buffer(11722) := X"148000C0";
        ram_buffer(11723) := X"00000000";
        ram_buffer(11724) := X"00031900";
        ram_buffer(11725) := X"00621021";
        ram_buffer(11726) := X"304200FF";
        ram_buffer(11727) := X"8E030014";
        ram_buffer(11728) := X"00000000";
        ram_buffer(11729) := X"8C640000";
        ram_buffer(11730) := X"00000000";
        ram_buffer(11731) := X"24850001";
        ram_buffer(11732) := X"AC650000";
        ram_buffer(11733) := X"A0820000";
        ram_buffer(11734) := X"8C620004";
        ram_buffer(11735) := X"00000000";
        ram_buffer(11736) := X"2442FFFF";
        ram_buffer(11737) := X"1440000D";
        ram_buffer(11738) := X"AC620004";
        ram_buffer(11739) := X"8C62000C";
        ram_buffer(11740) := X"00000000";
        ram_buffer(11741) := X"0040F809";
        ram_buffer(11742) := X"02002021";
        ram_buffer(11743) := X"14400007";
        ram_buffer(11744) := X"24040016";
        ram_buffer(11745) := X"8E020000";
        ram_buffer(11746) := X"00000000";
        ram_buffer(11747) := X"8C430000";
        ram_buffer(11748) := X"AC440014";
        ram_buffer(11749) := X"0060F809";
        ram_buffer(11750) := X"02002021";
        ram_buffer(11751) := X"8E020014";
        ram_buffer(11752) := X"8E040134";
        ram_buffer(11753) := X"8C430000";
        ram_buffer(11754) := X"00000000";
        ram_buffer(11755) := X"24650001";
        ram_buffer(11756) := X"AC450000";
        ram_buffer(11757) := X"A0640000";
        ram_buffer(11758) := X"8C430004";
        ram_buffer(11759) := X"00000000";
        ram_buffer(11760) := X"2463FFFF";
        ram_buffer(11761) := X"106000D1";
        ram_buffer(11762) := X"AC430004";
        ram_buffer(11763) := X"8E020014";
        ram_buffer(11764) := X"8E040138";
        ram_buffer(11765) := X"8C430000";
        ram_buffer(11766) := X"00000000";
        ram_buffer(11767) := X"24650001";
        ram_buffer(11768) := X"AC450000";
        ram_buffer(11769) := X"A0640000";
        ram_buffer(11770) := X"8C430004";
        ram_buffer(11771) := X"00000000";
        ram_buffer(11772) := X"2463FFFF";
        ram_buffer(11773) := X"106000B7";
        ram_buffer(11774) := X"AC430004";
        ram_buffer(11775) := X"8E030014";
        ram_buffer(11776) := X"8E02013C";
        ram_buffer(11777) := X"8E050140";
        ram_buffer(11778) := X"8C640000";
        ram_buffer(11779) := X"00021100";
        ram_buffer(11780) := X"00451021";
        ram_buffer(11781) := X"24850001";
        ram_buffer(11782) := X"AC650000";
        ram_buffer(11783) := X"A0820000";
        ram_buffer(11784) := X"8C620004";
        ram_buffer(11785) := X"00000000";
        ram_buffer(11786) := X"2442FFFF";
        ram_buffer(11787) := X"10400148";
        ram_buffer(11788) := X"AC620004";
        ram_buffer(11789) := X"8FBF001C";
        ram_buffer(11790) := X"8FB10018";
        ram_buffer(11791) := X"8FB00014";
        ram_buffer(11792) := X"03E00008";
        ram_buffer(11793) := X"27BD0020";
        ram_buffer(11794) := X"00031900";
        ram_buffer(11795) := X"00621021";
        ram_buffer(11796) := X"304200FF";
        ram_buffer(11797) := X"8E030014";
        ram_buffer(11798) := X"00000000";
        ram_buffer(11799) := X"8C640000";
        ram_buffer(11800) := X"00000000";
        ram_buffer(11801) := X"24850001";
        ram_buffer(11802) := X"AC650000";
        ram_buffer(11803) := X"A0820000";
        ram_buffer(11804) := X"8C620004";
        ram_buffer(11805) := X"00000000";
        ram_buffer(11806) := X"2442FFFF";
        ram_buffer(11807) := X"10400154";
        ram_buffer(11808) := X"AC620004";
        ram_buffer(11809) := X"8E0200EC";
        ram_buffer(11810) := X"00000000";
        ram_buffer(11811) := X"28420002";
        ram_buffer(11812) := X"1440FFC2";
        ram_buffer(11813) := X"00000000";
        ram_buffer(11814) := X"8E020014";
        ram_buffer(11815) := X"8E1100F4";
        ram_buffer(11816) := X"8C430000";
        ram_buffer(11817) := X"8E240000";
        ram_buffer(11818) := X"24650001";
        ram_buffer(11819) := X"AC450000";
        ram_buffer(11820) := X"A0640000";
        ram_buffer(11821) := X"8C430004";
        ram_buffer(11822) := X"00000000";
        ram_buffer(11823) := X"2463FFFF";
        ram_buffer(11824) := X"10600135";
        ram_buffer(11825) := X"AC430004";
        ram_buffer(11826) := X"8E0400DC";
        ram_buffer(11827) := X"8E230014";
        ram_buffer(11828) := X"8E220018";
        ram_buffer(11829) := X"10800022";
        ram_buffer(11830) := X"00000000";
        ram_buffer(11831) := X"8E040134";
        ram_buffer(11832) := X"00000000";
        ram_buffer(11833) := X"14800021";
        ram_buffer(11834) := X"304200FF";
        ram_buffer(11835) := X"8E02013C";
        ram_buffer(11836) := X"00000000";
        ram_buffer(11837) := X"1040017D";
        ram_buffer(11838) := X"00031100";
        ram_buffer(11839) := X"8E0200AC";
        ram_buffer(11840) := X"00000000";
        ram_buffer(11841) := X"14400178";
        ram_buffer(11842) := X"00000000";
        ram_buffer(11843) := X"10000017";
        ram_buffer(11844) := X"00001021";
        ram_buffer(11845) := X"8C42000C";
        ram_buffer(11846) := X"00000000";
        ram_buffer(11847) := X"0040F809";
        ram_buffer(11848) := X"02002021";
        ram_buffer(11849) := X"1440FF4A";
        ram_buffer(11850) := X"24040016";
        ram_buffer(11851) := X"8E020000";
        ram_buffer(11852) := X"00000000";
        ram_buffer(11853) := X"8C430000";
        ram_buffer(11854) := X"AC440014";
        ram_buffer(11855) := X"0060F809";
        ram_buffer(11856) := X"02002021";
        ram_buffer(11857) := X"8E0400DC";
        ram_buffer(11858) := X"8E230014";
        ram_buffer(11859) := X"8E220018";
        ram_buffer(11860) := X"1080FFBD";
        ram_buffer(11861) := X"00000000";
        ram_buffer(11862) := X"1000FF42";
        ram_buffer(11863) := X"00000000";
        ram_buffer(11864) := X"00031900";
        ram_buffer(11865) := X"00621021";
        ram_buffer(11866) := X"304200FF";
        ram_buffer(11867) := X"8E030014";
        ram_buffer(11868) := X"00000000";
        ram_buffer(11869) := X"8C640000";
        ram_buffer(11870) := X"00000000";
        ram_buffer(11871) := X"24850001";
        ram_buffer(11872) := X"AC650000";
        ram_buffer(11873) := X"A0820000";
        ram_buffer(11874) := X"8C620004";
        ram_buffer(11875) := X"00000000";
        ram_buffer(11876) := X"2442FFFF";
        ram_buffer(11877) := X"10400146";
        ram_buffer(11878) := X"AC620004";
        ram_buffer(11879) := X"8E0200EC";
        ram_buffer(11880) := X"00000000";
        ram_buffer(11881) := X"28420003";
        ram_buffer(11882) := X"1440FF7C";
        ram_buffer(11883) := X"00000000";
        ram_buffer(11884) := X"8E020014";
        ram_buffer(11885) := X"8E1100F8";
        ram_buffer(11886) := X"8C430000";
        ram_buffer(11887) := X"8E240000";
        ram_buffer(11888) := X"24650001";
        ram_buffer(11889) := X"AC450000";
        ram_buffer(11890) := X"A0640000";
        ram_buffer(11891) := X"8C430004";
        ram_buffer(11892) := X"00000000";
        ram_buffer(11893) := X"2463FFFF";
        ram_buffer(11894) := X"10600127";
        ram_buffer(11895) := X"AC430004";
        ram_buffer(11896) := X"8E0400DC";
        ram_buffer(11897) := X"8E230014";
        ram_buffer(11898) := X"8E220018";
        ram_buffer(11899) := X"1080FF2B";
        ram_buffer(11900) := X"00000000";
        ram_buffer(11901) := X"8E040134";
        ram_buffer(11902) := X"00000000";
        ram_buffer(11903) := X"1480FF2A";
        ram_buffer(11904) := X"304200FF";
        ram_buffer(11905) := X"8E02013C";
        ram_buffer(11906) := X"00000000";
        ram_buffer(11907) := X"1040013A";
        ram_buffer(11908) := X"00031100";
        ram_buffer(11909) := X"8E0200AC";
        ram_buffer(11910) := X"00000000";
        ram_buffer(11911) := X"14400135";
        ram_buffer(11912) := X"00000000";
        ram_buffer(11913) := X"1000FF20";
        ram_buffer(11914) := X"00001021";
        ram_buffer(11915) := X"8E040134";
        ram_buffer(11916) := X"00000000";
        ram_buffer(11917) := X"1480FF41";
        ram_buffer(11918) := X"304200FF";
        ram_buffer(11919) := X"8E02013C";
        ram_buffer(11920) := X"00000000";
        ram_buffer(11921) := X"104000D2";
        ram_buffer(11922) := X"00031100";
        ram_buffer(11923) := X"8E0200AC";
        ram_buffer(11924) := X"00000000";
        ram_buffer(11925) := X"144000CD";
        ram_buffer(11926) := X"00000000";
        ram_buffer(11927) := X"1000FF37";
        ram_buffer(11928) := X"00001021";
        ram_buffer(11929) := X"8C42000C";
        ram_buffer(11930) := X"00000000";
        ram_buffer(11931) := X"0040F809";
        ram_buffer(11932) := X"02002021";
        ram_buffer(11933) := X"1440FEE6";
        ram_buffer(11934) := X"24040016";
        ram_buffer(11935) := X"8E020000";
        ram_buffer(11936) := X"00000000";
        ram_buffer(11937) := X"8C430000";
        ram_buffer(11938) := X"AC440014";
        ram_buffer(11939) := X"0060F809";
        ram_buffer(11940) := X"02002021";
        ram_buffer(11941) := X"1000FEDE";
        ram_buffer(11942) := X"00000000";
        ram_buffer(11943) := X"8C42000C";
        ram_buffer(11944) := X"00000000";
        ram_buffer(11945) := X"0040F809";
        ram_buffer(11946) := X"02002021";
        ram_buffer(11947) := X"1440FECC";
        ram_buffer(11948) := X"24040016";
        ram_buffer(11949) := X"8E020000";
        ram_buffer(11950) := X"00000000";
        ram_buffer(11951) := X"8C430000";
        ram_buffer(11952) := X"AC440014";
        ram_buffer(11953) := X"0060F809";
        ram_buffer(11954) := X"02002021";
        ram_buffer(11955) := X"1000FEC4";
        ram_buffer(11956) := X"00000000";
        ram_buffer(11957) := X"8C42000C";
        ram_buffer(11958) := X"00000000";
        ram_buffer(11959) := X"0040F809";
        ram_buffer(11960) := X"02002021";
        ram_buffer(11961) := X"1440FF45";
        ram_buffer(11962) := X"24040016";
        ram_buffer(11963) := X"8E020000";
        ram_buffer(11964) := X"00000000";
        ram_buffer(11965) := X"8C430000";
        ram_buffer(11966) := X"AC440014";
        ram_buffer(11967) := X"0060F809";
        ram_buffer(11968) := X"02002021";
        ram_buffer(11969) := X"1000FF3D";
        ram_buffer(11970) := X"00000000";
        ram_buffer(11971) := X"8C42000C";
        ram_buffer(11972) := X"00000000";
        ram_buffer(11973) := X"0040F809";
        ram_buffer(11974) := X"02002021";
        ram_buffer(11975) := X"1440FF2B";
        ram_buffer(11976) := X"24040016";
        ram_buffer(11977) := X"8E020000";
        ram_buffer(11978) := X"00000000";
        ram_buffer(11979) := X"8C430000";
        ram_buffer(11980) := X"AC440014";
        ram_buffer(11981) := X"0060F809";
        ram_buffer(11982) := X"02002021";
        ram_buffer(11983) := X"1000FF23";
        ram_buffer(11984) := X"00000000";
        ram_buffer(11985) := X"8C42000C";
        ram_buffer(11986) := X"00000000";
        ram_buffer(11987) := X"0040F809";
        ram_buffer(11988) := X"02002021";
        ram_buffer(11989) := X"1440FE96";
        ram_buffer(11990) := X"24040016";
        ram_buffer(11991) := X"8E020000";
        ram_buffer(11992) := X"00000000";
        ram_buffer(11993) := X"8C430000";
        ram_buffer(11994) := X"AC440014";
        ram_buffer(11995) := X"0060F809";
        ram_buffer(11996) := X"02002021";
        ram_buffer(11997) := X"1000FE8E";
        ram_buffer(11998) := X"00000000";
        ram_buffer(11999) := X"8C42000C";
        ram_buffer(12000) := X"00000000";
        ram_buffer(12001) := X"0040F809";
        ram_buffer(12002) := X"02002021";
        ram_buffer(12003) := X"1440FE7A";
        ram_buffer(12004) := X"24040016";
        ram_buffer(12005) := X"8E020000";
        ram_buffer(12006) := X"00000000";
        ram_buffer(12007) := X"8C430000";
        ram_buffer(12008) := X"AC440014";
        ram_buffer(12009) := X"0060F809";
        ram_buffer(12010) := X"02002021";
        ram_buffer(12011) := X"1000FE72";
        ram_buffer(12012) := X"00000000";
        ram_buffer(12013) := X"8C42000C";
        ram_buffer(12014) := X"00000000";
        ram_buffer(12015) := X"0040F809";
        ram_buffer(12016) := X"02002021";
        ram_buffer(12017) := X"1440FE5F";
        ram_buffer(12018) := X"24040016";
        ram_buffer(12019) := X"8E020000";
        ram_buffer(12020) := X"00000000";
        ram_buffer(12021) := X"8C430000";
        ram_buffer(12022) := X"AC440014";
        ram_buffer(12023) := X"0060F809";
        ram_buffer(12024) := X"02002021";
        ram_buffer(12025) := X"1000FE57";
        ram_buffer(12026) := X"00000000";
        ram_buffer(12027) := X"8E020014";
        ram_buffer(12028) := X"00000000";
        ram_buffer(12029) := X"8C430000";
        ram_buffer(12030) := X"00000000";
        ram_buffer(12031) := X"24640001";
        ram_buffer(12032) := X"AC440000";
        ram_buffer(12033) := X"2404FFFF";
        ram_buffer(12034) := X"A0640000";
        ram_buffer(12035) := X"8C430004";
        ram_buffer(12036) := X"00000000";
        ram_buffer(12037) := X"2463FFFF";
        ram_buffer(12038) := X"106000F3";
        ram_buffer(12039) := X"AC430004";
        ram_buffer(12040) := X"8E020014";
        ram_buffer(12041) := X"00000000";
        ram_buffer(12042) := X"8C430000";
        ram_buffer(12043) := X"00000000";
        ram_buffer(12044) := X"24640001";
        ram_buffer(12045) := X"AC440000";
        ram_buffer(12046) := X"2404FFDD";
        ram_buffer(12047) := X"A0640000";
        ram_buffer(12048) := X"8C430004";
        ram_buffer(12049) := X"00000000";
        ram_buffer(12050) := X"2463FFFF";
        ram_buffer(12051) := X"1060011E";
        ram_buffer(12052) := X"AC430004";
        ram_buffer(12053) := X"8E020014";
        ram_buffer(12054) := X"00000000";
        ram_buffer(12055) := X"8C430000";
        ram_buffer(12056) := X"00000000";
        ram_buffer(12057) := X"24640001";
        ram_buffer(12058) := X"AC440000";
        ram_buffer(12059) := X"A0600000";
        ram_buffer(12060) := X"8C430004";
        ram_buffer(12061) := X"00000000";
        ram_buffer(12062) := X"2463FFFF";
        ram_buffer(12063) := X"10600104";
        ram_buffer(12064) := X"AC430004";
        ram_buffer(12065) := X"8E020014";
        ram_buffer(12066) := X"00000000";
        ram_buffer(12067) := X"8C430000";
        ram_buffer(12068) := X"00000000";
        ram_buffer(12069) := X"24640001";
        ram_buffer(12070) := X"AC440000";
        ram_buffer(12071) := X"24040004";
        ram_buffer(12072) := X"A0640000";
        ram_buffer(12073) := X"8C430004";
        ram_buffer(12074) := X"00000000";
        ram_buffer(12075) := X"2463FFFF";
        ram_buffer(12076) := X"106000E9";
        ram_buffer(12077) := X"AC430004";
        ram_buffer(12078) := X"8E020014";
        ram_buffer(12079) := X"8E1100C0";
        ram_buffer(12080) := X"8C430000";
        ram_buffer(12081) := X"00112203";
        ram_buffer(12082) := X"24650001";
        ram_buffer(12083) := X"AC450000";
        ram_buffer(12084) := X"A0640000";
        ram_buffer(12085) := X"8C430004";
        ram_buffer(12086) := X"00000000";
        ram_buffer(12087) := X"2463FFFF";
        ram_buffer(12088) := X"106000CF";
        ram_buffer(12089) := X"AC430004";
        ram_buffer(12090) := X"8E020014";
        ram_buffer(12091) := X"00000000";
        ram_buffer(12092) := X"8C430000";
        ram_buffer(12093) := X"00000000";
        ram_buffer(12094) := X"24640001";
        ram_buffer(12095) := X"AC440000";
        ram_buffer(12096) := X"A0710000";
        ram_buffer(12097) := X"8C430004";
        ram_buffer(12098) := X"00000000";
        ram_buffer(12099) := X"2463FFFF";
        ram_buffer(12100) := X"1460FDFF";
        ram_buffer(12101) := X"AC430004";
        ram_buffer(12102) := X"8C42000C";
        ram_buffer(12103) := X"00000000";
        ram_buffer(12104) := X"0040F809";
        ram_buffer(12105) := X"02002021";
        ram_buffer(12106) := X"1440FDF9";
        ram_buffer(12107) := X"24040016";
        ram_buffer(12108) := X"8E020000";
        ram_buffer(12109) := X"00000000";
        ram_buffer(12110) := X"8C430000";
        ram_buffer(12111) := X"AC440014";
        ram_buffer(12112) := X"0060F809";
        ram_buffer(12113) := X"02002021";
        ram_buffer(12114) := X"1000FDF1";
        ram_buffer(12115) := X"00000000";
        ram_buffer(12116) := X"8C62000C";
        ram_buffer(12117) := X"00000000";
        ram_buffer(12118) := X"0040F809";
        ram_buffer(12119) := X"02002021";
        ram_buffer(12120) := X"1440FEB4";
        ram_buffer(12121) := X"02002021";
        ram_buffer(12122) := X"8E020000";
        ram_buffer(12123) := X"8FBF001C";
        ram_buffer(12124) := X"8FB10018";
        ram_buffer(12125) := X"8C590000";
        ram_buffer(12126) := X"24030016";
        ram_buffer(12127) := X"8FB00014";
        ram_buffer(12128) := X"AC430014";
        ram_buffer(12129) := X"03200008";
        ram_buffer(12130) := X"27BD0020";
        ram_buffer(12131) := X"00031100";
        ram_buffer(12132) := X"1000FE6A";
        ram_buffer(12133) := X"304200FF";
        ram_buffer(12134) := X"8C42000C";
        ram_buffer(12135) := X"00000000";
        ram_buffer(12136) := X"0040F809";
        ram_buffer(12137) := X"02002021";
        ram_buffer(12138) := X"1440FEC7";
        ram_buffer(12139) := X"24040016";
        ram_buffer(12140) := X"8E020000";
        ram_buffer(12141) := X"00000000";
        ram_buffer(12142) := X"8C430000";
        ram_buffer(12143) := X"AC440014";
        ram_buffer(12144) := X"0060F809";
        ram_buffer(12145) := X"02002021";
        ram_buffer(12146) := X"1000FEBF";
        ram_buffer(12147) := X"00000000";
        ram_buffer(12148) := X"8C62000C";
        ram_buffer(12149) := X"00000000";
        ram_buffer(12150) := X"0040F809";
        ram_buffer(12151) := X"02002021";
        ram_buffer(12152) := X"1440FEA8";
        ram_buffer(12153) := X"24040016";
        ram_buffer(12154) := X"8E020000";
        ram_buffer(12155) := X"00000000";
        ram_buffer(12156) := X"8C430000";
        ram_buffer(12157) := X"AC440014";
        ram_buffer(12158) := X"0060F809";
        ram_buffer(12159) := X"02002021";
        ram_buffer(12160) := X"1000FEA0";
        ram_buffer(12161) := X"00000000";
        ram_buffer(12162) := X"8C42000C";
        ram_buffer(12163) := X"00000000";
        ram_buffer(12164) := X"0040F809";
        ram_buffer(12165) := X"02002021";
        ram_buffer(12166) := X"1440FE40";
        ram_buffer(12167) := X"24040016";
        ram_buffer(12168) := X"8E020000";
        ram_buffer(12169) := X"00000000";
        ram_buffer(12170) := X"8C430000";
        ram_buffer(12171) := X"AC440014";
        ram_buffer(12172) := X"0060F809";
        ram_buffer(12173) := X"02002021";
        ram_buffer(12174) := X"1000FE38";
        ram_buffer(12175) := X"00000000";
        ram_buffer(12176) := X"8C62000C";
        ram_buffer(12177) := X"00000000";
        ram_buffer(12178) := X"0040F809";
        ram_buffer(12179) := X"02002021";
        ram_buffer(12180) := X"1440FE21";
        ram_buffer(12181) := X"24040016";
        ram_buffer(12182) := X"8E020000";
        ram_buffer(12183) := X"00000000";
        ram_buffer(12184) := X"8C430000";
        ram_buffer(12185) := X"AC440014";
        ram_buffer(12186) := X"0060F809";
        ram_buffer(12187) := X"02002021";
        ram_buffer(12188) := X"1000FE19";
        ram_buffer(12189) := X"00000000";
        ram_buffer(12190) := X"8C42000C";
        ram_buffer(12191) := X"00000000";
        ram_buffer(12192) := X"0040F809";
        ram_buffer(12193) := X"02002021";
        ram_buffer(12194) := X"1440FED5";
        ram_buffer(12195) := X"24040016";
        ram_buffer(12196) := X"8E020000";
        ram_buffer(12197) := X"00000000";
        ram_buffer(12198) := X"8C430000";
        ram_buffer(12199) := X"AC440014";
        ram_buffer(12200) := X"0060F809";
        ram_buffer(12201) := X"02002021";
        ram_buffer(12202) := X"1000FECD";
        ram_buffer(12203) := X"00000000";
        ram_buffer(12204) := X"8C62000C";
        ram_buffer(12205) := X"00000000";
        ram_buffer(12206) := X"0040F809";
        ram_buffer(12207) := X"02002021";
        ram_buffer(12208) := X"1440FEB6";
        ram_buffer(12209) := X"24040016";
        ram_buffer(12210) := X"8E020000";
        ram_buffer(12211) := X"00000000";
        ram_buffer(12212) := X"8C430000";
        ram_buffer(12213) := X"AC440014";
        ram_buffer(12214) := X"0060F809";
        ram_buffer(12215) := X"02002021";
        ram_buffer(12216) := X"1000FEAE";
        ram_buffer(12217) := X"00000000";
        ram_buffer(12218) := X"00031100";
        ram_buffer(12219) := X"1000FE9F";
        ram_buffer(12220) := X"304200FF";
        ram_buffer(12221) := X"00031100";
        ram_buffer(12222) := X"1000FDEB";
        ram_buffer(12223) := X"304200FF";
        ram_buffer(12224) := X"00031100";
        ram_buffer(12225) := X"1000FE53";
        ram_buffer(12226) := X"304200FF";
        ram_buffer(12227) := X"8E250014";
        ram_buffer(12228) := X"0C022BF7";
        ram_buffer(12229) := X"00003021";
        ram_buffer(12230) := X"8E0200EC";
        ram_buffer(12231) := X"00000000";
        ram_buffer(12232) := X"28430002";
        ram_buffer(12233) := X"1460FD76";
        ram_buffer(12234) := X"00000000";
        ram_buffer(12235) := X"8E0300DC";
        ram_buffer(12236) := X"8E1100F4";
        ram_buffer(12237) := X"10600072";
        ram_buffer(12238) := X"02002021";
        ram_buffer(12239) := X"8E030134";
        ram_buffer(12240) := X"00000000";
        ram_buffer(12241) := X"1060FD58";
        ram_buffer(12242) := X"00000000";
        ram_buffer(12243) := X"8E250018";
        ram_buffer(12244) := X"24060001";
        ram_buffer(12245) := X"0C022BF7";
        ram_buffer(12246) := X"02002021";
        ram_buffer(12247) := X"8E0200EC";
        ram_buffer(12248) := X"00000000";
        ram_buffer(12249) := X"28430003";
        ram_buffer(12250) := X"1460FD65";
        ram_buffer(12251) := X"00000000";
        ram_buffer(12252) := X"8E0300DC";
        ram_buffer(12253) := X"8E1100F8";
        ram_buffer(12254) := X"10600070";
        ram_buffer(12255) := X"00000000";
        ram_buffer(12256) := X"8E030134";
        ram_buffer(12257) := X"00000000";
        ram_buffer(12258) := X"1060FD4F";
        ram_buffer(12259) := X"00000000";
        ram_buffer(12260) := X"8E250018";
        ram_buffer(12261) := X"24060001";
        ram_buffer(12262) := X"0C022BF7";
        ram_buffer(12263) := X"02002021";
        ram_buffer(12264) := X"8E0200EC";
        ram_buffer(12265) := X"00000000";
        ram_buffer(12266) := X"28420004";
        ram_buffer(12267) := X"1440FD54";
        ram_buffer(12268) := X"00000000";
        ram_buffer(12269) := X"8E0200DC";
        ram_buffer(12270) := X"8E1100FC";
        ram_buffer(12271) := X"10400055";
        ram_buffer(12272) := X"00000000";
        ram_buffer(12273) := X"8E030134";
        ram_buffer(12274) := X"00000000";
        ram_buffer(12275) := X"1060FD45";
        ram_buffer(12276) := X"24060001";
        ram_buffer(12277) := X"8E250018";
        ram_buffer(12278) := X"0C022BF7";
        ram_buffer(12279) := X"02002021";
        ram_buffer(12280) := X"1000FD47";
        ram_buffer(12281) := X"00000000";
        ram_buffer(12282) := X"8C42000C";
        ram_buffer(12283) := X"00000000";
        ram_buffer(12284) := X"0040F809";
        ram_buffer(12285) := X"02002021";
        ram_buffer(12286) := X"1440FF09";
        ram_buffer(12287) := X"24040016";
        ram_buffer(12288) := X"8E020000";
        ram_buffer(12289) := X"00000000";
        ram_buffer(12290) := X"8C430000";
        ram_buffer(12291) := X"AC440014";
        ram_buffer(12292) := X"0060F809";
        ram_buffer(12293) := X"02002021";
        ram_buffer(12294) := X"1000FF01";
        ram_buffer(12295) := X"00000000";
        ram_buffer(12296) := X"8C42000C";
        ram_buffer(12297) := X"00000000";
        ram_buffer(12298) := X"0040F809";
        ram_buffer(12299) := X"02002021";
        ram_buffer(12300) := X"1440FF2D";
        ram_buffer(12301) := X"24040016";
        ram_buffer(12302) := X"8E020000";
        ram_buffer(12303) := X"00000000";
        ram_buffer(12304) := X"8C430000";
        ram_buffer(12305) := X"AC440014";
        ram_buffer(12306) := X"0060F809";
        ram_buffer(12307) := X"02002021";
        ram_buffer(12308) := X"1000FF25";
        ram_buffer(12309) := X"00000000";
        ram_buffer(12310) := X"8C42000C";
        ram_buffer(12311) := X"00000000";
        ram_buffer(12312) := X"0040F809";
        ram_buffer(12313) := X"02002021";
        ram_buffer(12314) := X"1440FF13";
        ram_buffer(12315) := X"24040016";
        ram_buffer(12316) := X"8E020000";
        ram_buffer(12317) := X"00000000";
        ram_buffer(12318) := X"8C430000";
        ram_buffer(12319) := X"AC440014";
        ram_buffer(12320) := X"0060F809";
        ram_buffer(12321) := X"02002021";
        ram_buffer(12322) := X"1000FF0B";
        ram_buffer(12323) := X"00000000";
        ram_buffer(12324) := X"8C42000C";
        ram_buffer(12325) := X"00000000";
        ram_buffer(12326) := X"0040F809";
        ram_buffer(12327) := X"02002021";
        ram_buffer(12328) := X"1440FEF8";
        ram_buffer(12329) := X"24040016";
        ram_buffer(12330) := X"8E020000";
        ram_buffer(12331) := X"00000000";
        ram_buffer(12332) := X"8C430000";
        ram_buffer(12333) := X"AC440014";
        ram_buffer(12334) := X"0060F809";
        ram_buffer(12335) := X"02002021";
        ram_buffer(12336) := X"1000FEF0";
        ram_buffer(12337) := X"00000000";
        ram_buffer(12338) := X"8C42000C";
        ram_buffer(12339) := X"00000000";
        ram_buffer(12340) := X"0040F809";
        ram_buffer(12341) := X"02002021";
        ram_buffer(12342) := X"1440FEDE";
        ram_buffer(12343) := X"24040016";
        ram_buffer(12344) := X"8E020000";
        ram_buffer(12345) := X"00000000";
        ram_buffer(12346) := X"8C430000";
        ram_buffer(12347) := X"AC440014";
        ram_buffer(12348) := X"0060F809";
        ram_buffer(12349) := X"02002021";
        ram_buffer(12350) := X"1000FED6";
        ram_buffer(12351) := X"00000000";
        ram_buffer(12352) := X"8E250014";
        ram_buffer(12353) := X"0C022BF7";
        ram_buffer(12354) := X"00003021";
        ram_buffer(12355) := X"1000FF8F";
        ram_buffer(12356) := X"00000000";
        ram_buffer(12357) := X"8E250014";
        ram_buffer(12358) := X"02002021";
        ram_buffer(12359) := X"0C022BF7";
        ram_buffer(12360) := X"00003021";
        ram_buffer(12361) := X"8E250018";
        ram_buffer(12362) := X"24060001";
        ram_buffer(12363) := X"0C022BF7";
        ram_buffer(12364) := X"02002021";
        ram_buffer(12365) := X"1000FCF2";
        ram_buffer(12366) := X"00000000";
        ram_buffer(12367) := X"8E250014";
        ram_buffer(12368) := X"02002021";
        ram_buffer(12369) := X"0C022BF7";
        ram_buffer(12370) := X"00003021";
        ram_buffer(12371) := X"1000FF90";
        ram_buffer(12372) := X"00000000";
        ram_buffer(12373) := X"8E250014";
        ram_buffer(12374) := X"0C022BF7";
        ram_buffer(12375) := X"00003021";
        ram_buffer(12376) := X"8E250018";
        ram_buffer(12377) := X"24060001";
        ram_buffer(12378) := X"0C022BF7";
        ram_buffer(12379) := X"02002021";
        ram_buffer(12380) := X"8E0200EC";
        ram_buffer(12381) := X"1000FF6B";
        ram_buffer(12382) := X"28430002";
        ram_buffer(12383) := X"8E250018";
        ram_buffer(12384) := X"0C022BF7";
        ram_buffer(12385) := X"24060001";
        ram_buffer(12386) := X"8E0200EC";
        ram_buffer(12387) := X"1000FF65";
        ram_buffer(12388) := X"28430002";
        ram_buffer(12389) := X"8E250014";
        ram_buffer(12390) := X"00003021";
        ram_buffer(12391) := X"0C022BF7";
        ram_buffer(12392) := X"02002021";
        ram_buffer(12393) := X"8E0200EC";
        ram_buffer(12394) := X"1000FF80";
        ram_buffer(12395) := X"28420004";
        ram_buffer(12396) := X"8E250014";
        ram_buffer(12397) := X"0C022BF7";
        ram_buffer(12398) := X"02002021";
        ram_buffer(12399) := X"8E0200EC";
        ram_buffer(12400) := X"1000FF69";
        ram_buffer(12401) := X"28430003";
        ram_buffer(12402) := X"24A20010";
        ram_buffer(12403) := X"00021080";
        ram_buffer(12404) := X"27BDFFD0";
        ram_buffer(12405) := X"00821021";
        ram_buffer(12406) := X"AFB10014";
        ram_buffer(12407) := X"8C510000";
        ram_buffer(12408) := X"AFB50024";
        ram_buffer(12409) := X"AFB20018";
        ram_buffer(12410) := X"AFBF002C";
        ram_buffer(12411) := X"AFB60028";
        ram_buffer(12412) := X"AFB40020";
        ram_buffer(12413) := X"AFB3001C";
        ram_buffer(12414) := X"AFB00010";
        ram_buffer(12415) := X"00A09021";
        ram_buffer(12416) := X"122000F4";
        ram_buffer(12417) := X"0080A821";
        ram_buffer(12418) := X"02201021";
        ram_buffer(12419) := X"26260080";
        ram_buffer(12420) := X"00002021";
        ram_buffer(12421) := X"94430000";
        ram_buffer(12422) := X"00000000";
        ram_buffer(12423) := X"2C630100";
        ram_buffer(12424) := X"14600002";
        ram_buffer(12425) := X"00808021";
        ram_buffer(12426) := X"24100001";
        ram_buffer(12427) := X"24420002";
        ram_buffer(12428) := X"14C2FFF8";
        ram_buffer(12429) := X"02002021";
        ram_buffer(12430) := X"8E220080";
        ram_buffer(12431) := X"00000000";
        ram_buffer(12432) := X"1040000C";
        ram_buffer(12433) := X"00000000";
        ram_buffer(12434) := X"8FBF002C";
        ram_buffer(12435) := X"02001021";
        ram_buffer(12436) := X"8FB60028";
        ram_buffer(12437) := X"8FB50024";
        ram_buffer(12438) := X"8FB40020";
        ram_buffer(12439) := X"8FB3001C";
        ram_buffer(12440) := X"8FB20018";
        ram_buffer(12441) := X"8FB10014";
        ram_buffer(12442) := X"8FB00010";
        ram_buffer(12443) := X"03E00008";
        ram_buffer(12444) := X"27BD0030";
        ram_buffer(12445) := X"8EA20014";
        ram_buffer(12446) := X"00000000";
        ram_buffer(12447) := X"8C430000";
        ram_buffer(12448) := X"00000000";
        ram_buffer(12449) := X"24640001";
        ram_buffer(12450) := X"AC440000";
        ram_buffer(12451) := X"2404FFFF";
        ram_buffer(12452) := X"A0640000";
        ram_buffer(12453) := X"8C430004";
        ram_buffer(12454) := X"00000000";
        ram_buffer(12455) := X"2463FFFF";
        ram_buffer(12456) := X"106000A2";
        ram_buffer(12457) := X"AC430004";
        ram_buffer(12458) := X"8EA20014";
        ram_buffer(12459) := X"00000000";
        ram_buffer(12460) := X"8C430000";
        ram_buffer(12461) := X"00000000";
        ram_buffer(12462) := X"24640001";
        ram_buffer(12463) := X"AC440000";
        ram_buffer(12464) := X"2404FFDB";
        ram_buffer(12465) := X"A0640000";
        ram_buffer(12466) := X"8C430004";
        ram_buffer(12467) := X"00000000";
        ram_buffer(12468) := X"2463FFFF";
        ram_buffer(12469) := X"10600087";
        ram_buffer(12470) := X"AC430004";
        ram_buffer(12471) := X"1200006B";
        ram_buffer(12472) := X"24130043";
        ram_buffer(12473) := X"8EA20014";
        ram_buffer(12474) := X"24130083";
        ram_buffer(12475) := X"8C430000";
        ram_buffer(12476) := X"00000000";
        ram_buffer(12477) := X"24640001";
        ram_buffer(12478) := X"AC440000";
        ram_buffer(12479) := X"A0600000";
        ram_buffer(12480) := X"8C430004";
        ram_buffer(12481) := X"00000000";
        ram_buffer(12482) := X"2463FFFF";
        ram_buffer(12483) := X"1060006B";
        ram_buffer(12484) := X"AC430004";
        ram_buffer(12485) := X"8EA20014";
        ram_buffer(12486) := X"00000000";
        ram_buffer(12487) := X"8C430000";
        ram_buffer(12488) := X"00000000";
        ram_buffer(12489) := X"24640001";
        ram_buffer(12490) := X"AC440000";
        ram_buffer(12491) := X"A0730000";
        ram_buffer(12492) := X"8C430004";
        ram_buffer(12493) := X"00000000";
        ram_buffer(12494) := X"2463FFFF";
        ram_buffer(12495) := X"10600097";
        ram_buffer(12496) := X"AC430004";
        ram_buffer(12497) := X"8EA30014";
        ram_buffer(12498) := X"00101100";
        ram_buffer(12499) := X"8C640000";
        ram_buffer(12500) := X"00529021";
        ram_buffer(12501) := X"24820001";
        ram_buffer(12502) := X"AC620000";
        ram_buffer(12503) := X"A0920000";
        ram_buffer(12504) := X"8C620004";
        ram_buffer(12505) := X"00000000";
        ram_buffer(12506) := X"2442FFFF";
        ram_buffer(12507) := X"1040007D";
        ram_buffer(12508) := X"AC620004";
        ram_buffer(12509) := X"3C14100D";
        ram_buffer(12510) := X"3C12100D";
        ram_buffer(12511) := X"26948968";
        ram_buffer(12512) := X"26528A68";
        ram_buffer(12513) := X"24130016";
        ram_buffer(12514) := X"8E820000";
        ram_buffer(12515) := X"00000000";
        ram_buffer(12516) := X"00021040";
        ram_buffer(12517) := X"02221021";
        ram_buffer(12518) := X"94560000";
        ram_buffer(12519) := X"16000021";
        ram_buffer(12520) := X"26940004";
        ram_buffer(12521) := X"8EA20014";
        ram_buffer(12522) := X"00000000";
        ram_buffer(12523) := X"8C430000";
        ram_buffer(12524) := X"00000000";
        ram_buffer(12525) := X"24640001";
        ram_buffer(12526) := X"AC440000";
        ram_buffer(12527) := X"A0760000";
        ram_buffer(12528) := X"8C430004";
        ram_buffer(12529) := X"00000000";
        ram_buffer(12530) := X"2463FFFF";
        ram_buffer(12531) := X"10600005";
        ram_buffer(12532) := X"AC430004";
        ram_buffer(12533) := X"1654FFEC";
        ram_buffer(12534) := X"24020001";
        ram_buffer(12535) := X"1000FF9A";
        ram_buffer(12536) := X"AE220080";
        ram_buffer(12537) := X"8C42000C";
        ram_buffer(12538) := X"00000000";
        ram_buffer(12539) := X"0040F809";
        ram_buffer(12540) := X"02A02021";
        ram_buffer(12541) := X"1440FFF7";
        ram_buffer(12542) := X"02A02021";
        ram_buffer(12543) := X"8EA20000";
        ram_buffer(12544) := X"00000000";
        ram_buffer(12545) := X"8C430000";
        ram_buffer(12546) := X"00000000";
        ram_buffer(12547) := X"0060F809";
        ram_buffer(12548) := X"AC530014";
        ram_buffer(12549) := X"1654FFDC";
        ram_buffer(12550) := X"24020001";
        ram_buffer(12551) := X"1000FF8A";
        ram_buffer(12552) := X"AE220080";
        ram_buffer(12553) := X"8EA20014";
        ram_buffer(12554) := X"00161A02";
        ram_buffer(12555) := X"8C440000";
        ram_buffer(12556) := X"00000000";
        ram_buffer(12557) := X"24850001";
        ram_buffer(12558) := X"AC450000";
        ram_buffer(12559) := X"A0830000";
        ram_buffer(12560) := X"8C430004";
        ram_buffer(12561) := X"00000000";
        ram_buffer(12562) := X"2463FFFF";
        ram_buffer(12563) := X"1460FFD5";
        ram_buffer(12564) := X"AC430004";
        ram_buffer(12565) := X"8C42000C";
        ram_buffer(12566) := X"00000000";
        ram_buffer(12567) := X"0040F809";
        ram_buffer(12568) := X"02A02021";
        ram_buffer(12569) := X"1440FFCF";
        ram_buffer(12570) := X"02A02021";
        ram_buffer(12571) := X"8EA20000";
        ram_buffer(12572) := X"00000000";
        ram_buffer(12573) := X"8C430000";
        ram_buffer(12574) := X"00000000";
        ram_buffer(12575) := X"0060F809";
        ram_buffer(12576) := X"AC530014";
        ram_buffer(12577) := X"1000FFC7";
        ram_buffer(12578) := X"00000000";
        ram_buffer(12579) := X"8EA20014";
        ram_buffer(12580) := X"00000000";
        ram_buffer(12581) := X"8C430000";
        ram_buffer(12582) := X"00000000";
        ram_buffer(12583) := X"24640001";
        ram_buffer(12584) := X"AC440000";
        ram_buffer(12585) := X"A0600000";
        ram_buffer(12586) := X"8C430004";
        ram_buffer(12587) := X"00000000";
        ram_buffer(12588) := X"2463FFFF";
        ram_buffer(12589) := X"1460FF97";
        ram_buffer(12590) := X"AC430004";
        ram_buffer(12591) := X"8C42000C";
        ram_buffer(12592) := X"00000000";
        ram_buffer(12593) := X"0040F809";
        ram_buffer(12594) := X"02A02021";
        ram_buffer(12595) := X"1440FF91";
        ram_buffer(12596) := X"24040016";
        ram_buffer(12597) := X"8EA20000";
        ram_buffer(12598) := X"00000000";
        ram_buffer(12599) := X"8C430000";
        ram_buffer(12600) := X"AC440014";
        ram_buffer(12601) := X"0060F809";
        ram_buffer(12602) := X"02A02021";
        ram_buffer(12603) := X"1000FF89";
        ram_buffer(12604) := X"00000000";
        ram_buffer(12605) := X"8C42000C";
        ram_buffer(12606) := X"00000000";
        ram_buffer(12607) := X"0040F809";
        ram_buffer(12608) := X"02A02021";
        ram_buffer(12609) := X"1440FF75";
        ram_buffer(12610) := X"24040016";
        ram_buffer(12611) := X"8EA20000";
        ram_buffer(12612) := X"00000000";
        ram_buffer(12613) := X"8C430000";
        ram_buffer(12614) := X"AC440014";
        ram_buffer(12615) := X"0060F809";
        ram_buffer(12616) := X"02A02021";
        ram_buffer(12617) := X"1000FF6D";
        ram_buffer(12618) := X"00000000";
        ram_buffer(12619) := X"8C42000C";
        ram_buffer(12620) := X"00000000";
        ram_buffer(12621) := X"0040F809";
        ram_buffer(12622) := X"02A02021";
        ram_buffer(12623) := X"1440FF5A";
        ram_buffer(12624) := X"24040016";
        ram_buffer(12625) := X"8EA20000";
        ram_buffer(12626) := X"00000000";
        ram_buffer(12627) := X"8C430000";
        ram_buffer(12628) := X"AC440014";
        ram_buffer(12629) := X"0060F809";
        ram_buffer(12630) := X"02A02021";
        ram_buffer(12631) := X"1000FF52";
        ram_buffer(12632) := X"00000000";
        ram_buffer(12633) := X"8C62000C";
        ram_buffer(12634) := X"00000000";
        ram_buffer(12635) := X"0040F809";
        ram_buffer(12636) := X"02A02021";
        ram_buffer(12637) := X"1440FF7F";
        ram_buffer(12638) := X"24040016";
        ram_buffer(12639) := X"8EA20000";
        ram_buffer(12640) := X"00000000";
        ram_buffer(12641) := X"8C430000";
        ram_buffer(12642) := X"AC440014";
        ram_buffer(12643) := X"0060F809";
        ram_buffer(12644) := X"02A02021";
        ram_buffer(12645) := X"1000FF78";
        ram_buffer(12646) := X"3C14100D";
        ram_buffer(12647) := X"8C42000C";
        ram_buffer(12648) := X"00000000";
        ram_buffer(12649) := X"0040F809";
        ram_buffer(12650) := X"02A02021";
        ram_buffer(12651) := X"1440FF65";
        ram_buffer(12652) := X"24040016";
        ram_buffer(12653) := X"8EA20000";
        ram_buffer(12654) := X"00000000";
        ram_buffer(12655) := X"8C430000";
        ram_buffer(12656) := X"AC440014";
        ram_buffer(12657) := X"0060F809";
        ram_buffer(12658) := X"02A02021";
        ram_buffer(12659) := X"1000FF5D";
        ram_buffer(12660) := X"00000000";
        ram_buffer(12661) := X"8C820000";
        ram_buffer(12662) := X"00000000";
        ram_buffer(12663) := X"AC450018";
        ram_buffer(12664) := X"8C830000";
        ram_buffer(12665) := X"24050033";
        ram_buffer(12666) := X"AC450014";
        ram_buffer(12667) := X"8C620000";
        ram_buffer(12668) := X"00000000";
        ram_buffer(12669) := X"0040F809";
        ram_buffer(12670) := X"00000000";
        ram_buffer(12671) := X"1000FF03";
        ram_buffer(12672) := X"02201021";
        ram_buffer(12673) := X"8C830034";
        ram_buffer(12674) := X"27BDFFD8";
        ram_buffer(12675) := X"AFB30020";
        ram_buffer(12676) := X"AFB2001C";
        ram_buffer(12677) := X"AFB00014";
        ram_buffer(12678) := X"AFBF0024";
        ram_buffer(12679) := X"AFB10018";
        ram_buffer(12680) := X"00809021";
        ram_buffer(12681) := X"8C90003C";
        ram_buffer(12682) := X"1860000B";
        ram_buffer(12683) := X"00009821";
        ram_buffer(12684) := X"00008821";
        ram_buffer(12685) := X"8E050010";
        ram_buffer(12686) := X"0C023072";
        ram_buffer(12687) := X"02402021";
        ram_buffer(12688) := X"8E430034";
        ram_buffer(12689) := X"26310001";
        ram_buffer(12690) := X"0223202A";
        ram_buffer(12691) := X"02629821";
        ram_buffer(12692) := X"1480FFF8";
        ram_buffer(12693) := X"26100054";
        ram_buffer(12694) := X"8E4200AC";
        ram_buffer(12695) := X"00000000";
        ram_buffer(12696) := X"1040000A";
        ram_buffer(12697) := X"00000000";
        ram_buffer(12698) := X"8FBF0024";
        ram_buffer(12699) := X"8FB30020";
        ram_buffer(12700) := X"8FB10018";
        ram_buffer(12701) := X"8FB00014";
        ram_buffer(12702) := X"02402021";
        ram_buffer(12703) := X"8FB2001C";
        ram_buffer(12704) := X"240500C9";
        ram_buffer(12705) := X"08022A29";
        ram_buffer(12706) := X"27BD0028";
        ram_buffer(12707) := X"8E4200DC";
        ram_buffer(12708) := X"00000000";
        ram_buffer(12709) := X"1040000A";
        ram_buffer(12710) := X"24020008";
        ram_buffer(12711) := X"8FBF0024";
        ram_buffer(12712) := X"8FB30020";
        ram_buffer(12713) := X"8FB10018";
        ram_buffer(12714) := X"8FB00014";
        ram_buffer(12715) := X"02402021";
        ram_buffer(12716) := X"8FB2001C";
        ram_buffer(12717) := X"240500C2";
        ram_buffer(12718) := X"08022A29";
        ram_buffer(12719) := X"27BD0028";
        ram_buffer(12720) := X"8E440030";
        ram_buffer(12721) := X"00000000";
        ram_buffer(12722) := X"1082000A";
        ram_buffer(12723) := X"00000000";
        ram_buffer(12724) := X"240500C1";
        ram_buffer(12725) := X"8FBF0024";
        ram_buffer(12726) := X"8FB30020";
        ram_buffer(12727) := X"8FB10018";
        ram_buffer(12728) := X"8FB00014";
        ram_buffer(12729) := X"02402021";
        ram_buffer(12730) := X"8FB2001C";
        ram_buffer(12731) := X"08022A29";
        ram_buffer(12732) := X"27BD0028";
        ram_buffer(12733) := X"8E44003C";
        ram_buffer(12734) := X"18600031";
        ram_buffer(12735) := X"24060001";
        ram_buffer(12736) := X"00002821";
        ram_buffer(12737) := X"8C820014";
        ram_buffer(12738) := X"00000000";
        ram_buffer(12739) := X"28420002";
        ram_buffer(12740) := X"1440001A";
        ram_buffer(12741) := X"00000000";
        ram_buffer(12742) := X"00003021";
        ram_buffer(12743) := X"24A50001";
        ram_buffer(12744) := X"14A3FFF8";
        ram_buffer(12745) := X"24840054";
        ram_buffer(12746) := X"1260001B";
        ram_buffer(12747) := X"00000000";
        ram_buffer(12748) := X"10C0FFE8";
        ram_buffer(12749) := X"240500C1";
        ram_buffer(12750) := X"8E420000";
        ram_buffer(12751) := X"2404004A";
        ram_buffer(12752) := X"8C430004";
        ram_buffer(12753) := X"AC440014";
        ram_buffer(12754) := X"00002821";
        ram_buffer(12755) := X"0060F809";
        ram_buffer(12756) := X"02402021";
        ram_buffer(12757) := X"8E4200AC";
        ram_buffer(12758) := X"00000000";
        ram_buffer(12759) := X"1440FFC2";
        ram_buffer(12760) := X"00000000";
        ram_buffer(12761) := X"8E4200DC";
        ram_buffer(12762) := X"00000000";
        ram_buffer(12763) := X"1440FFCB";
        ram_buffer(12764) := X"240500C1";
        ram_buffer(12765) := X"1000FFD7";
        ram_buffer(12766) := X"00000000";
        ram_buffer(12767) := X"8C820018";
        ram_buffer(12768) := X"00000000";
        ram_buffer(12769) := X"28420002";
        ram_buffer(12770) := X"1040FFE3";
        ram_buffer(12771) := X"00000000";
        ram_buffer(12772) := X"1000FFE3";
        ram_buffer(12773) := X"24A50001";
        ram_buffer(12774) := X"10C0FFCD";
        ram_buffer(12775) := X"240500C0";
        ram_buffer(12776) := X"8FBF0024";
        ram_buffer(12777) := X"8FB30020";
        ram_buffer(12778) := X"8FB10018";
        ram_buffer(12779) := X"8FB00014";
        ram_buffer(12780) := X"02402021";
        ram_buffer(12781) := X"8FB2001C";
        ram_buffer(12782) := X"08022A29";
        ram_buffer(12783) := X"27BD0028";
        ram_buffer(12784) := X"1660FFDD";
        ram_buffer(12785) := X"240500C0";
        ram_buffer(12786) := X"1000FFF5";
        ram_buffer(12787) := X"00000000";
        ram_buffer(12788) := X"8C820014";
        ram_buffer(12789) := X"27BDFFD8";
        ram_buffer(12790) := X"8C430000";
        ram_buffer(12791) := X"AFB00014";
        ram_buffer(12792) := X"24650001";
        ram_buffer(12793) := X"AFBF0024";
        ram_buffer(12794) := X"AFB30020";
        ram_buffer(12795) := X"AFB2001C";
        ram_buffer(12796) := X"AFB10018";
        ram_buffer(12797) := X"AC450000";
        ram_buffer(12798) := X"2405FFFF";
        ram_buffer(12799) := X"A0650000";
        ram_buffer(12800) := X"8C430004";
        ram_buffer(12801) := X"00808021";
        ram_buffer(12802) := X"2463FFFF";
        ram_buffer(12803) := X"10600053";
        ram_buffer(12804) := X"AC430004";
        ram_buffer(12805) := X"8E020014";
        ram_buffer(12806) := X"00000000";
        ram_buffer(12807) := X"8C430000";
        ram_buffer(12808) := X"00000000";
        ram_buffer(12809) := X"24640001";
        ram_buffer(12810) := X"AC440000";
        ram_buffer(12811) := X"2404FFD8";
        ram_buffer(12812) := X"A0640000";
        ram_buffer(12813) := X"8C430004";
        ram_buffer(12814) := X"00000000";
        ram_buffer(12815) := X"2463FFFF";
        ram_buffer(12816) := X"1060005F";
        ram_buffer(12817) := X"AC430004";
        ram_buffer(12818) := X"26120040";
        ram_buffer(12819) := X"00008821";
        ram_buffer(12820) := X"24130004";
        ram_buffer(12821) := X"8E420000";
        ram_buffer(12822) := X"02202821";
        ram_buffer(12823) := X"02002021";
        ram_buffer(12824) := X"10400003";
        ram_buffer(12825) := X"26310001";
        ram_buffer(12826) := X"0C023072";
        ram_buffer(12827) := X"00000000";
        ram_buffer(12828) := X"1633FFF8";
        ram_buffer(12829) := X"26520004";
        ram_buffer(12830) := X"8E0200AC";
        ram_buffer(12831) := X"00000000";
        ram_buffer(12832) := X"14400015";
        ram_buffer(12833) := X"00000000";
        ram_buffer(12834) := X"26120050";
        ram_buffer(12835) := X"00008821";
        ram_buffer(12836) := X"24130004";
        ram_buffer(12837) := X"8E420000";
        ram_buffer(12838) := X"02202821";
        ram_buffer(12839) := X"02002021";
        ram_buffer(12840) := X"10400003";
        ram_buffer(12841) := X"00003021";
        ram_buffer(12842) := X"0C022BF7";
        ram_buffer(12843) := X"00000000";
        ram_buffer(12844) := X"8E420010";
        ram_buffer(12845) := X"02202821";
        ram_buffer(12846) := X"24060001";
        ram_buffer(12847) := X"26310001";
        ram_buffer(12848) := X"10400003";
        ram_buffer(12849) := X"02002021";
        ram_buffer(12850) := X"0C022BF7";
        ram_buffer(12851) := X"00000000";
        ram_buffer(12852) := X"1633FFF0";
        ram_buffer(12853) := X"26520004";
        ram_buffer(12854) := X"8E020014";
        ram_buffer(12855) := X"00000000";
        ram_buffer(12856) := X"8C430000";
        ram_buffer(12857) := X"00000000";
        ram_buffer(12858) := X"24640001";
        ram_buffer(12859) := X"AC440000";
        ram_buffer(12860) := X"2404FFFF";
        ram_buffer(12861) := X"A0640000";
        ram_buffer(12862) := X"8C430004";
        ram_buffer(12863) := X"00000000";
        ram_buffer(12864) := X"2463FFFF";
        ram_buffer(12865) := X"1060004D";
        ram_buffer(12866) := X"AC430004";
        ram_buffer(12867) := X"8E020014";
        ram_buffer(12868) := X"00000000";
        ram_buffer(12869) := X"8C430000";
        ram_buffer(12870) := X"00000000";
        ram_buffer(12871) := X"24640001";
        ram_buffer(12872) := X"AC440000";
        ram_buffer(12873) := X"2404FFD9";
        ram_buffer(12874) := X"A0640000";
        ram_buffer(12875) := X"8C430004";
        ram_buffer(12876) := X"00000000";
        ram_buffer(12877) := X"2463FFFF";
        ram_buffer(12878) := X"1060002F";
        ram_buffer(12879) := X"AC430004";
        ram_buffer(12880) := X"8FBF0024";
        ram_buffer(12881) := X"8FB30020";
        ram_buffer(12882) := X"8FB2001C";
        ram_buffer(12883) := X"8FB10018";
        ram_buffer(12884) := X"8FB00014";
        ram_buffer(12885) := X"03E00008";
        ram_buffer(12886) := X"27BD0028";
        ram_buffer(12887) := X"8C42000C";
        ram_buffer(12888) := X"00000000";
        ram_buffer(12889) := X"0040F809";
        ram_buffer(12890) := X"00000000";
        ram_buffer(12891) := X"1440FFA9";
        ram_buffer(12892) := X"24040016";
        ram_buffer(12893) := X"8E020000";
        ram_buffer(12894) := X"00000000";
        ram_buffer(12895) := X"8C430000";
        ram_buffer(12896) := X"AC440014";
        ram_buffer(12897) := X"0060F809";
        ram_buffer(12898) := X"02002021";
        ram_buffer(12899) := X"8E020014";
        ram_buffer(12900) := X"00000000";
        ram_buffer(12901) := X"8C430000";
        ram_buffer(12902) := X"00000000";
        ram_buffer(12903) := X"24640001";
        ram_buffer(12904) := X"AC440000";
        ram_buffer(12905) := X"2404FFD8";
        ram_buffer(12906) := X"A0640000";
        ram_buffer(12907) := X"8C430004";
        ram_buffer(12908) := X"00000000";
        ram_buffer(12909) := X"2463FFFF";
        ram_buffer(12910) := X"1460FFA3";
        ram_buffer(12911) := X"AC430004";
        ram_buffer(12912) := X"8C42000C";
        ram_buffer(12913) := X"00000000";
        ram_buffer(12914) := X"0040F809";
        ram_buffer(12915) := X"02002021";
        ram_buffer(12916) := X"1440FF9D";
        ram_buffer(12917) := X"24040016";
        ram_buffer(12918) := X"8E020000";
        ram_buffer(12919) := X"00000000";
        ram_buffer(12920) := X"8C430000";
        ram_buffer(12921) := X"AC440014";
        ram_buffer(12922) := X"0060F809";
        ram_buffer(12923) := X"02002021";
        ram_buffer(12924) := X"1000FF96";
        ram_buffer(12925) := X"26120040";
        ram_buffer(12926) := X"8C42000C";
        ram_buffer(12927) := X"00000000";
        ram_buffer(12928) := X"0040F809";
        ram_buffer(12929) := X"02002021";
        ram_buffer(12930) := X"1440FFCD";
        ram_buffer(12931) := X"24030016";
        ram_buffer(12932) := X"8E020000";
        ram_buffer(12933) := X"8FBF0024";
        ram_buffer(12934) := X"8FB30020";
        ram_buffer(12935) := X"8FB2001C";
        ram_buffer(12936) := X"8FB10018";
        ram_buffer(12937) := X"8C590000";
        ram_buffer(12938) := X"02002021";
        ram_buffer(12939) := X"8FB00014";
        ram_buffer(12940) := X"AC430014";
        ram_buffer(12941) := X"03200008";
        ram_buffer(12942) := X"27BD0028";
        ram_buffer(12943) := X"8C42000C";
        ram_buffer(12944) := X"00000000";
        ram_buffer(12945) := X"0040F809";
        ram_buffer(12946) := X"02002021";
        ram_buffer(12947) := X"1440FFAF";
        ram_buffer(12948) := X"24040016";
        ram_buffer(12949) := X"8E020000";
        ram_buffer(12950) := X"00000000";
        ram_buffer(12951) := X"8C430000";
        ram_buffer(12952) := X"AC440014";
        ram_buffer(12953) := X"0060F809";
        ram_buffer(12954) := X"02002021";
        ram_buffer(12955) := X"1000FFA7";
        ram_buffer(12956) := X"00000000";
        ram_buffer(12957) := X"8C820014";
        ram_buffer(12958) := X"27BDFFE0";
        ram_buffer(12959) := X"8C430000";
        ram_buffer(12960) := X"AFB00014";
        ram_buffer(12961) := X"24650001";
        ram_buffer(12962) := X"AFBF001C";
        ram_buffer(12963) := X"AFB10018";
        ram_buffer(12964) := X"AC450000";
        ram_buffer(12965) := X"2405FFFF";
        ram_buffer(12966) := X"A0650000";
        ram_buffer(12967) := X"8C430004";
        ram_buffer(12968) := X"00808021";
        ram_buffer(12969) := X"2463FFFF";
        ram_buffer(12970) := X"1060001B";
        ram_buffer(12971) := X"AC430004";
        ram_buffer(12972) := X"8E020014";
        ram_buffer(12973) := X"00000000";
        ram_buffer(12974) := X"8C430000";
        ram_buffer(12975) := X"00000000";
        ram_buffer(12976) := X"24640001";
        ram_buffer(12977) := X"AC440000";
        ram_buffer(12978) := X"2404FFD8";
        ram_buffer(12979) := X"A0640000";
        ram_buffer(12980) := X"8C430004";
        ram_buffer(12981) := X"00000000";
        ram_buffer(12982) := X"2463FFFF";
        ram_buffer(12983) := X"10600027";
        ram_buffer(12984) := X"AC430004";
        ram_buffer(12985) := X"8E0200C8";
        ram_buffer(12986) := X"00000000";
        ram_buffer(12987) := X"14400033";
        ram_buffer(12988) := X"00000000";
        ram_buffer(12989) := X"8E0200D4";
        ram_buffer(12990) := X"00000000";
        ram_buffer(12991) := X"1440011E";
        ram_buffer(12992) := X"00000000";
        ram_buffer(12993) := X"8FBF001C";
        ram_buffer(12994) := X"8FB10018";
        ram_buffer(12995) := X"8FB00014";
        ram_buffer(12996) := X"03E00008";
        ram_buffer(12997) := X"27BD0020";
        ram_buffer(12998) := X"8C42000C";
        ram_buffer(12999) := X"00000000";
        ram_buffer(13000) := X"0040F809";
        ram_buffer(13001) := X"00000000";
        ram_buffer(13002) := X"1440FFE1";
        ram_buffer(13003) := X"24040016";
        ram_buffer(13004) := X"8E020000";
        ram_buffer(13005) := X"00000000";
        ram_buffer(13006) := X"8C430000";
        ram_buffer(13007) := X"AC440014";
        ram_buffer(13008) := X"0060F809";
        ram_buffer(13009) := X"02002021";
        ram_buffer(13010) := X"8E020014";
        ram_buffer(13011) := X"00000000";
        ram_buffer(13012) := X"8C430000";
        ram_buffer(13013) := X"00000000";
        ram_buffer(13014) := X"24640001";
        ram_buffer(13015) := X"AC440000";
        ram_buffer(13016) := X"2404FFD8";
        ram_buffer(13017) := X"A0640000";
        ram_buffer(13018) := X"8C430004";
        ram_buffer(13019) := X"00000000";
        ram_buffer(13020) := X"2463FFFF";
        ram_buffer(13021) := X"1460FFDB";
        ram_buffer(13022) := X"AC430004";
        ram_buffer(13023) := X"8C42000C";
        ram_buffer(13024) := X"00000000";
        ram_buffer(13025) := X"0040F809";
        ram_buffer(13026) := X"02002021";
        ram_buffer(13027) := X"1440FFD5";
        ram_buffer(13028) := X"24040016";
        ram_buffer(13029) := X"8E020000";
        ram_buffer(13030) := X"00000000";
        ram_buffer(13031) := X"8C430000";
        ram_buffer(13032) := X"AC440014";
        ram_buffer(13033) := X"0060F809";
        ram_buffer(13034) := X"02002021";
        ram_buffer(13035) := X"8E0200C8";
        ram_buffer(13036) := X"00000000";
        ram_buffer(13037) := X"1040FFCF";
        ram_buffer(13038) := X"00000000";
        ram_buffer(13039) := X"8E020014";
        ram_buffer(13040) := X"00000000";
        ram_buffer(13041) := X"8C430000";
        ram_buffer(13042) := X"00000000";
        ram_buffer(13043) := X"24640001";
        ram_buffer(13044) := X"AC440000";
        ram_buffer(13045) := X"2404FFFF";
        ram_buffer(13046) := X"A0640000";
        ram_buffer(13047) := X"8C430004";
        ram_buffer(13048) := X"00000000";
        ram_buffer(13049) := X"2463FFFF";
        ram_buffer(13050) := X"106002B1";
        ram_buffer(13051) := X"AC430004";
        ram_buffer(13052) := X"8E020014";
        ram_buffer(13053) := X"00000000";
        ram_buffer(13054) := X"8C430000";
        ram_buffer(13055) := X"00000000";
        ram_buffer(13056) := X"24640001";
        ram_buffer(13057) := X"AC440000";
        ram_buffer(13058) := X"2404FFE0";
        ram_buffer(13059) := X"A0640000";
        ram_buffer(13060) := X"8C430004";
        ram_buffer(13061) := X"00000000";
        ram_buffer(13062) := X"2463FFFF";
        ram_buffer(13063) := X"10600296";
        ram_buffer(13064) := X"AC430004";
        ram_buffer(13065) := X"8E020014";
        ram_buffer(13066) := X"00000000";
        ram_buffer(13067) := X"8C430000";
        ram_buffer(13068) := X"00000000";
        ram_buffer(13069) := X"24640001";
        ram_buffer(13070) := X"AC440000";
        ram_buffer(13071) := X"A0600000";
        ram_buffer(13072) := X"8C430004";
        ram_buffer(13073) := X"00000000";
        ram_buffer(13074) := X"2463FFFF";
        ram_buffer(13075) := X"1060027C";
        ram_buffer(13076) := X"AC430004";
        ram_buffer(13077) := X"8E020014";
        ram_buffer(13078) := X"00000000";
        ram_buffer(13079) := X"8C430000";
        ram_buffer(13080) := X"00000000";
        ram_buffer(13081) := X"24640001";
        ram_buffer(13082) := X"AC440000";
        ram_buffer(13083) := X"24040010";
        ram_buffer(13084) := X"A0640000";
        ram_buffer(13085) := X"8C430004";
        ram_buffer(13086) := X"00000000";
        ram_buffer(13087) := X"2463FFFF";
        ram_buffer(13088) := X"10600261";
        ram_buffer(13089) := X"AC430004";
        ram_buffer(13090) := X"8E020014";
        ram_buffer(13091) := X"00000000";
        ram_buffer(13092) := X"8C430000";
        ram_buffer(13093) := X"00000000";
        ram_buffer(13094) := X"24640001";
        ram_buffer(13095) := X"AC440000";
        ram_buffer(13096) := X"2404004A";
        ram_buffer(13097) := X"A0640000";
        ram_buffer(13098) := X"8C430004";
        ram_buffer(13099) := X"00000000";
        ram_buffer(13100) := X"2463FFFF";
        ram_buffer(13101) := X"10600246";
        ram_buffer(13102) := X"AC430004";
        ram_buffer(13103) := X"8E020014";
        ram_buffer(13104) := X"00000000";
        ram_buffer(13105) := X"8C430000";
        ram_buffer(13106) := X"00000000";
        ram_buffer(13107) := X"24640001";
        ram_buffer(13108) := X"AC440000";
        ram_buffer(13109) := X"24040046";
        ram_buffer(13110) := X"A0640000";
        ram_buffer(13111) := X"8C430004";
        ram_buffer(13112) := X"00000000";
        ram_buffer(13113) := X"2463FFFF";
        ram_buffer(13114) := X"1060022B";
        ram_buffer(13115) := X"AC430004";
        ram_buffer(13116) := X"8E020014";
        ram_buffer(13117) := X"00000000";
        ram_buffer(13118) := X"8C430000";
        ram_buffer(13119) := X"00000000";
        ram_buffer(13120) := X"24640001";
        ram_buffer(13121) := X"AC440000";
        ram_buffer(13122) := X"24040049";
        ram_buffer(13123) := X"A0640000";
        ram_buffer(13124) := X"8C430004";
        ram_buffer(13125) := X"00000000";
        ram_buffer(13126) := X"2463FFFF";
        ram_buffer(13127) := X"10600210";
        ram_buffer(13128) := X"AC430004";
        ram_buffer(13129) := X"8E020014";
        ram_buffer(13130) := X"00000000";
        ram_buffer(13131) := X"8C430000";
        ram_buffer(13132) := X"00000000";
        ram_buffer(13133) := X"24640001";
        ram_buffer(13134) := X"AC440000";
        ram_buffer(13135) := X"24040046";
        ram_buffer(13136) := X"A0640000";
        ram_buffer(13137) := X"8C430004";
        ram_buffer(13138) := X"00000000";
        ram_buffer(13139) := X"2463FFFF";
        ram_buffer(13140) := X"106001F5";
        ram_buffer(13141) := X"AC430004";
        ram_buffer(13142) := X"8E020014";
        ram_buffer(13143) := X"00000000";
        ram_buffer(13144) := X"8C430000";
        ram_buffer(13145) := X"00000000";
        ram_buffer(13146) := X"24640001";
        ram_buffer(13147) := X"AC440000";
        ram_buffer(13148) := X"A0600000";
        ram_buffer(13149) := X"8C430004";
        ram_buffer(13150) := X"00000000";
        ram_buffer(13151) := X"2463FFFF";
        ram_buffer(13152) := X"106001DB";
        ram_buffer(13153) := X"AC430004";
        ram_buffer(13154) := X"8E020014";
        ram_buffer(13155) := X"00000000";
        ram_buffer(13156) := X"8C430000";
        ram_buffer(13157) := X"00000000";
        ram_buffer(13158) := X"24640001";
        ram_buffer(13159) := X"AC440000";
        ram_buffer(13160) := X"24040001";
        ram_buffer(13161) := X"A0640000";
        ram_buffer(13162) := X"8C430004";
        ram_buffer(13163) := X"00000000";
        ram_buffer(13164) := X"2463FFFF";
        ram_buffer(13165) := X"106001C0";
        ram_buffer(13166) := X"AC430004";
        ram_buffer(13167) := X"8E020014";
        ram_buffer(13168) := X"00000000";
        ram_buffer(13169) := X"8C430000";
        ram_buffer(13170) := X"00000000";
        ram_buffer(13171) := X"24640001";
        ram_buffer(13172) := X"AC440000";
        ram_buffer(13173) := X"24040001";
        ram_buffer(13174) := X"A0640000";
        ram_buffer(13175) := X"8C430004";
        ram_buffer(13176) := X"00000000";
        ram_buffer(13177) := X"2463FFFF";
        ram_buffer(13178) := X"106001A5";
        ram_buffer(13179) := X"AC430004";
        ram_buffer(13180) := X"8E020014";
        ram_buffer(13181) := X"920400CC";
        ram_buffer(13182) := X"8C430000";
        ram_buffer(13183) := X"00000000";
        ram_buffer(13184) := X"24650001";
        ram_buffer(13185) := X"AC450000";
        ram_buffer(13186) := X"A0640000";
        ram_buffer(13187) := X"8C430004";
        ram_buffer(13188) := X"00000000";
        ram_buffer(13189) := X"2463FFFF";
        ram_buffer(13190) := X"1060018B";
        ram_buffer(13191) := X"AC430004";
        ram_buffer(13192) := X"8E020014";
        ram_buffer(13193) := X"961100CE";
        ram_buffer(13194) := X"8C430000";
        ram_buffer(13195) := X"00112203";
        ram_buffer(13196) := X"24650001";
        ram_buffer(13197) := X"AC450000";
        ram_buffer(13198) := X"A0640000";
        ram_buffer(13199) := X"8C430004";
        ram_buffer(13200) := X"00000000";
        ram_buffer(13201) := X"2463FFFF";
        ram_buffer(13202) := X"10600171";
        ram_buffer(13203) := X"AC430004";
        ram_buffer(13204) := X"8E020014";
        ram_buffer(13205) := X"00000000";
        ram_buffer(13206) := X"8C430000";
        ram_buffer(13207) := X"00000000";
        ram_buffer(13208) := X"24640001";
        ram_buffer(13209) := X"AC440000";
        ram_buffer(13210) := X"A0710000";
        ram_buffer(13211) := X"8C430004";
        ram_buffer(13212) := X"00000000";
        ram_buffer(13213) := X"2463FFFF";
        ram_buffer(13214) := X"10600157";
        ram_buffer(13215) := X"AC430004";
        ram_buffer(13216) := X"8E020014";
        ram_buffer(13217) := X"961100D0";
        ram_buffer(13218) := X"8C430000";
        ram_buffer(13219) := X"00112203";
        ram_buffer(13220) := X"24650001";
        ram_buffer(13221) := X"AC450000";
        ram_buffer(13222) := X"A0640000";
        ram_buffer(13223) := X"8C430004";
        ram_buffer(13224) := X"00000000";
        ram_buffer(13225) := X"2463FFFF";
        ram_buffer(13226) := X"1060013D";
        ram_buffer(13227) := X"AC430004";
        ram_buffer(13228) := X"8E020014";
        ram_buffer(13229) := X"00000000";
        ram_buffer(13230) := X"8C430000";
        ram_buffer(13231) := X"00000000";
        ram_buffer(13232) := X"24640001";
        ram_buffer(13233) := X"AC440000";
        ram_buffer(13234) := X"A0710000";
        ram_buffer(13235) := X"8C430004";
        ram_buffer(13236) := X"00000000";
        ram_buffer(13237) := X"2463FFFF";
        ram_buffer(13238) := X"10600123";
        ram_buffer(13239) := X"AC430004";
        ram_buffer(13240) := X"8E020014";
        ram_buffer(13241) := X"00000000";
        ram_buffer(13242) := X"8C430000";
        ram_buffer(13243) := X"00000000";
        ram_buffer(13244) := X"24640001";
        ram_buffer(13245) := X"AC440000";
        ram_buffer(13246) := X"A0600000";
        ram_buffer(13247) := X"8C430004";
        ram_buffer(13248) := X"00000000";
        ram_buffer(13249) := X"2463FFFF";
        ram_buffer(13250) := X"10600109";
        ram_buffer(13251) := X"AC430004";
        ram_buffer(13252) := X"8E020014";
        ram_buffer(13253) := X"00000000";
        ram_buffer(13254) := X"8C430000";
        ram_buffer(13255) := X"00000000";
        ram_buffer(13256) := X"24640001";
        ram_buffer(13257) := X"AC440000";
        ram_buffer(13258) := X"A0600000";
        ram_buffer(13259) := X"8C430004";
        ram_buffer(13260) := X"00000000";
        ram_buffer(13261) := X"2463FFFF";
        ram_buffer(13262) := X"1460FEEE";
        ram_buffer(13263) := X"AC430004";
        ram_buffer(13264) := X"8C42000C";
        ram_buffer(13265) := X"00000000";
        ram_buffer(13266) := X"0040F809";
        ram_buffer(13267) := X"02002021";
        ram_buffer(13268) := X"1440FEE8";
        ram_buffer(13269) := X"24040016";
        ram_buffer(13270) := X"8E020000";
        ram_buffer(13271) := X"00000000";
        ram_buffer(13272) := X"8C430000";
        ram_buffer(13273) := X"AC440014";
        ram_buffer(13274) := X"0060F809";
        ram_buffer(13275) := X"02002021";
        ram_buffer(13276) := X"1000FEE0";
        ram_buffer(13277) := X"00000000";
        ram_buffer(13278) := X"8E020014";
        ram_buffer(13279) := X"00000000";
        ram_buffer(13280) := X"8C430000";
        ram_buffer(13281) := X"00000000";
        ram_buffer(13282) := X"24640001";
        ram_buffer(13283) := X"AC440000";
        ram_buffer(13284) := X"2404FFFF";
        ram_buffer(13285) := X"A0640000";
        ram_buffer(13286) := X"8C430004";
        ram_buffer(13287) := X"00000000";
        ram_buffer(13288) := X"2463FFFF";
        ram_buffer(13289) := X"106001EC";
        ram_buffer(13290) := X"AC430004";
        ram_buffer(13291) := X"8E020014";
        ram_buffer(13292) := X"00000000";
        ram_buffer(13293) := X"8C430000";
        ram_buffer(13294) := X"00000000";
        ram_buffer(13295) := X"24640001";
        ram_buffer(13296) := X"AC440000";
        ram_buffer(13297) := X"2404FFEE";
        ram_buffer(13298) := X"A0640000";
        ram_buffer(13299) := X"8C430004";
        ram_buffer(13300) := X"00000000";
        ram_buffer(13301) := X"2463FFFF";
        ram_buffer(13302) := X"10600217";
        ram_buffer(13303) := X"AC430004";
        ram_buffer(13304) := X"8E020014";
        ram_buffer(13305) := X"00000000";
        ram_buffer(13306) := X"8C430000";
        ram_buffer(13307) := X"00000000";
        ram_buffer(13308) := X"24640001";
        ram_buffer(13309) := X"AC440000";
        ram_buffer(13310) := X"A0600000";
        ram_buffer(13311) := X"8C430004";
        ram_buffer(13312) := X"00000000";
        ram_buffer(13313) := X"2463FFFF";
        ram_buffer(13314) := X"106001FD";
        ram_buffer(13315) := X"AC430004";
        ram_buffer(13316) := X"8E020014";
        ram_buffer(13317) := X"00000000";
        ram_buffer(13318) := X"8C430000";
        ram_buffer(13319) := X"00000000";
        ram_buffer(13320) := X"24640001";
        ram_buffer(13321) := X"AC440000";
        ram_buffer(13322) := X"2404000E";
        ram_buffer(13323) := X"A0640000";
        ram_buffer(13324) := X"8C430004";
        ram_buffer(13325) := X"00000000";
        ram_buffer(13326) := X"2463FFFF";
        ram_buffer(13327) := X"106001E2";
        ram_buffer(13328) := X"AC430004";
        ram_buffer(13329) := X"8E020014";
        ram_buffer(13330) := X"00000000";
        ram_buffer(13331) := X"8C430000";
        ram_buffer(13332) := X"00000000";
        ram_buffer(13333) := X"24640001";
        ram_buffer(13334) := X"AC440000";
        ram_buffer(13335) := X"24040041";
        ram_buffer(13336) := X"A0640000";
        ram_buffer(13337) := X"8C430004";
        ram_buffer(13338) := X"00000000";
        ram_buffer(13339) := X"2463FFFF";
        ram_buffer(13340) := X"106001C7";
        ram_buffer(13341) := X"AC430004";
        ram_buffer(13342) := X"8E020014";
        ram_buffer(13343) := X"00000000";
        ram_buffer(13344) := X"8C430000";
        ram_buffer(13345) := X"00000000";
        ram_buffer(13346) := X"24640001";
        ram_buffer(13347) := X"AC440000";
        ram_buffer(13348) := X"24040064";
        ram_buffer(13349) := X"A0640000";
        ram_buffer(13350) := X"8C430004";
        ram_buffer(13351) := X"00000000";
        ram_buffer(13352) := X"2463FFFF";
        ram_buffer(13353) := X"10600254";
        ram_buffer(13354) := X"AC430004";
        ram_buffer(13355) := X"8E020014";
        ram_buffer(13356) := X"00000000";
        ram_buffer(13357) := X"8C430000";
        ram_buffer(13358) := X"00000000";
        ram_buffer(13359) := X"24640001";
        ram_buffer(13360) := X"AC440000";
        ram_buffer(13361) := X"2404006F";
        ram_buffer(13362) := X"A0640000";
        ram_buffer(13363) := X"8C430004";
        ram_buffer(13364) := X"00000000";
        ram_buffer(13365) := X"2463FFFF";
        ram_buffer(13366) := X"10600239";
        ram_buffer(13367) := X"AC430004";
        ram_buffer(13368) := X"8E020014";
        ram_buffer(13369) := X"00000000";
        ram_buffer(13370) := X"8C430000";
        ram_buffer(13371) := X"00000000";
        ram_buffer(13372) := X"24640001";
        ram_buffer(13373) := X"AC440000";
        ram_buffer(13374) := X"24040062";
        ram_buffer(13375) := X"A0640000";
        ram_buffer(13376) := X"8C430004";
        ram_buffer(13377) := X"00000000";
        ram_buffer(13378) := X"2463FFFF";
        ram_buffer(13379) := X"1060021E";
        ram_buffer(13380) := X"AC430004";
        ram_buffer(13381) := X"8E020014";
        ram_buffer(13382) := X"00000000";
        ram_buffer(13383) := X"8C430000";
        ram_buffer(13384) := X"00000000";
        ram_buffer(13385) := X"24640001";
        ram_buffer(13386) := X"AC440000";
        ram_buffer(13387) := X"24040065";
        ram_buffer(13388) := X"A0640000";
        ram_buffer(13389) := X"8C430004";
        ram_buffer(13390) := X"00000000";
        ram_buffer(13391) := X"2463FFFF";
        ram_buffer(13392) := X"10600203";
        ram_buffer(13393) := X"AC430004";
        ram_buffer(13394) := X"8E020014";
        ram_buffer(13395) := X"00000000";
        ram_buffer(13396) := X"8C430000";
        ram_buffer(13397) := X"00000000";
        ram_buffer(13398) := X"24640001";
        ram_buffer(13399) := X"AC440000";
        ram_buffer(13400) := X"A0600000";
        ram_buffer(13401) := X"8C430004";
        ram_buffer(13402) := X"00000000";
        ram_buffer(13403) := X"2463FFFF";
        ram_buffer(13404) := X"106001E9";
        ram_buffer(13405) := X"AC430004";
        ram_buffer(13406) := X"8E020014";
        ram_buffer(13407) := X"00000000";
        ram_buffer(13408) := X"8C430000";
        ram_buffer(13409) := X"00000000";
        ram_buffer(13410) := X"24640001";
        ram_buffer(13411) := X"AC440000";
        ram_buffer(13412) := X"24040064";
        ram_buffer(13413) := X"A0640000";
        ram_buffer(13414) := X"8C430004";
        ram_buffer(13415) := X"00000000";
        ram_buffer(13416) := X"2463FFFF";
        ram_buffer(13417) := X"106001CE";
        ram_buffer(13418) := X"AC430004";
        ram_buffer(13419) := X"8E020014";
        ram_buffer(13420) := X"00000000";
        ram_buffer(13421) := X"8C430000";
        ram_buffer(13422) := X"00000000";
        ram_buffer(13423) := X"24640001";
        ram_buffer(13424) := X"AC440000";
        ram_buffer(13425) := X"A0600000";
        ram_buffer(13426) := X"8C430004";
        ram_buffer(13427) := X"00000000";
        ram_buffer(13428) := X"2463FFFF";
        ram_buffer(13429) := X"106001B4";
        ram_buffer(13430) := X"AC430004";
        ram_buffer(13431) := X"8E020014";
        ram_buffer(13432) := X"00000000";
        ram_buffer(13433) := X"8C430000";
        ram_buffer(13434) := X"00000000";
        ram_buffer(13435) := X"24640001";
        ram_buffer(13436) := X"AC440000";
        ram_buffer(13437) := X"A0600000";
        ram_buffer(13438) := X"8C430004";
        ram_buffer(13439) := X"00000000";
        ram_buffer(13440) := X"2463FFFF";
        ram_buffer(13441) := X"1060019A";
        ram_buffer(13442) := X"AC430004";
        ram_buffer(13443) := X"8E020014";
        ram_buffer(13444) := X"00000000";
        ram_buffer(13445) := X"8C430000";
        ram_buffer(13446) := X"00000000";
        ram_buffer(13447) := X"24640001";
        ram_buffer(13448) := X"AC440000";
        ram_buffer(13449) := X"A0600000";
        ram_buffer(13450) := X"8C430004";
        ram_buffer(13451) := X"00000000";
        ram_buffer(13452) := X"2463FFFF";
        ram_buffer(13453) := X"1060013A";
        ram_buffer(13454) := X"AC430004";
        ram_buffer(13455) := X"8E020014";
        ram_buffer(13456) := X"00000000";
        ram_buffer(13457) := X"8C430000";
        ram_buffer(13458) := X"00000000";
        ram_buffer(13459) := X"24640001";
        ram_buffer(13460) := X"AC440000";
        ram_buffer(13461) := X"A0600000";
        ram_buffer(13462) := X"8C430004";
        ram_buffer(13463) := X"00000000";
        ram_buffer(13464) := X"2463FFFF";
        ram_buffer(13465) := X"10600120";
        ram_buffer(13466) := X"AC430004";
        ram_buffer(13467) := X"8E020038";
        ram_buffer(13468) := X"24030003";
        ram_buffer(13469) := X"104301EE";
        ram_buffer(13470) := X"00000000";
        ram_buffer(13471) := X"24030005";
        ram_buffer(13472) := X"1443001D";
        ram_buffer(13473) := X"00000000";
        ram_buffer(13474) := X"8E020014";
        ram_buffer(13475) := X"00000000";
        ram_buffer(13476) := X"8C430000";
        ram_buffer(13477) := X"00000000";
        ram_buffer(13478) := X"24640001";
        ram_buffer(13479) := X"AC440000";
        ram_buffer(13480) := X"24040002";
        ram_buffer(13481) := X"A0640000";
        ram_buffer(13482) := X"8C430004";
        ram_buffer(13483) := X"00000000";
        ram_buffer(13484) := X"2463FFFF";
        ram_buffer(13485) := X"1460FE13";
        ram_buffer(13486) := X"AC430004";
        ram_buffer(13487) := X"8C42000C";
        ram_buffer(13488) := X"00000000";
        ram_buffer(13489) := X"0040F809";
        ram_buffer(13490) := X"02002021";
        ram_buffer(13491) := X"1440FE0D";
        ram_buffer(13492) := X"24030016";
        ram_buffer(13493) := X"8E020000";
        ram_buffer(13494) := X"8FBF001C";
        ram_buffer(13495) := X"8FB10018";
        ram_buffer(13496) := X"8C590000";
        ram_buffer(13497) := X"02002021";
        ram_buffer(13498) := X"8FB00014";
        ram_buffer(13499) := X"AC430014";
        ram_buffer(13500) := X"03200008";
        ram_buffer(13501) := X"27BD0020";
        ram_buffer(13502) := X"8E020014";
        ram_buffer(13503) := X"00000000";
        ram_buffer(13504) := X"8C430000";
        ram_buffer(13505) := X"00000000";
        ram_buffer(13506) := X"24640001";
        ram_buffer(13507) := X"AC440000";
        ram_buffer(13508) := X"A0600000";
        ram_buffer(13509) := X"8C430004";
        ram_buffer(13510) := X"00000000";
        ram_buffer(13511) := X"2463FFFF";
        ram_buffer(13512) := X"1460FDF8";
        ram_buffer(13513) := X"AC430004";
        ram_buffer(13514) := X"1000FFE4";
        ram_buffer(13515) := X"00000000";
        ram_buffer(13516) := X"8C42000C";
        ram_buffer(13517) := X"00000000";
        ram_buffer(13518) := X"0040F809";
        ram_buffer(13519) := X"02002021";
        ram_buffer(13520) := X"1440FEF3";
        ram_buffer(13521) := X"24040016";
        ram_buffer(13522) := X"8E020000";
        ram_buffer(13523) := X"00000000";
        ram_buffer(13524) := X"8C430000";
        ram_buffer(13525) := X"AC440014";
        ram_buffer(13526) := X"0060F809";
        ram_buffer(13527) := X"02002021";
        ram_buffer(13528) := X"1000FEEB";
        ram_buffer(13529) := X"00000000";
        ram_buffer(13530) := X"8C42000C";
        ram_buffer(13531) := X"00000000";
        ram_buffer(13532) := X"0040F809";
        ram_buffer(13533) := X"02002021";
        ram_buffer(13534) := X"1440FED9";
        ram_buffer(13535) := X"24040016";
        ram_buffer(13536) := X"8E020000";
        ram_buffer(13537) := X"00000000";
        ram_buffer(13538) := X"8C430000";
        ram_buffer(13539) := X"AC440014";
        ram_buffer(13540) := X"0060F809";
        ram_buffer(13541) := X"02002021";
        ram_buffer(13542) := X"1000FED1";
        ram_buffer(13543) := X"00000000";
        ram_buffer(13544) := X"8C42000C";
        ram_buffer(13545) := X"00000000";
        ram_buffer(13546) := X"0040F809";
        ram_buffer(13547) := X"02002021";
        ram_buffer(13548) := X"1440FEBF";
        ram_buffer(13549) := X"24040016";
        ram_buffer(13550) := X"8E020000";
        ram_buffer(13551) := X"00000000";
        ram_buffer(13552) := X"8C430000";
        ram_buffer(13553) := X"AC440014";
        ram_buffer(13554) := X"0060F809";
        ram_buffer(13555) := X"02002021";
        ram_buffer(13556) := X"1000FEB7";
        ram_buffer(13557) := X"00000000";
        ram_buffer(13558) := X"8C42000C";
        ram_buffer(13559) := X"00000000";
        ram_buffer(13560) := X"0040F809";
        ram_buffer(13561) := X"02002021";
        ram_buffer(13562) := X"1440FEA5";
        ram_buffer(13563) := X"24040016";
        ram_buffer(13564) := X"8E020000";
        ram_buffer(13565) := X"00000000";
        ram_buffer(13566) := X"8C430000";
        ram_buffer(13567) := X"AC440014";
        ram_buffer(13568) := X"0060F809";
        ram_buffer(13569) := X"02002021";
        ram_buffer(13570) := X"1000FE9D";
        ram_buffer(13571) := X"00000000";
        ram_buffer(13572) := X"8C42000C";
        ram_buffer(13573) := X"00000000";
        ram_buffer(13574) := X"0040F809";
        ram_buffer(13575) := X"02002021";
        ram_buffer(13576) := X"1440FE8B";
        ram_buffer(13577) := X"24040016";
        ram_buffer(13578) := X"8E020000";
        ram_buffer(13579) := X"00000000";
        ram_buffer(13580) := X"8C430000";
        ram_buffer(13581) := X"AC440014";
        ram_buffer(13582) := X"0060F809";
        ram_buffer(13583) := X"02002021";
        ram_buffer(13584) := X"1000FE83";
        ram_buffer(13585) := X"00000000";
        ram_buffer(13586) := X"8C42000C";
        ram_buffer(13587) := X"00000000";
        ram_buffer(13588) := X"0040F809";
        ram_buffer(13589) := X"02002021";
        ram_buffer(13590) := X"1440FE71";
        ram_buffer(13591) := X"24040016";
        ram_buffer(13592) := X"8E020000";
        ram_buffer(13593) := X"00000000";
        ram_buffer(13594) := X"8C430000";
        ram_buffer(13595) := X"AC440014";
        ram_buffer(13596) := X"0060F809";
        ram_buffer(13597) := X"02002021";
        ram_buffer(13598) := X"1000FE69";
        ram_buffer(13599) := X"00000000";
        ram_buffer(13600) := X"8C42000C";
        ram_buffer(13601) := X"00000000";
        ram_buffer(13602) := X"0040F809";
        ram_buffer(13603) := X"02002021";
        ram_buffer(13604) := X"1440FE57";
        ram_buffer(13605) := X"24040016";
        ram_buffer(13606) := X"8E020000";
        ram_buffer(13607) := X"00000000";
        ram_buffer(13608) := X"8C430000";
        ram_buffer(13609) := X"AC440014";
        ram_buffer(13610) := X"0060F809";
        ram_buffer(13611) := X"02002021";
        ram_buffer(13612) := X"1000FE4F";
        ram_buffer(13613) := X"00000000";
        ram_buffer(13614) := X"8C42000C";
        ram_buffer(13615) := X"00000000";
        ram_buffer(13616) := X"0040F809";
        ram_buffer(13617) := X"02002021";
        ram_buffer(13618) := X"1440FE3C";
        ram_buffer(13619) := X"24040016";
        ram_buffer(13620) := X"8E020000";
        ram_buffer(13621) := X"00000000";
        ram_buffer(13622) := X"8C430000";
        ram_buffer(13623) := X"AC440014";
        ram_buffer(13624) := X"0060F809";
        ram_buffer(13625) := X"02002021";
        ram_buffer(13626) := X"1000FE34";
        ram_buffer(13627) := X"00000000";
        ram_buffer(13628) := X"8C42000C";
        ram_buffer(13629) := X"00000000";
        ram_buffer(13630) := X"0040F809";
        ram_buffer(13631) := X"02002021";
        ram_buffer(13632) := X"1440FE21";
        ram_buffer(13633) := X"24040016";
        ram_buffer(13634) := X"8E020000";
        ram_buffer(13635) := X"00000000";
        ram_buffer(13636) := X"8C430000";
        ram_buffer(13637) := X"AC440014";
        ram_buffer(13638) := X"0060F809";
        ram_buffer(13639) := X"02002021";
        ram_buffer(13640) := X"1000FE19";
        ram_buffer(13641) := X"00000000";
        ram_buffer(13642) := X"8C42000C";
        ram_buffer(13643) := X"00000000";
        ram_buffer(13644) := X"0040F809";
        ram_buffer(13645) := X"02002021";
        ram_buffer(13646) := X"1440FE07";
        ram_buffer(13647) := X"24040016";
        ram_buffer(13648) := X"8E020000";
        ram_buffer(13649) := X"00000000";
        ram_buffer(13650) := X"8C430000";
        ram_buffer(13651) := X"AC440014";
        ram_buffer(13652) := X"0060F809";
        ram_buffer(13653) := X"02002021";
        ram_buffer(13654) := X"1000FDFF";
        ram_buffer(13655) := X"00000000";
        ram_buffer(13656) := X"8C42000C";
        ram_buffer(13657) := X"00000000";
        ram_buffer(13658) := X"0040F809";
        ram_buffer(13659) := X"02002021";
        ram_buffer(13660) := X"1440FDEC";
        ram_buffer(13661) := X"24040016";
        ram_buffer(13662) := X"8E020000";
        ram_buffer(13663) := X"00000000";
        ram_buffer(13664) := X"8C430000";
        ram_buffer(13665) := X"AC440014";
        ram_buffer(13666) := X"0060F809";
        ram_buffer(13667) := X"02002021";
        ram_buffer(13668) := X"1000FDE4";
        ram_buffer(13669) := X"00000000";
        ram_buffer(13670) := X"8C42000C";
        ram_buffer(13671) := X"00000000";
        ram_buffer(13672) := X"0040F809";
        ram_buffer(13673) := X"02002021";
        ram_buffer(13674) := X"1440FDD1";
        ram_buffer(13675) := X"24040016";
        ram_buffer(13676) := X"8E020000";
        ram_buffer(13677) := X"00000000";
        ram_buffer(13678) := X"8C430000";
        ram_buffer(13679) := X"AC440014";
        ram_buffer(13680) := X"0060F809";
        ram_buffer(13681) := X"02002021";
        ram_buffer(13682) := X"1000FDC9";
        ram_buffer(13683) := X"00000000";
        ram_buffer(13684) := X"8C42000C";
        ram_buffer(13685) := X"00000000";
        ram_buffer(13686) := X"0040F809";
        ram_buffer(13687) := X"02002021";
        ram_buffer(13688) := X"1440FDB6";
        ram_buffer(13689) := X"24040016";
        ram_buffer(13690) := X"8E020000";
        ram_buffer(13691) := X"00000000";
        ram_buffer(13692) := X"8C430000";
        ram_buffer(13693) := X"AC440014";
        ram_buffer(13694) := X"0060F809";
        ram_buffer(13695) := X"02002021";
        ram_buffer(13696) := X"1000FDAE";
        ram_buffer(13697) := X"00000000";
        ram_buffer(13698) := X"8C42000C";
        ram_buffer(13699) := X"00000000";
        ram_buffer(13700) := X"0040F809";
        ram_buffer(13701) := X"02002021";
        ram_buffer(13702) := X"1440FD9B";
        ram_buffer(13703) := X"24040016";
        ram_buffer(13704) := X"8E020000";
        ram_buffer(13705) := X"00000000";
        ram_buffer(13706) := X"8C430000";
        ram_buffer(13707) := X"AC440014";
        ram_buffer(13708) := X"0060F809";
        ram_buffer(13709) := X"02002021";
        ram_buffer(13710) := X"1000FD93";
        ram_buffer(13711) := X"00000000";
        ram_buffer(13712) := X"8C42000C";
        ram_buffer(13713) := X"00000000";
        ram_buffer(13714) := X"0040F809";
        ram_buffer(13715) := X"02002021";
        ram_buffer(13716) := X"1440FD80";
        ram_buffer(13717) := X"24040016";
        ram_buffer(13718) := X"8E020000";
        ram_buffer(13719) := X"00000000";
        ram_buffer(13720) := X"8C430000";
        ram_buffer(13721) := X"AC440014";
        ram_buffer(13722) := X"0060F809";
        ram_buffer(13723) := X"02002021";
        ram_buffer(13724) := X"1000FD78";
        ram_buffer(13725) := X"00000000";
        ram_buffer(13726) := X"8C42000C";
        ram_buffer(13727) := X"00000000";
        ram_buffer(13728) := X"0040F809";
        ram_buffer(13729) := X"02002021";
        ram_buffer(13730) := X"1440FD66";
        ram_buffer(13731) := X"24040016";
        ram_buffer(13732) := X"8E020000";
        ram_buffer(13733) := X"00000000";
        ram_buffer(13734) := X"8C430000";
        ram_buffer(13735) := X"AC440014";
        ram_buffer(13736) := X"0060F809";
        ram_buffer(13737) := X"02002021";
        ram_buffer(13738) := X"1000FD5E";
        ram_buffer(13739) := X"00000000";
        ram_buffer(13740) := X"8C42000C";
        ram_buffer(13741) := X"00000000";
        ram_buffer(13742) := X"0040F809";
        ram_buffer(13743) := X"02002021";
        ram_buffer(13744) := X"1440FD4B";
        ram_buffer(13745) := X"24040016";
        ram_buffer(13746) := X"8E020000";
        ram_buffer(13747) := X"00000000";
        ram_buffer(13748) := X"8C430000";
        ram_buffer(13749) := X"AC440014";
        ram_buffer(13750) := X"0060F809";
        ram_buffer(13751) := X"02002021";
        ram_buffer(13752) := X"1000FD43";
        ram_buffer(13753) := X"00000000";
        ram_buffer(13754) := X"8C42000C";
        ram_buffer(13755) := X"00000000";
        ram_buffer(13756) := X"0040F809";
        ram_buffer(13757) := X"02002021";
        ram_buffer(13758) := X"1440FEDC";
        ram_buffer(13759) := X"24040016";
        ram_buffer(13760) := X"8E020000";
        ram_buffer(13761) := X"00000000";
        ram_buffer(13762) := X"8C430000";
        ram_buffer(13763) := X"AC440014";
        ram_buffer(13764) := X"0060F809";
        ram_buffer(13765) := X"02002021";
        ram_buffer(13766) := X"1000FED4";
        ram_buffer(13767) := X"00000000";
        ram_buffer(13768) := X"8C42000C";
        ram_buffer(13769) := X"00000000";
        ram_buffer(13770) := X"0040F809";
        ram_buffer(13771) := X"02002021";
        ram_buffer(13772) := X"1440FEC2";
        ram_buffer(13773) := X"24040016";
        ram_buffer(13774) := X"8E020000";
        ram_buffer(13775) := X"00000000";
        ram_buffer(13776) := X"8C430000";
        ram_buffer(13777) := X"AC440014";
        ram_buffer(13778) := X"0060F809";
        ram_buffer(13779) := X"02002021";
        ram_buffer(13780) := X"1000FEBA";
        ram_buffer(13781) := X"00000000";
        ram_buffer(13782) := X"8C42000C";
        ram_buffer(13783) := X"00000000";
        ram_buffer(13784) := X"0040F809";
        ram_buffer(13785) := X"02002021";
        ram_buffer(13786) := X"1440FE10";
        ram_buffer(13787) := X"24040016";
        ram_buffer(13788) := X"8E020000";
        ram_buffer(13789) := X"00000000";
        ram_buffer(13790) := X"8C430000";
        ram_buffer(13791) := X"AC440014";
        ram_buffer(13792) := X"0060F809";
        ram_buffer(13793) := X"02002021";
        ram_buffer(13794) := X"1000FE08";
        ram_buffer(13795) := X"00000000";
        ram_buffer(13796) := X"8C42000C";
        ram_buffer(13797) := X"00000000";
        ram_buffer(13798) := X"0040F809";
        ram_buffer(13799) := X"02002021";
        ram_buffer(13800) := X"1440FE35";
        ram_buffer(13801) := X"24040016";
        ram_buffer(13802) := X"8E020000";
        ram_buffer(13803) := X"00000000";
        ram_buffer(13804) := X"8C430000";
        ram_buffer(13805) := X"AC440014";
        ram_buffer(13806) := X"0060F809";
        ram_buffer(13807) := X"02002021";
        ram_buffer(13808) := X"1000FE2D";
        ram_buffer(13809) := X"00000000";
        ram_buffer(13810) := X"8C42000C";
        ram_buffer(13811) := X"00000000";
        ram_buffer(13812) := X"0040F809";
        ram_buffer(13813) := X"02002021";
        ram_buffer(13814) := X"1440FE1A";
        ram_buffer(13815) := X"24040016";
        ram_buffer(13816) := X"8E020000";
        ram_buffer(13817) := X"00000000";
        ram_buffer(13818) := X"8C430000";
        ram_buffer(13819) := X"AC440014";
        ram_buffer(13820) := X"0060F809";
        ram_buffer(13821) := X"02002021";
        ram_buffer(13822) := X"1000FE12";
        ram_buffer(13823) := X"00000000";
        ram_buffer(13824) := X"8C42000C";
        ram_buffer(13825) := X"00000000";
        ram_buffer(13826) := X"0040F809";
        ram_buffer(13827) := X"02002021";
        ram_buffer(13828) := X"1440FDFF";
        ram_buffer(13829) := X"24040016";
        ram_buffer(13830) := X"8E020000";
        ram_buffer(13831) := X"00000000";
        ram_buffer(13832) := X"8C430000";
        ram_buffer(13833) := X"AC440014";
        ram_buffer(13834) := X"0060F809";
        ram_buffer(13835) := X"02002021";
        ram_buffer(13836) := X"1000FDF7";
        ram_buffer(13837) := X"00000000";
        ram_buffer(13838) := X"8C42000C";
        ram_buffer(13839) := X"00000000";
        ram_buffer(13840) := X"0040F809";
        ram_buffer(13841) := X"02002021";
        ram_buffer(13842) := X"1440FDE5";
        ram_buffer(13843) := X"24040016";
        ram_buffer(13844) := X"8E020000";
        ram_buffer(13845) := X"00000000";
        ram_buffer(13846) := X"8C430000";
        ram_buffer(13847) := X"AC440014";
        ram_buffer(13848) := X"0060F809";
        ram_buffer(13849) := X"02002021";
        ram_buffer(13850) := X"1000FDDD";
        ram_buffer(13851) := X"00000000";
        ram_buffer(13852) := X"8C42000C";
        ram_buffer(13853) := X"00000000";
        ram_buffer(13854) := X"0040F809";
        ram_buffer(13855) := X"02002021";
        ram_buffer(13856) := X"1440FE62";
        ram_buffer(13857) := X"24040016";
        ram_buffer(13858) := X"8E020000";
        ram_buffer(13859) := X"00000000";
        ram_buffer(13860) := X"8C430000";
        ram_buffer(13861) := X"AC440014";
        ram_buffer(13862) := X"0060F809";
        ram_buffer(13863) := X"02002021";
        ram_buffer(13864) := X"1000FE5A";
        ram_buffer(13865) := X"00000000";
        ram_buffer(13866) := X"8C42000C";
        ram_buffer(13867) := X"00000000";
        ram_buffer(13868) := X"0040F809";
        ram_buffer(13869) := X"02002021";
        ram_buffer(13870) := X"1440FE48";
        ram_buffer(13871) := X"24040016";
        ram_buffer(13872) := X"8E020000";
        ram_buffer(13873) := X"00000000";
        ram_buffer(13874) := X"8C430000";
        ram_buffer(13875) := X"AC440014";
        ram_buffer(13876) := X"0060F809";
        ram_buffer(13877) := X"02002021";
        ram_buffer(13878) := X"1000FE40";
        ram_buffer(13879) := X"00000000";
        ram_buffer(13880) := X"8C42000C";
        ram_buffer(13881) := X"00000000";
        ram_buffer(13882) := X"0040F809";
        ram_buffer(13883) := X"02002021";
        ram_buffer(13884) := X"1440FE2E";
        ram_buffer(13885) := X"24040016";
        ram_buffer(13886) := X"8E020000";
        ram_buffer(13887) := X"00000000";
        ram_buffer(13888) := X"8C430000";
        ram_buffer(13889) := X"AC440014";
        ram_buffer(13890) := X"0060F809";
        ram_buffer(13891) := X"02002021";
        ram_buffer(13892) := X"1000FE26";
        ram_buffer(13893) := X"00000000";
        ram_buffer(13894) := X"8C42000C";
        ram_buffer(13895) := X"00000000";
        ram_buffer(13896) := X"0040F809";
        ram_buffer(13897) := X"02002021";
        ram_buffer(13898) := X"1440FE13";
        ram_buffer(13899) := X"24040016";
        ram_buffer(13900) := X"8E020000";
        ram_buffer(13901) := X"00000000";
        ram_buffer(13902) := X"8C430000";
        ram_buffer(13903) := X"AC440014";
        ram_buffer(13904) := X"0060F809";
        ram_buffer(13905) := X"02002021";
        ram_buffer(13906) := X"1000FE0B";
        ram_buffer(13907) := X"00000000";
        ram_buffer(13908) := X"8C42000C";
        ram_buffer(13909) := X"00000000";
        ram_buffer(13910) := X"0040F809";
        ram_buffer(13911) := X"02002021";
        ram_buffer(13912) := X"1440FDF9";
        ram_buffer(13913) := X"24040016";
        ram_buffer(13914) := X"8E020000";
        ram_buffer(13915) := X"00000000";
        ram_buffer(13916) := X"8C430000";
        ram_buffer(13917) := X"AC440014";
        ram_buffer(13918) := X"0060F809";
        ram_buffer(13919) := X"02002021";
        ram_buffer(13920) := X"1000FDF1";
        ram_buffer(13921) := X"00000000";
        ram_buffer(13922) := X"8C42000C";
        ram_buffer(13923) := X"00000000";
        ram_buffer(13924) := X"0040F809";
        ram_buffer(13925) := X"02002021";
        ram_buffer(13926) := X"1440FDDE";
        ram_buffer(13927) := X"24040016";
        ram_buffer(13928) := X"8E020000";
        ram_buffer(13929) := X"00000000";
        ram_buffer(13930) := X"8C430000";
        ram_buffer(13931) := X"AC440014";
        ram_buffer(13932) := X"0060F809";
        ram_buffer(13933) := X"02002021";
        ram_buffer(13934) := X"1000FDD6";
        ram_buffer(13935) := X"00000000";
        ram_buffer(13936) := X"8C42000C";
        ram_buffer(13937) := X"00000000";
        ram_buffer(13938) := X"0040F809";
        ram_buffer(13939) := X"02002021";
        ram_buffer(13940) := X"1440FDC3";
        ram_buffer(13941) := X"24040016";
        ram_buffer(13942) := X"8E020000";
        ram_buffer(13943) := X"00000000";
        ram_buffer(13944) := X"8C430000";
        ram_buffer(13945) := X"AC440014";
        ram_buffer(13946) := X"0060F809";
        ram_buffer(13947) := X"02002021";
        ram_buffer(13948) := X"1000FDBB";
        ram_buffer(13949) := X"00000000";
        ram_buffer(13950) := X"8C42000C";
        ram_buffer(13951) := X"00000000";
        ram_buffer(13952) := X"0040F809";
        ram_buffer(13953) := X"02002021";
        ram_buffer(13954) := X"1440FDA8";
        ram_buffer(13955) := X"24040016";
        ram_buffer(13956) := X"8E020000";
        ram_buffer(13957) := X"00000000";
        ram_buffer(13958) := X"8C430000";
        ram_buffer(13959) := X"AC440014";
        ram_buffer(13960) := X"0060F809";
        ram_buffer(13961) := X"02002021";
        ram_buffer(13962) := X"1000FDA0";
        ram_buffer(13963) := X"00000000";
        ram_buffer(13964) := X"8E020014";
        ram_buffer(13965) := X"00000000";
        ram_buffer(13966) := X"8C430000";
        ram_buffer(13967) := X"00000000";
        ram_buffer(13968) := X"24640001";
        ram_buffer(13969) := X"AC440000";
        ram_buffer(13970) := X"1000FE16";
        ram_buffer(13971) := X"24040001";
        ram_buffer(13972) := X"8C820004";
        ram_buffer(13973) := X"27BDFFE8";
        ram_buffer(13974) := X"8C420000";
        ram_buffer(13975) := X"24060018";
        ram_buffer(13976) := X"AFBF0014";
        ram_buffer(13977) := X"AFB00010";
        ram_buffer(13978) := X"24050001";
        ram_buffer(13979) := X"0040F809";
        ram_buffer(13980) := X"00808021";
        ram_buffer(13981) := X"3C031009";
        ram_buffer(13982) := X"2463A62C";
        ram_buffer(13983) := X"AE020154";
        ram_buffer(13984) := X"AC430000";
        ram_buffer(13985) := X"3C031009";
        ram_buffer(13986) := X"2463CA74";
        ram_buffer(13987) := X"AC430004";
        ram_buffer(13988) := X"3C031009";
        ram_buffer(13989) := X"2463C604";
        ram_buffer(13990) := X"AC430008";
        ram_buffer(13991) := X"3C031009";
        ram_buffer(13992) := X"2463B440";
        ram_buffer(13993) := X"AC43000C";
        ram_buffer(13994) := X"3C031009";
        ram_buffer(13995) := X"2463A514";
        ram_buffer(13996) := X"AC430010";
        ram_buffer(13997) := X"8FBF0014";
        ram_buffer(13998) := X"3C031009";
        ram_buffer(13999) := X"2463C7D0";
        ram_buffer(14000) := X"8FB00010";
        ram_buffer(14001) := X"AC430014";
        ram_buffer(14002) := X"03E00008";
        ram_buffer(14003) := X"27BD0018";
        ram_buffer(14004) := X"27BDFFB8";
        ram_buffer(14005) := X"AFB00024";
        ram_buffer(14006) := X"8C900148";
        ram_buffer(14007) := X"8C8300E8";
        ram_buffer(14008) := X"8E020008";
        ram_buffer(14009) := X"AFBF0044";
        ram_buffer(14010) := X"0043102B";
        ram_buffer(14011) := X"AFB70040";
        ram_buffer(14012) := X"AFB6003C";
        ram_buffer(14013) := X"AFB50038";
        ram_buffer(14014) := X"AFB40034";
        ram_buffer(14015) := X"AFB30030";
        ram_buffer(14016) := X"AFB2002C";
        ram_buffer(14017) := X"10400033";
        ram_buffer(14018) := X"AFB10028";
        ram_buffer(14019) := X"8E02000C";
        ram_buffer(14020) := X"00E0A821";
        ram_buffer(14021) := X"2C430008";
        ram_buffer(14022) := X"00C08821";
        ram_buffer(14023) := X"00A0A021";
        ram_buffer(14024) := X"0080B821";
        ram_buffer(14025) := X"24120008";
        ram_buffer(14026) := X"2616000C";
        ram_buffer(14027) := X"1460001B";
        ram_buffer(14028) := X"26130018";
        ram_buffer(14029) := X"14520027";
        ram_buffer(14030) := X"00000000";
        ram_buffer(14031) := X"8EE20150";
        ram_buffer(14032) := X"02602821";
        ram_buffer(14033) := X"8C420004";
        ram_buffer(14034) := X"00000000";
        ram_buffer(14035) := X"0040F809";
        ram_buffer(14036) := X"02E02021";
        ram_buffer(14037) := X"1040002A";
        ram_buffer(14038) := X"00000000";
        ram_buffer(14039) := X"8E020010";
        ram_buffer(14040) := X"00000000";
        ram_buffer(14041) := X"10400006";
        ram_buffer(14042) := X"00000000";
        ram_buffer(14043) := X"8E220000";
        ram_buffer(14044) := X"00000000";
        ram_buffer(14045) := X"24420001";
        ram_buffer(14046) := X"AE220000";
        ram_buffer(14047) := X"AE000010";
        ram_buffer(14048) := X"8E020008";
        ram_buffer(14049) := X"8EE300E8";
        ram_buffer(14050) := X"24420001";
        ram_buffer(14051) := X"0043182B";
        ram_buffer(14052) := X"AE00000C";
        ram_buffer(14053) := X"1060000F";
        ram_buffer(14054) := X"AE020008";
        ram_buffer(14055) := X"8EE2014C";
        ram_buffer(14056) := X"AFB20018";
        ram_buffer(14057) := X"AFB60014";
        ram_buffer(14058) := X"AFB30010";
        ram_buffer(14059) := X"8C420004";
        ram_buffer(14060) := X"02A03821";
        ram_buffer(14061) := X"02203021";
        ram_buffer(14062) := X"02802821";
        ram_buffer(14063) := X"0040F809";
        ram_buffer(14064) := X"02E02021";
        ram_buffer(14065) := X"8E02000C";
        ram_buffer(14066) := X"00000000";
        ram_buffer(14067) := X"1052FFDB";
        ram_buffer(14068) := X"00000000";
        ram_buffer(14069) := X"8FBF0044";
        ram_buffer(14070) := X"8FB70040";
        ram_buffer(14071) := X"8FB6003C";
        ram_buffer(14072) := X"8FB50038";
        ram_buffer(14073) := X"8FB40034";
        ram_buffer(14074) := X"8FB30030";
        ram_buffer(14075) := X"8FB2002C";
        ram_buffer(14076) := X"8FB10028";
        ram_buffer(14077) := X"8FB00024";
        ram_buffer(14078) := X"03E00008";
        ram_buffer(14079) := X"27BD0048";
        ram_buffer(14080) := X"8E020010";
        ram_buffer(14081) := X"00000000";
        ram_buffer(14082) := X"1440FFF2";
        ram_buffer(14083) := X"00000000";
        ram_buffer(14084) := X"8E220000";
        ram_buffer(14085) := X"00000000";
        ram_buffer(14086) := X"2442FFFF";
        ram_buffer(14087) := X"AE220000";
        ram_buffer(14088) := X"24020001";
        ram_buffer(14089) := X"1000FFEB";
        ram_buffer(14090) := X"AE020010";
        ram_buffer(14091) := X"8C8200A8";
        ram_buffer(14092) := X"00000000";
        ram_buffer(14093) := X"1440000C";
        ram_buffer(14094) := X"00000000";
        ram_buffer(14095) := X"8C820148";
        ram_buffer(14096) := X"00000000";
        ram_buffer(14097) := X"AC400008";
        ram_buffer(14098) := X"AC40000C";
        ram_buffer(14099) := X"AC400010";
        ram_buffer(14100) := X"14A00007";
        ram_buffer(14101) := X"AC450014";
        ram_buffer(14102) := X"3C031009";
        ram_buffer(14103) := X"2463DAD0";
        ram_buffer(14104) := X"03E00008";
        ram_buffer(14105) := X"AC430004";
        ram_buffer(14106) := X"03E00008";
        ram_buffer(14107) := X"00000000";
        ram_buffer(14108) := X"8C820000";
        ram_buffer(14109) := X"24030004";
        ram_buffer(14110) := X"8C590000";
        ram_buffer(14111) := X"00000000";
        ram_buffer(14112) := X"03200008";
        ram_buffer(14113) := X"AC430014";
        ram_buffer(14114) := X"8C820004";
        ram_buffer(14115) := X"27BDFFD8";
        ram_buffer(14116) := X"8C420000";
        ram_buffer(14117) := X"24060040";
        ram_buffer(14118) := X"AFB10018";
        ram_buffer(14119) := X"AFB00014";
        ram_buffer(14120) := X"00808821";
        ram_buffer(14121) := X"AFBF0024";
        ram_buffer(14122) := X"AFB30020";
        ram_buffer(14123) := X"AFB2001C";
        ram_buffer(14124) := X"00A08021";
        ram_buffer(14125) := X"0040F809";
        ram_buffer(14126) := X"24050001";
        ram_buffer(14127) := X"8E2400A8";
        ram_buffer(14128) := X"3C031009";
        ram_buffer(14129) := X"2463DC2C";
        ram_buffer(14130) := X"AE220148";
        ram_buffer(14131) := X"14800018";
        ram_buffer(14132) := X"AC430000";
        ram_buffer(14133) := X"1600001D";
        ram_buffer(14134) := X"24030004";
        ram_buffer(14135) := X"8E230034";
        ram_buffer(14136) := X"8E30003C";
        ram_buffer(14137) := X"18600012";
        ram_buffer(14138) := X"24520018";
        ram_buffer(14139) := X"00009821";
        ram_buffer(14140) := X"8E220004";
        ram_buffer(14141) := X"8E07000C";
        ram_buffer(14142) := X"8E06001C";
        ram_buffer(14143) := X"8C420008";
        ram_buffer(14144) := X"000738C0";
        ram_buffer(14145) := X"000630C0";
        ram_buffer(14146) := X"24050001";
        ram_buffer(14147) := X"0040F809";
        ram_buffer(14148) := X"02202021";
        ram_buffer(14149) := X"8E230034";
        ram_buffer(14150) := X"26730001";
        ram_buffer(14151) := X"0263182A";
        ram_buffer(14152) := X"AE420000";
        ram_buffer(14153) := X"26100054";
        ram_buffer(14154) := X"1460FFF1";
        ram_buffer(14155) := X"26520004";
        ram_buffer(14156) := X"8FBF0024";
        ram_buffer(14157) := X"8FB30020";
        ram_buffer(14158) := X"8FB2001C";
        ram_buffer(14159) := X"8FB10018";
        ram_buffer(14160) := X"8FB00014";
        ram_buffer(14161) := X"03E00008";
        ram_buffer(14162) := X"27BD0028";
        ram_buffer(14163) := X"8E220000";
        ram_buffer(14164) := X"8FBF0024";
        ram_buffer(14165) := X"8FB30020";
        ram_buffer(14166) := X"8FB2001C";
        ram_buffer(14167) := X"8FB00014";
        ram_buffer(14168) := X"8C590000";
        ram_buffer(14169) := X"02202021";
        ram_buffer(14170) := X"8FB10018";
        ram_buffer(14171) := X"AC430014";
        ram_buffer(14172) := X"03200008";
        ram_buffer(14173) := X"27BD0028";
        ram_buffer(14174) := X"27BDFFE0";
        ram_buffer(14175) := X"AFB10018";
        ram_buffer(14176) := X"AFB00014";
        ram_buffer(14177) := X"AFBF001C";
        ram_buffer(14178) := X"8C90014C";
        ram_buffer(14179) := X"10A00007";
        ram_buffer(14180) := X"00808821";
        ram_buffer(14181) := X"8C820000";
        ram_buffer(14182) := X"24050004";
        ram_buffer(14183) := X"8C430000";
        ram_buffer(14184) := X"00000000";
        ram_buffer(14185) := X"0060F809";
        ram_buffer(14186) := X"AC450014";
        ram_buffer(14187) := X"8E2200E4";
        ram_buffer(14188) := X"8E23001C";
        ram_buffer(14189) := X"8FBF001C";
        ram_buffer(14190) := X"00021040";
        ram_buffer(14191) := X"AE030030";
        ram_buffer(14192) := X"AE000034";
        ram_buffer(14193) := X"AE000038";
        ram_buffer(14194) := X"AE02003C";
        ram_buffer(14195) := X"8FB10018";
        ram_buffer(14196) := X"8FB00014";
        ram_buffer(14197) := X"03E00008";
        ram_buffer(14198) := X"27BD0020";
        ram_buffer(14199) := X"27BDFFB8";
        ram_buffer(14200) := X"AFB50034";
        ram_buffer(14201) := X"8C95014C";
        ram_buffer(14202) := X"AFB40030";
        ram_buffer(14203) := X"26A20008";
        ram_buffer(14204) := X"AFB3002C";
        ram_buffer(14205) := X"AFBF0044";
        ram_buffer(14206) := X"AFBE0040";
        ram_buffer(14207) := X"AFB7003C";
        ram_buffer(14208) := X"AFB60038";
        ram_buffer(14209) := X"AFB20028";
        ram_buffer(14210) := X"AFB10024";
        ram_buffer(14211) := X"AFB00020";
        ram_buffer(14212) := X"0080A021";
        ram_buffer(14213) := X"AFA5004C";
        ram_buffer(14214) := X"AFA60050";
        ram_buffer(14215) := X"AFA70054";
        ram_buffer(14216) := X"AFA2001C";
        ram_buffer(14217) := X"24130001";
        ram_buffer(14218) := X"8FA20050";
        ram_buffer(14219) := X"00000000";
        ram_buffer(14220) := X"8C450000";
        ram_buffer(14221) := X"8FA20054";
        ram_buffer(14222) := X"00000000";
        ram_buffer(14223) := X"00A2102B";
        ram_buffer(14224) := X"10400059";
        ram_buffer(14225) := X"00000000";
        ram_buffer(14226) := X"8FA2005C";
        ram_buffer(14227) := X"8FA30060";
        ram_buffer(14228) := X"8C420000";
        ram_buffer(14229) := X"00000000";
        ram_buffer(14230) := X"0043102B";
        ram_buffer(14231) := X"10400052";
        ram_buffer(14232) := X"00000000";
        ram_buffer(14233) := X"8EA70034";
        ram_buffer(14234) := X"8E9000E4";
        ram_buffer(14235) := X"8FA20054";
        ram_buffer(14236) := X"02078023";
        ram_buffer(14237) := X"00451023";
        ram_buffer(14238) := X"0050182B";
        ram_buffer(14239) := X"10600002";
        ram_buffer(14240) := X"00000000";
        ram_buffer(14241) := X"00408021";
        ram_buffer(14242) := X"8E820158";
        ram_buffer(14243) := X"8FA3004C";
        ram_buffer(14244) := X"AFB00010";
        ram_buffer(14245) := X"8FB7001C";
        ram_buffer(14246) := X"8C420004";
        ram_buffer(14247) := X"00052880";
        ram_buffer(14248) := X"00652821";
        ram_buffer(14249) := X"02E03021";
        ram_buffer(14250) := X"0040F809";
        ram_buffer(14251) := X"02802021";
        ram_buffer(14252) := X"8FA20050";
        ram_buffer(14253) := X"8FA30050";
        ram_buffer(14254) := X"8C420000";
        ram_buffer(14255) := X"00000000";
        ram_buffer(14256) := X"00501021";
        ram_buffer(14257) := X"AC620000";
        ram_buffer(14258) := X"8EA20034";
        ram_buffer(14259) := X"8EA30030";
        ram_buffer(14260) := X"02021021";
        ram_buffer(14261) := X"00708023";
        ram_buffer(14262) := X"AEA20034";
        ram_buffer(14263) := X"16000026";
        ram_buffer(14264) := X"AEB00030";
        ram_buffer(14265) := X"8E9000E4";
        ram_buffer(14266) := X"00000000";
        ram_buffer(14267) := X"0050182A";
        ram_buffer(14268) := X"10600082";
        ram_buffer(14269) := X"00000000";
        ram_buffer(14270) := X"8E850034";
        ram_buffer(14271) := X"00000000";
        ram_buffer(14272) := X"18A00035";
        ram_buffer(14273) := X"0040F021";
        ram_buffer(14274) := X"AFA00018";
        ram_buffer(14275) := X"03D0202A";
        ram_buffer(14276) := X"8EF60000";
        ram_buffer(14277) := X"8E910018";
        ram_buffer(14278) := X"1080000D";
        ram_buffer(14279) := X"03C03821";
        ram_buffer(14280) := X"27D2FFFF";
        ram_buffer(14281) := X"AFB10014";
        ram_buffer(14282) := X"27DE0001";
        ram_buffer(14283) := X"AFB30010";
        ram_buffer(14284) := X"02C03021";
        ram_buffer(14285) := X"02402821";
        ram_buffer(14286) := X"0C0264BB";
        ram_buffer(14287) := X"02C02021";
        ram_buffer(14288) := X"17D0FFF8";
        ram_buffer(14289) := X"03C03821";
        ram_buffer(14290) := X"8E9000E4";
        ram_buffer(14291) := X"8E850034";
        ram_buffer(14292) := X"8FA20018";
        ram_buffer(14293) := X"00000000";
        ram_buffer(14294) := X"24420001";
        ram_buffer(14295) := X"AFA20018";
        ram_buffer(14296) := X"0045102A";
        ram_buffer(14297) := X"1040001C";
        ram_buffer(14298) := X"26F70004";
        ram_buffer(14299) := X"8EBE0034";
        ram_buffer(14300) := X"1000FFE7";
        ram_buffer(14301) := X"03D0202A";
        ram_buffer(14302) := X"8E8300E4";
        ram_buffer(14303) := X"00000000";
        ram_buffer(14304) := X"10430016";
        ram_buffer(14305) := X"00000000";
        ram_buffer(14306) := X"8FA20050";
        ram_buffer(14307) := X"00000000";
        ram_buffer(14308) := X"8C450000";
        ram_buffer(14309) := X"8FA20054";
        ram_buffer(14310) := X"00000000";
        ram_buffer(14311) := X"00A2102B";
        ram_buffer(14312) := X"1440FFA9";
        ram_buffer(14313) := X"00000000";
        ram_buffer(14314) := X"8FBF0044";
        ram_buffer(14315) := X"8FBE0040";
        ram_buffer(14316) := X"8FB7003C";
        ram_buffer(14317) := X"8FB60038";
        ram_buffer(14318) := X"8FB50034";
        ram_buffer(14319) := X"8FB40030";
        ram_buffer(14320) := X"8FB3002C";
        ram_buffer(14321) := X"8FB20028";
        ram_buffer(14322) := X"8FB10024";
        ram_buffer(14323) := X"8FB00020";
        ram_buffer(14324) := X"03E00008";
        ram_buffer(14325) := X"27BD0048";
        ram_buffer(14326) := X"AEB00034";
        ram_buffer(14327) := X"8FA2005C";
        ram_buffer(14328) := X"8FA70058";
        ram_buffer(14329) := X"8C430000";
        ram_buffer(14330) := X"8E82015C";
        ram_buffer(14331) := X"AFA30010";
        ram_buffer(14332) := X"8C420004";
        ram_buffer(14333) := X"8FA5001C";
        ram_buffer(14334) := X"00003021";
        ram_buffer(14335) := X"0040F809";
        ram_buffer(14336) := X"02802021";
        ram_buffer(14337) := X"8FA2005C";
        ram_buffer(14338) := X"AEA00034";
        ram_buffer(14339) := X"8C420000";
        ram_buffer(14340) := X"8FA3005C";
        ram_buffer(14341) := X"24420001";
        ram_buffer(14342) := X"AC620000";
        ram_buffer(14343) := X"8EA30030";
        ram_buffer(14344) := X"00000000";
        ram_buffer(14345) := X"1460FF80";
        ram_buffer(14346) := X"00000000";
        ram_buffer(14347) := X"8FA30060";
        ram_buffer(14348) := X"00000000";
        ram_buffer(14349) := X"0043182B";
        ram_buffer(14350) := X"1060FF7B";
        ram_buffer(14351) := X"00000000";
        ram_buffer(14352) := X"8E830034";
        ram_buffer(14353) := X"8E96003C";
        ram_buffer(14354) := X"18600033";
        ram_buffer(14355) := X"0000B821";
        ram_buffer(14356) := X"8FA40058";
        ram_buffer(14357) := X"00000000";
        ram_buffer(14358) := X"AFA40018";
        ram_buffer(14359) := X"24130001";
        ram_buffer(14360) := X"8ED0000C";
        ram_buffer(14361) := X"8ED1001C";
        ram_buffer(14362) := X"02020018";
        ram_buffer(14363) := X"8FA20018";
        ram_buffer(14364) := X"00000000";
        ram_buffer(14365) := X"8C550000";
        ram_buffer(14366) := X"8FA20060";
        ram_buffer(14367) := X"0000F012";
        ram_buffer(14368) := X"00000000";
        ram_buffer(14369) := X"00000000";
        ram_buffer(14370) := X"00500018";
        ram_buffer(14371) := X"00008012";
        ram_buffer(14372) := X"03D0202A";
        ram_buffer(14373) := X"1080000D";
        ram_buffer(14374) := X"001188C0";
        ram_buffer(14375) := X"27D2FFFF";
        ram_buffer(14376) := X"03C03821";
        ram_buffer(14377) := X"AFB10014";
        ram_buffer(14378) := X"27DE0001";
        ram_buffer(14379) := X"AFB30010";
        ram_buffer(14380) := X"02A03021";
        ram_buffer(14381) := X"02402821";
        ram_buffer(14382) := X"0C0264BB";
        ram_buffer(14383) := X"02A02021";
        ram_buffer(14384) := X"161EFFF8";
        ram_buffer(14385) := X"03C03821";
        ram_buffer(14386) := X"8E830034";
        ram_buffer(14387) := X"8FA40018";
        ram_buffer(14388) := X"26F70001";
        ram_buffer(14389) := X"24840004";
        ram_buffer(14390) := X"02E3102A";
        ram_buffer(14391) := X"26D60054";
        ram_buffer(14392) := X"1040000D";
        ram_buffer(14393) := X"AFA40018";
        ram_buffer(14394) := X"8FA2005C";
        ram_buffer(14395) := X"00000000";
        ram_buffer(14396) := X"8C420000";
        ram_buffer(14397) := X"1000FFDA";
        ram_buffer(14398) := X"00000000";
        ram_buffer(14399) := X"1050FFB7";
        ram_buffer(14400) := X"00000000";
        ram_buffer(14401) := X"8FA2005C";
        ram_buffer(14402) := X"00000000";
        ram_buffer(14403) := X"8C420000";
        ram_buffer(14404) := X"1000FFC6";
        ram_buffer(14405) := X"00000000";
        ram_buffer(14406) := X"8FA2005C";
        ram_buffer(14407) := X"8FA30060";
        ram_buffer(14408) := X"1000FFA1";
        ram_buffer(14409) := X"AC430000";
        ram_buffer(14410) := X"8C8200E4";
        ram_buffer(14411) := X"27BDFFB0";
        ram_buffer(14412) := X"00021840";
        ram_buffer(14413) := X"AFB5003C";
        ram_buffer(14414) := X"8C95014C";
        ram_buffer(14415) := X"00621021";
        ram_buffer(14416) := X"AFA20020";
        ram_buffer(14417) := X"26A20008";
        ram_buffer(14418) := X"AFB40038";
        ram_buffer(14419) := X"AFB1002C";
        ram_buffer(14420) := X"AFBF004C";
        ram_buffer(14421) := X"AFBE0048";
        ram_buffer(14422) := X"AFB70044";
        ram_buffer(14423) := X"AFB60040";
        ram_buffer(14424) := X"AFB30034";
        ram_buffer(14425) := X"AFB20030";
        ram_buffer(14426) := X"AFB00028";
        ram_buffer(14427) := X"0080A021";
        ram_buffer(14428) := X"AFA50054";
        ram_buffer(14429) := X"AFA60058";
        ram_buffer(14430) := X"AFA7005C";
        ram_buffer(14431) := X"AFA2001C";
        ram_buffer(14432) := X"24110001";
        ram_buffer(14433) := X"8FA20064";
        ram_buffer(14434) := X"00000000";
        ram_buffer(14435) := X"8C440000";
        ram_buffer(14436) := X"8FA20068";
        ram_buffer(14437) := X"00000000";
        ram_buffer(14438) := X"0082102B";
        ram_buffer(14439) := X"10400060";
        ram_buffer(14440) := X"00000000";
        ram_buffer(14441) := X"8FA20058";
        ram_buffer(14442) := X"8FA3005C";
        ram_buffer(14443) := X"8C420000";
        ram_buffer(14444) := X"00000000";
        ram_buffer(14445) := X"0043182B";
        ram_buffer(14446) := X"1460002C";
        ram_buffer(14447) := X"00000000";
        ram_buffer(14448) := X"8EA20030";
        ram_buffer(14449) := X"00000000";
        ram_buffer(14450) := X"14400055";
        ram_buffer(14451) := X"00000000";
        ram_buffer(14452) := X"8EA20034";
        ram_buffer(14453) := X"8EB0003C";
        ram_buffer(14454) := X"00000000";
        ram_buffer(14455) := X"0050182A";
        ram_buffer(14456) := X"10600048";
        ram_buffer(14457) := X"00000000";
        ram_buffer(14458) := X"8E850034";
        ram_buffer(14459) := X"00000000";
        ram_buffer(14460) := X"18A00057";
        ram_buffer(14461) := X"0040F021";
        ram_buffer(14462) := X"8FB7001C";
        ram_buffer(14463) := X"AFA00018";
        ram_buffer(14464) := X"03D0202A";
        ram_buffer(14465) := X"8EF60000";
        ram_buffer(14466) := X"8E920018";
        ram_buffer(14467) := X"1080000D";
        ram_buffer(14468) := X"03C03821";
        ram_buffer(14469) := X"27D3FFFF";
        ram_buffer(14470) := X"AFB20014";
        ram_buffer(14471) := X"27DE0001";
        ram_buffer(14472) := X"AFB10010";
        ram_buffer(14473) := X"02C03021";
        ram_buffer(14474) := X"02602821";
        ram_buffer(14475) := X"0C0264BB";
        ram_buffer(14476) := X"02C02021";
        ram_buffer(14477) := X"17D0FFF8";
        ram_buffer(14478) := X"03C03821";
        ram_buffer(14479) := X"8EB0003C";
        ram_buffer(14480) := X"8E850034";
        ram_buffer(14481) := X"8FA20018";
        ram_buffer(14482) := X"00000000";
        ram_buffer(14483) := X"24420001";
        ram_buffer(14484) := X"AFA20018";
        ram_buffer(14485) := X"0045102A";
        ram_buffer(14486) := X"1040003D";
        ram_buffer(14487) := X"26F70004";
        ram_buffer(14488) := X"8EBE0034";
        ram_buffer(14489) := X"1000FFE7";
        ram_buffer(14490) := X"03D0202A";
        ram_buffer(14491) := X"8EA70034";
        ram_buffer(14492) := X"8EB3003C";
        ram_buffer(14493) := X"8FA3005C";
        ram_buffer(14494) := X"02679823";
        ram_buffer(14495) := X"00621823";
        ram_buffer(14496) := X"0073202B";
        ram_buffer(14497) := X"10800002";
        ram_buffer(14498) := X"00000000";
        ram_buffer(14499) := X"00609821";
        ram_buffer(14500) := X"8E830158";
        ram_buffer(14501) := X"00022880";
        ram_buffer(14502) := X"AFB30010";
        ram_buffer(14503) := X"8FA20054";
        ram_buffer(14504) := X"8C630004";
        ram_buffer(14505) := X"8FA6001C";
        ram_buffer(14506) := X"00452821";
        ram_buffer(14507) := X"0060F809";
        ram_buffer(14508) := X"02802021";
        ram_buffer(14509) := X"8EA30030";
        ram_buffer(14510) := X"8E82001C";
        ram_buffer(14511) := X"00000000";
        ram_buffer(14512) := X"10620047";
        ram_buffer(14513) := X"00000000";
        ram_buffer(14514) := X"8FA20058";
        ram_buffer(14515) := X"8FA30058";
        ram_buffer(14516) := X"8C420000";
        ram_buffer(14517) := X"00000000";
        ram_buffer(14518) := X"00531021";
        ram_buffer(14519) := X"AC620000";
        ram_buffer(14520) := X"8EA30030";
        ram_buffer(14521) := X"8EA20034";
        ram_buffer(14522) := X"8EB0003C";
        ram_buffer(14523) := X"02621021";
        ram_buffer(14524) := X"00739823";
        ram_buffer(14525) := X"8FA30064";
        ram_buffer(14526) := X"AEA20034";
        ram_buffer(14527) := X"AEB30030";
        ram_buffer(14528) := X"8C640000";
        ram_buffer(14529) := X"10500015";
        ram_buffer(14530) := X"00000000";
        ram_buffer(14531) := X"8FA20068";
        ram_buffer(14532) := X"00000000";
        ram_buffer(14533) := X"0082102B";
        ram_buffer(14534) := X"1440FFA2";
        ram_buffer(14535) := X"00000000";
        ram_buffer(14536) := X"8FBF004C";
        ram_buffer(14537) := X"8FBE0048";
        ram_buffer(14538) := X"8FB70044";
        ram_buffer(14539) := X"8FB60040";
        ram_buffer(14540) := X"8FB5003C";
        ram_buffer(14541) := X"8FB40038";
        ram_buffer(14542) := X"8FB30034";
        ram_buffer(14543) := X"8FB20030";
        ram_buffer(14544) := X"8FB1002C";
        ram_buffer(14545) := X"8FB00028";
        ram_buffer(14546) := X"03E00008";
        ram_buffer(14547) := X"27BD0050";
        ram_buffer(14548) := X"8FA20064";
        ram_buffer(14549) := X"AEB00034";
        ram_buffer(14550) := X"8C440000";
        ram_buffer(14551) := X"8E82015C";
        ram_buffer(14552) := X"8EA60038";
        ram_buffer(14553) := X"AFA40010";
        ram_buffer(14554) := X"8C420004";
        ram_buffer(14555) := X"8FA70060";
        ram_buffer(14556) := X"8FA5001C";
        ram_buffer(14557) := X"0040F809";
        ram_buffer(14558) := X"02802021";
        ram_buffer(14559) := X"8FA20064";
        ram_buffer(14560) := X"8FA30064";
        ram_buffer(14561) := X"8C420000";
        ram_buffer(14562) := X"8FA40020";
        ram_buffer(14563) := X"24420001";
        ram_buffer(14564) := X"AC620000";
        ram_buffer(14565) := X"8E8200E4";
        ram_buffer(14566) := X"8EA30038";
        ram_buffer(14567) := X"00000000";
        ram_buffer(14568) := X"00431821";
        ram_buffer(14569) := X"0064202A";
        ram_buffer(14570) := X"10800029";
        ram_buffer(14571) := X"00000000";
        ram_buffer(14572) := X"AEA30038";
        ram_buffer(14573) := X"8EA30034";
        ram_buffer(14574) := X"8FA40020";
        ram_buffer(14575) := X"00000000";
        ram_buffer(14576) := X"0064202A";
        ram_buffer(14577) := X"14800003";
        ram_buffer(14578) := X"00000000";
        ram_buffer(14579) := X"AEA00034";
        ram_buffer(14580) := X"00001821";
        ram_buffer(14581) := X"00431021";
        ram_buffer(14582) := X"1000FF6A";
        ram_buffer(14583) := X"AEA2003C";
        ram_buffer(14584) := X"8E830034";
        ram_buffer(14585) := X"00000000";
        ram_buffer(14586) := X"1860FFB7";
        ram_buffer(14587) := X"00009021";
        ram_buffer(14588) := X"8E8200E4";
        ram_buffer(14589) := X"8FB0001C";
        ram_buffer(14590) := X"1840000F";
        ram_buffer(14591) := X"24160001";
        ram_buffer(14592) := X"8E060000";
        ram_buffer(14593) := X"8E820018";
        ram_buffer(14594) := X"00163823";
        ram_buffer(14595) := X"AFA20014";
        ram_buffer(14596) := X"AFB10010";
        ram_buffer(14597) := X"00002821";
        ram_buffer(14598) := X"0C0264BB";
        ram_buffer(14599) := X"00C02021";
        ram_buffer(14600) := X"8E8200E4";
        ram_buffer(14601) := X"26D60001";
        ram_buffer(14602) := X"0056182A";
        ram_buffer(14603) := X"1060FFF4";
        ram_buffer(14604) := X"00000000";
        ram_buffer(14605) := X"8E830034";
        ram_buffer(14606) := X"26520001";
        ram_buffer(14607) := X"0243202A";
        ram_buffer(14608) := X"1480FFED";
        ram_buffer(14609) := X"26100004";
        ram_buffer(14610) := X"1000FF9F";
        ram_buffer(14611) := X"00000000";
        ram_buffer(14612) := X"1000FFD8";
        ram_buffer(14613) := X"AEA00038";
        ram_buffer(14614) := X"27BDFFB0";
        ram_buffer(14615) := X"AFB70044";
        ram_buffer(14616) := X"AFBF004C";
        ram_buffer(14617) := X"AFBE0048";
        ram_buffer(14618) := X"AFB60040";
        ram_buffer(14619) := X"AFB5003C";
        ram_buffer(14620) := X"AFB40038";
        ram_buffer(14621) := X"AFB30034";
        ram_buffer(14622) := X"AFB20030";
        ram_buffer(14623) := X"AFB1002C";
        ram_buffer(14624) := X"AFB00028";
        ram_buffer(14625) := X"14A0003E";
        ram_buffer(14626) := X"0080B821";
        ram_buffer(14627) := X"8EE20004";
        ram_buffer(14628) := X"24060040";
        ram_buffer(14629) := X"8C420000";
        ram_buffer(14630) := X"24050001";
        ram_buffer(14631) := X"0040F809";
        ram_buffer(14632) := X"02E02021";
        ram_buffer(14633) := X"0040B021";
        ram_buffer(14634) := X"8EE2015C";
        ram_buffer(14635) := X"00000000";
        ram_buffer(14636) := X"8C430008";
        ram_buffer(14637) := X"3C021009";
        ram_buffer(14638) := X"2442DD78";
        ram_buffer(14639) := X"AEF6014C";
        ram_buffer(14640) := X"14600037";
        ram_buffer(14641) := X"AEC20000";
        ram_buffer(14642) := X"8EE30034";
        ram_buffer(14643) := X"3C021009";
        ram_buffer(14644) := X"2442DDDC";
        ram_buffer(14645) := X"AEC20004";
        ram_buffer(14646) := X"8EF0003C";
        ram_buffer(14647) := X"1860001C";
        ram_buffer(14648) := X"26D10008";
        ram_buffer(14649) := X"00009021";
        ram_buffer(14650) := X"8E02001C";
        ram_buffer(14651) := X"8EE600E0";
        ram_buffer(14652) := X"000210C0";
        ram_buffer(14653) := X"00460018";
        ram_buffer(14654) := X"8E020008";
        ram_buffer(14655) := X"8EE30004";
        ram_buffer(14656) := X"8EE700E4";
        ram_buffer(14657) := X"8C630008";
        ram_buffer(14658) := X"24050001";
        ram_buffer(14659) := X"02E02021";
        ram_buffer(14660) := X"26520001";
        ram_buffer(14661) := X"26310004";
        ram_buffer(14662) := X"00003012";
        ram_buffer(14663) := X"00000000";
        ram_buffer(14664) := X"00000000";
        ram_buffer(14665) := X"14400002";
        ram_buffer(14666) := X"00C2001A";
        ram_buffer(14667) := X"0007000D";
        ram_buffer(14668) := X"00003012";
        ram_buffer(14669) := X"0060F809";
        ram_buffer(14670) := X"26100054";
        ram_buffer(14671) := X"8EE30034";
        ram_buffer(14672) := X"00000000";
        ram_buffer(14673) := X"0243182A";
        ram_buffer(14674) := X"1460FFE7";
        ram_buffer(14675) := X"AE22FFFC";
        ram_buffer(14676) := X"8FBF004C";
        ram_buffer(14677) := X"8FBE0048";
        ram_buffer(14678) := X"8FB70044";
        ram_buffer(14679) := X"8FB60040";
        ram_buffer(14680) := X"8FB5003C";
        ram_buffer(14681) := X"8FB40038";
        ram_buffer(14682) := X"8FB30034";
        ram_buffer(14683) := X"8FB20030";
        ram_buffer(14684) := X"8FB1002C";
        ram_buffer(14685) := X"8FB00028";
        ram_buffer(14686) := X"03E00008";
        ram_buffer(14687) := X"27BD0050";
        ram_buffer(14688) := X"8C820000";
        ram_buffer(14689) := X"24050004";
        ram_buffer(14690) := X"8C430000";
        ram_buffer(14691) := X"00000000";
        ram_buffer(14692) := X"0060F809";
        ram_buffer(14693) := X"AC450014";
        ram_buffer(14694) := X"1000FFBC";
        ram_buffer(14695) := X"00000000";
        ram_buffer(14696) := X"8EE60034";
        ram_buffer(14697) := X"8EF100E4";
        ram_buffer(14698) := X"00061080";
        ram_buffer(14699) := X"00463021";
        ram_buffer(14700) := X"00D10018";
        ram_buffer(14701) := X"8EE20004";
        ram_buffer(14702) := X"24050001";
        ram_buffer(14703) := X"8C430000";
        ram_buffer(14704) := X"3C021009";
        ram_buffer(14705) := X"2442E128";
        ram_buffer(14706) := X"AEC20004";
        ram_buffer(14707) := X"02E02021";
        ram_buffer(14708) := X"00003012";
        ram_buffer(14709) := X"0060F809";
        ram_buffer(14710) := X"00063080";
        ram_buffer(14711) := X"00408021";
        ram_buffer(14712) := X"8EE20034";
        ram_buffer(14713) := X"8EF3003C";
        ram_buffer(14714) := X"1840FFD9";
        ram_buffer(14715) := X"00119040";
        ram_buffer(14716) := X"02511821";
        ram_buffer(14717) := X"00111080";
        ram_buffer(14718) := X"0011A900";
        ram_buffer(14719) := X"AFA20018";
        ram_buffer(14720) := X"AFA30010";
        ram_buffer(14721) := X"02A21023";
        ram_buffer(14722) := X"001118C0";
        ram_buffer(14723) := X"26D20008";
        ram_buffer(14724) := X"AFA20014";
        ram_buffer(14725) := X"AFA3001C";
        ram_buffer(14726) := X"0000B021";
        ram_buffer(14727) := X"AFA20020";
        ram_buffer(14728) := X"8E62001C";
        ram_buffer(14729) := X"8EE600E0";
        ram_buffer(14730) := X"000210C0";
        ram_buffer(14731) := X"00460018";
        ram_buffer(14732) := X"8E620008";
        ram_buffer(14733) := X"8EE30004";
        ram_buffer(14734) := X"8FA80018";
        ram_buffer(14735) := X"8C630008";
        ram_buffer(14736) := X"8FA70010";
        ram_buffer(14737) := X"24050001";
        ram_buffer(14738) := X"02E02021";
        ram_buffer(14739) := X"00003012";
        ram_buffer(14740) := X"00000000";
        ram_buffer(14741) := X"00000000";
        ram_buffer(14742) := X"14400002";
        ram_buffer(14743) := X"00C2001A";
        ram_buffer(14744) := X"0007000D";
        ram_buffer(14745) := X"00003012";
        ram_buffer(14746) := X"0060F809";
        ram_buffer(14747) := X"0208A021";
        ram_buffer(14748) := X"8FA60014";
        ram_buffer(14749) := X"00402821";
        ram_buffer(14750) := X"02802021";
        ram_buffer(14751) := X"0C027F93";
        ram_buffer(14752) := X"0040F021";
        ram_buffer(14753) := X"1A200010";
        ram_buffer(14754) := X"00000000";
        ram_buffer(14755) := X"8FA2001C";
        ram_buffer(14756) := X"8FA40020";
        ram_buffer(14757) := X"03C22821";
        ram_buffer(14758) := X"02001821";
        ram_buffer(14759) := X"03C01021";
        ram_buffer(14760) := X"02842021";
        ram_buffer(14761) := X"8CA60000";
        ram_buffer(14762) := X"24630004";
        ram_buffer(14763) := X"AC66FFFC";
        ram_buffer(14764) := X"8C460000";
        ram_buffer(14765) := X"24A50004";
        ram_buffer(14766) := X"AC860000";
        ram_buffer(14767) := X"24420004";
        ram_buffer(14768) := X"1683FFF8";
        ram_buffer(14769) := X"24840004";
        ram_buffer(14770) := X"8EE20034";
        ram_buffer(14771) := X"26D60001";
        ram_buffer(14772) := X"02C2102A";
        ram_buffer(14773) := X"AE540000";
        ram_buffer(14774) := X"02958021";
        ram_buffer(14775) := X"26730054";
        ram_buffer(14776) := X"1440FFCF";
        ram_buffer(14777) := X"26520004";
        ram_buffer(14778) := X"1000FF99";
        ram_buffer(14779) := X"00000000";
        ram_buffer(14780) := X"27BDFFE8";
        ram_buffer(14781) := X"8C8200EC";
        ram_buffer(14782) := X"AFB00010";
        ram_buffer(14783) := X"8C900150";
        ram_buffer(14784) := X"28420002";
        ram_buffer(14785) := X"AFBF0014";
        ram_buffer(14786) := X"14400024";
        ram_buffer(14787) := X"AE000008";
        ram_buffer(14788) := X"24020001";
        ram_buffer(14789) := X"AE020014";
        ram_buffer(14790) := X"24020002";
        ram_buffer(14791) := X"AE00000C";
        ram_buffer(14792) := X"10A2002A";
        ram_buffer(14793) := X"AE000010";
        ram_buffer(14794) := X"24020003";
        ram_buffer(14795) := X"10A20032";
        ram_buffer(14796) := X"00000000";
        ram_buffer(14797) := X"10A00008";
        ram_buffer(14798) := X"24030004";
        ram_buffer(14799) := X"8C820000";
        ram_buffer(14800) := X"8FBF0014";
        ram_buffer(14801) := X"8FB00010";
        ram_buffer(14802) := X"8C590000";
        ram_buffer(14803) := X"AC430014";
        ram_buffer(14804) := X"03200008";
        ram_buffer(14805) := X"27BD0018";
        ram_buffer(14806) := X"8E020040";
        ram_buffer(14807) := X"00000000";
        ram_buffer(14808) := X"10400007";
        ram_buffer(14809) := X"24050004";
        ram_buffer(14810) := X"8C820000";
        ram_buffer(14811) := X"00000000";
        ram_buffer(14812) := X"8C430000";
        ram_buffer(14813) := X"00000000";
        ram_buffer(14814) := X"0060F809";
        ram_buffer(14815) := X"AC450014";
        ram_buffer(14816) := X"8FBF0014";
        ram_buffer(14817) := X"3C021009";
        ram_buffer(14818) := X"2442F200";
        ram_buffer(14819) := X"AE020004";
        ram_buffer(14820) := X"8FB00010";
        ram_buffer(14821) := X"03E00008";
        ram_buffer(14822) := X"27BD0018";
        ram_buffer(14823) := X"8C8300E8";
        ram_buffer(14824) := X"24020001";
        ram_buffer(14825) := X"1062001F";
        ram_buffer(14826) := X"00000000";
        ram_buffer(14827) := X"8C8200F0";
        ram_buffer(14828) := X"00000000";
        ram_buffer(14829) := X"8C42000C";
        ram_buffer(14830) := X"AE00000C";
        ram_buffer(14831) := X"AE020014";
        ram_buffer(14832) := X"24020002";
        ram_buffer(14833) := X"14A2FFD8";
        ram_buffer(14834) := X"AE000010";
        ram_buffer(14835) := X"8E020040";
        ram_buffer(14836) := X"00000000";
        ram_buffer(14837) := X"10400018";
        ram_buffer(14838) := X"00000000";
        ram_buffer(14839) := X"8FBF0014";
        ram_buffer(14840) := X"3C021009";
        ram_buffer(14841) := X"2442E878";
        ram_buffer(14842) := X"AE020004";
        ram_buffer(14843) := X"8FB00010";
        ram_buffer(14844) := X"03E00008";
        ram_buffer(14845) := X"27BD0018";
        ram_buffer(14846) := X"8E020040";
        ram_buffer(14847) := X"00000000";
        ram_buffer(14848) := X"10400015";
        ram_buffer(14849) := X"24050004";
        ram_buffer(14850) := X"8FBF0014";
        ram_buffer(14851) := X"3C021009";
        ram_buffer(14852) := X"2442EEF4";
        ram_buffer(14853) := X"AE020004";
        ram_buffer(14854) := X"8FB00010";
        ram_buffer(14855) := X"03E00008";
        ram_buffer(14856) := X"27BD0018";
        ram_buffer(14857) := X"8C8200F0";
        ram_buffer(14858) := X"00000000";
        ram_buffer(14859) := X"8C420048";
        ram_buffer(14860) := X"1000FFB9";
        ram_buffer(14861) := X"AE020014";
        ram_buffer(14862) := X"8C820000";
        ram_buffer(14863) := X"24050004";
        ram_buffer(14864) := X"8C430000";
        ram_buffer(14865) := X"00000000";
        ram_buffer(14866) := X"0060F809";
        ram_buffer(14867) := X"AC450014";
        ram_buffer(14868) := X"1000FFE2";
        ram_buffer(14869) := X"00000000";
        ram_buffer(14870) := X"8C820000";
        ram_buffer(14871) := X"00000000";
        ram_buffer(14872) := X"8C430000";
        ram_buffer(14873) := X"00000000";
        ram_buffer(14874) := X"0060F809";
        ram_buffer(14875) := X"AC450014";
        ram_buffer(14876) := X"1000FFE5";
        ram_buffer(14877) := X"00000000";
        ram_buffer(14878) := X"8C8300EC";
        ram_buffer(14879) := X"27BDFFA0";
        ram_buffer(14880) := X"AFB1003C";
        ram_buffer(14881) := X"AFB00038";
        ram_buffer(14882) := X"AFBF005C";
        ram_buffer(14883) := X"AFBE0058";
        ram_buffer(14884) := X"AFB70054";
        ram_buffer(14885) := X"AFB60050";
        ram_buffer(14886) := X"AFB5004C";
        ram_buffer(14887) := X"AFB40048";
        ram_buffer(14888) := X"AFB30044";
        ram_buffer(14889) := X"AFB20040";
        ram_buffer(14890) := X"8C900150";
        ram_buffer(14891) := X"1860001B";
        ram_buffer(14892) := X"00808821";
        ram_buffer(14893) := X"249400F0";
        ram_buffer(14894) := X"27B30018";
        ram_buffer(14895) := X"00009021";
        ram_buffer(14896) := X"8E820000";
        ram_buffer(14897) := X"8E060008";
        ram_buffer(14898) := X"8C47000C";
        ram_buffer(14899) := X"8C420004";
        ram_buffer(14900) := X"00E60018";
        ram_buffer(14901) := X"24420010";
        ram_buffer(14902) := X"00021080";
        ram_buffer(14903) := X"8E230004";
        ram_buffer(14904) := X"02021021";
        ram_buffer(14905) := X"8C450000";
        ram_buffer(14906) := X"AFA00010";
        ram_buffer(14907) := X"8C620020";
        ram_buffer(14908) := X"02202021";
        ram_buffer(14909) := X"26520001";
        ram_buffer(14910) := X"26940004";
        ram_buffer(14911) := X"00003012";
        ram_buffer(14912) := X"0040F809";
        ram_buffer(14913) := X"26730004";
        ram_buffer(14914) := X"8E2300EC";
        ram_buffer(14915) := X"AE62FFFC";
        ram_buffer(14916) := X"0243102A";
        ram_buffer(14917) := X"1440FFEA";
        ram_buffer(14918) := X"00000000";
        ram_buffer(14919) := X"8E130010";
        ram_buffer(14920) := X"8E040014";
        ram_buffer(14921) := X"00000000";
        ram_buffer(14922) := X"0264102A";
        ram_buffer(14923) := X"10400147";
        ram_buffer(14924) := X"26620003";
        ram_buffer(14925) := X"00021080";
        ram_buffer(14926) := X"00402821";
        ram_buffer(14927) := X"24B5FFF4";
        ram_buffer(14928) := X"24A5FFF8";
        ram_buffer(14929) := X"AFA5002C";
        ram_buffer(14930) := X"26050018";
        ram_buffer(14931) := X"AFA50030";
        ram_buffer(14932) := X"3C057FFF";
        ram_buffer(14933) := X"AFA20028";
        ram_buffer(14934) := X"34A5FFFF";
        ram_buffer(14935) := X"8E12000C";
        ram_buffer(14936) := X"8E220100";
        ram_buffer(14937) := X"24140001";
        ram_buffer(14938) := X"AFA50034";
        ram_buffer(14939) := X"0242282B";
        ram_buffer(14940) := X"10A0012A";
        ram_buffer(14941) := X"24160003";
        ram_buffer(14942) := X"1860004E";
        ram_buffer(14943) := X"27B90018";
        ram_buffer(14944) := X"00031880";
        ram_buffer(14945) := X"263F00F0";
        ram_buffer(14946) := X"0323B821";
        ram_buffer(14947) := X"00002021";
        ram_buffer(14948) := X"240B0004";
        ram_buffer(14949) := X"24180005";
        ram_buffer(14950) := X"240F0006";
        ram_buffer(14951) := X"240E0007";
        ram_buffer(14952) := X"240D0008";
        ram_buffer(14953) := X"240C0009";
        ram_buffer(14954) := X"8FE20000";
        ram_buffer(14955) := X"00000000";
        ram_buffer(14956) := X"8C450034";
        ram_buffer(14957) := X"8C420038";
        ram_buffer(14958) := X"00000000";
        ram_buffer(14959) := X"1840003A";
        ram_buffer(14960) := X"000549C0";
        ram_buffer(14961) := X"02490018";
        ram_buffer(14962) := X"8F230000";
        ram_buffer(14963) := X"00004812";
        ram_buffer(14964) := X"18A00035";
        ram_buffer(14965) := X"00000000";
        ram_buffer(14966) := X"10B40048";
        ram_buffer(14967) := X"24060002";
        ram_buffer(14968) := X"10A600D4";
        ram_buffer(14969) := X"00753021";
        ram_buffer(14970) := X"10B60098";
        ram_buffer(14971) := X"02625021";
        ram_buffer(14972) := X"000A5080";
        ram_buffer(14973) := X"00753021";
        ram_buffer(14974) := X"1000001A";
        ram_buffer(14975) := X"006A5021";
        ram_buffer(14976) := X"249E0005";
        ram_buffer(14977) := X"24680280";
        ram_buffer(14978) := X"10B80024";
        ram_buffer(14979) := X"AC470028";
        ram_buffer(14980) := X"249E0006";
        ram_buffer(14981) := X"24670300";
        ram_buffer(14982) := X"10AF0020";
        ram_buffer(14983) := X"AC48002C";
        ram_buffer(14984) := X"249E0007";
        ram_buffer(14985) := X"24680380";
        ram_buffer(14986) := X"10AE001C";
        ram_buffer(14987) := X"AC470030";
        ram_buffer(14988) := X"249E0008";
        ram_buffer(14989) := X"24670400";
        ram_buffer(14990) := X"10AD0018";
        ram_buffer(14991) := X"AC480034";
        ram_buffer(14992) := X"24880009";
        ram_buffer(14993) := X"24630480";
        ram_buffer(14994) := X"10AC002A";
        ram_buffer(14995) := X"AC470038";
        ram_buffer(14996) := X"2484000A";
        ram_buffer(14997) := X"AC43003C";
        ram_buffer(14998) := X"24C60004";
        ram_buffer(14999) := X"10CA0012";
        ram_buffer(15000) := X"00000000";
        ram_buffer(15001) := X"8CC30000";
        ram_buffer(15002) := X"00041080";
        ram_buffer(15003) := X"00691821";
        ram_buffer(15004) := X"02021021";
        ram_buffer(15005) := X"247E0080";
        ram_buffer(15006) := X"24670100";
        ram_buffer(15007) := X"24680180";
        ram_buffer(15008) := X"AC5E001C";
        ram_buffer(15009) := X"AC470020";
        ram_buffer(15010) := X"AC430018";
        ram_buffer(15011) := X"249E0004";
        ram_buffer(15012) := X"24670200";
        ram_buffer(15013) := X"14ABFFDA";
        ram_buffer(15014) := X"AC480024";
        ram_buffer(15015) := X"24C60004";
        ram_buffer(15016) := X"14CAFFF0";
        ram_buffer(15017) := X"03C02021";
        ram_buffer(15018) := X"27390004";
        ram_buffer(15019) := X"1737FFBE";
        ram_buffer(15020) := X"27FF0004";
        ram_buffer(15021) := X"8E220164";
        ram_buffer(15022) := X"8FA50030";
        ram_buffer(15023) := X"8C420004";
        ram_buffer(15024) := X"00000000";
        ram_buffer(15025) := X"0040F809";
        ram_buffer(15026) := X"02202021";
        ram_buffer(15027) := X"104000EB";
        ram_buffer(15028) := X"00000000";
        ram_buffer(15029) := X"8E220100";
        ram_buffer(15030) := X"26520001";
        ram_buffer(15031) := X"0242182B";
        ram_buffer(15032) := X"106000CC";
        ram_buffer(15033) := X"00000000";
        ram_buffer(15034) := X"8E2300EC";
        ram_buffer(15035) := X"1000FFA2";
        ram_buffer(15036) := X"00000000";
        ram_buffer(15037) := X"1000FFD8";
        ram_buffer(15038) := X"01002021";
        ram_buffer(15039) := X"00752821";
        ram_buffer(15040) := X"8CA70000";
        ram_buffer(15041) := X"24860006";
        ram_buffer(15042) := X"00063080";
        ram_buffer(15043) := X"02063021";
        ram_buffer(15044) := X"00E93821";
        ram_buffer(15045) := X"10540047";
        ram_buffer(15046) := X"ACC70000";
        ram_buffer(15047) := X"8FA6002C";
        ram_buffer(15048) := X"00000000";
        ram_buffer(15049) := X"00663021";
        ram_buffer(15050) := X"8CC80000";
        ram_buffer(15051) := X"24860007";
        ram_buffer(15052) := X"00063880";
        ram_buffer(15053) := X"02073821";
        ram_buffer(15054) := X"01094021";
        ram_buffer(15055) := X"ACE80000";
        ram_buffer(15056) := X"24070002";
        ram_buffer(15057) := X"1047003B";
        ram_buffer(15058) := X"00000000";
        ram_buffer(15059) := X"8CA80008";
        ram_buffer(15060) := X"24870008";
        ram_buffer(15061) := X"00073880";
        ram_buffer(15062) := X"02073821";
        ram_buffer(15063) := X"01094021";
        ram_buffer(15064) := X"10560034";
        ram_buffer(15065) := X"ACE80000";
        ram_buffer(15066) := X"8FA70028";
        ram_buffer(15067) := X"00000000";
        ram_buffer(15068) := X"00671821";
        ram_buffer(15069) := X"8C670000";
        ram_buffer(15070) := X"24830009";
        ram_buffer(15071) := X"00031880";
        ram_buffer(15072) := X"02031821";
        ram_buffer(15073) := X"00E93821";
        ram_buffer(15074) := X"104B002A";
        ram_buffer(15075) := X"AC670000";
        ram_buffer(15076) := X"8CA70010";
        ram_buffer(15077) := X"2483000A";
        ram_buffer(15078) := X"00031880";
        ram_buffer(15079) := X"02031821";
        ram_buffer(15080) := X"00E93821";
        ram_buffer(15081) := X"10580023";
        ram_buffer(15082) := X"AC670000";
        ram_buffer(15083) := X"8CA70014";
        ram_buffer(15084) := X"2483000B";
        ram_buffer(15085) := X"00031880";
        ram_buffer(15086) := X"02031821";
        ram_buffer(15087) := X"00E93821";
        ram_buffer(15088) := X"104F001C";
        ram_buffer(15089) := X"AC670000";
        ram_buffer(15090) := X"8CA70018";
        ram_buffer(15091) := X"2483000C";
        ram_buffer(15092) := X"00031880";
        ram_buffer(15093) := X"02031821";
        ram_buffer(15094) := X"00E93821";
        ram_buffer(15095) := X"104E0015";
        ram_buffer(15096) := X"AC670000";
        ram_buffer(15097) := X"8CA7001C";
        ram_buffer(15098) := X"2483000D";
        ram_buffer(15099) := X"00031880";
        ram_buffer(15100) := X"02031821";
        ram_buffer(15101) := X"00E93821";
        ram_buffer(15102) := X"104D000E";
        ram_buffer(15103) := X"AC670000";
        ram_buffer(15104) := X"8CA60020";
        ram_buffer(15105) := X"2483000E";
        ram_buffer(15106) := X"00031880";
        ram_buffer(15107) := X"02031821";
        ram_buffer(15108) := X"00C93021";
        ram_buffer(15109) := X"104C0007";
        ram_buffer(15110) := X"AC660000";
        ram_buffer(15111) := X"8CA50024";
        ram_buffer(15112) := X"2483000F";
        ram_buffer(15113) := X"00031880";
        ram_buffer(15114) := X"02031821";
        ram_buffer(15115) := X"00A94821";
        ram_buffer(15116) := X"AC690000";
        ram_buffer(15117) := X"00442021";
        ram_buffer(15118) := X"27390004";
        ram_buffer(15119) := X"1737FF5A";
        ram_buffer(15120) := X"27FF0004";
        ram_buffer(15121) := X"1000FF9B";
        ram_buffer(15122) := X"00000000";
        ram_buffer(15123) := X"00753821";
        ram_buffer(15124) := X"8CE60000";
        ram_buffer(15125) := X"00042880";
        ram_buffer(15126) := X"00C93021";
        ram_buffer(15127) := X"02052821";
        ram_buffer(15128) := X"24CA0080";
        ram_buffer(15129) := X"24C80100";
        ram_buffer(15130) := X"ACAA001C";
        ram_buffer(15131) := X"ACA60018";
        ram_buffer(15132) := X"248A0003";
        ram_buffer(15133) := X"10540027";
        ram_buffer(15134) := X"ACA80020";
        ram_buffer(15135) := X"8FA5002C";
        ram_buffer(15136) := X"00000000";
        ram_buffer(15137) := X"00652821";
        ram_buffer(15138) := X"8CA60000";
        ram_buffer(15139) := X"000A2880";
        ram_buffer(15140) := X"00C93021";
        ram_buffer(15141) := X"02052821";
        ram_buffer(15142) := X"24CA0080";
        ram_buffer(15143) := X"24C80100";
        ram_buffer(15144) := X"ACA60018";
        ram_buffer(15145) := X"ACAA001C";
        ram_buffer(15146) := X"ACA80020";
        ram_buffer(15147) := X"24050002";
        ram_buffer(15148) := X"10450018";
        ram_buffer(15149) := X"24860006";
        ram_buffer(15150) := X"8CE50008";
        ram_buffer(15151) := X"00063080";
        ram_buffer(15152) := X"00A92821";
        ram_buffer(15153) := X"02063021";
        ram_buffer(15154) := X"24A80080";
        ram_buffer(15155) := X"24A70100";
        ram_buffer(15156) := X"ACC50018";
        ram_buffer(15157) := X"ACC8001C";
        ram_buffer(15158) := X"24850009";
        ram_buffer(15159) := X"1056000D";
        ram_buffer(15160) := X"ACC70020";
        ram_buffer(15161) := X"8FA60028";
        ram_buffer(15162) := X"00000000";
        ram_buffer(15163) := X"00661821";
        ram_buffer(15164) := X"8C660000";
        ram_buffer(15165) := X"00051880";
        ram_buffer(15166) := X"00C94821";
        ram_buffer(15167) := X"02031821";
        ram_buffer(15168) := X"25260080";
        ram_buffer(15169) := X"25250100";
        ram_buffer(15170) := X"AC690018";
        ram_buffer(15171) := X"AC66001C";
        ram_buffer(15172) := X"AC650020";
        ram_buffer(15173) := X"00021840";
        ram_buffer(15174) := X"00621021";
        ram_buffer(15175) := X"27390004";
        ram_buffer(15176) := X"00442021";
        ram_buffer(15177) := X"1737FF20";
        ram_buffer(15178) := X"27FF0004";
        ram_buffer(15179) := X"1000FF61";
        ram_buffer(15180) := X"00000000";
        ram_buffer(15181) := X"8CC70000";
        ram_buffer(15182) := X"00042880";
        ram_buffer(15183) := X"00E93821";
        ram_buffer(15184) := X"02052821";
        ram_buffer(15185) := X"24E80080";
        ram_buffer(15186) := X"ACA70018";
        ram_buffer(15187) := X"248A0002";
        ram_buffer(15188) := X"10540029";
        ram_buffer(15189) := X"ACA8001C";
        ram_buffer(15190) := X"8FA5002C";
        ram_buffer(15191) := X"00000000";
        ram_buffer(15192) := X"00652821";
        ram_buffer(15193) := X"8CA70000";
        ram_buffer(15194) := X"000A2880";
        ram_buffer(15195) := X"00E93821";
        ram_buffer(15196) := X"02052821";
        ram_buffer(15197) := X"24E80080";
        ram_buffer(15198) := X"ACA70018";
        ram_buffer(15199) := X"ACA8001C";
        ram_buffer(15200) := X"24050002";
        ram_buffer(15201) := X"1045001C";
        ram_buffer(15202) := X"24870004";
        ram_buffer(15203) := X"8CC50008";
        ram_buffer(15204) := X"00073880";
        ram_buffer(15205) := X"00A92821";
        ram_buffer(15206) := X"02073821";
        ram_buffer(15207) := X"24A80080";
        ram_buffer(15208) := X"ACE50018";
        ram_buffer(15209) := X"ACE8001C";
        ram_buffer(15210) := X"10560013";
        ram_buffer(15211) := X"24850006";
        ram_buffer(15212) := X"8FA70028";
        ram_buffer(15213) := X"00052880";
        ram_buffer(15214) := X"00671821";
        ram_buffer(15215) := X"8C630000";
        ram_buffer(15216) := X"02052821";
        ram_buffer(15217) := X"00691821";
        ram_buffer(15218) := X"24670080";
        ram_buffer(15219) := X"ACA30018";
        ram_buffer(15220) := X"ACA7001C";
        ram_buffer(15221) := X"104B0008";
        ram_buffer(15222) := X"24830008";
        ram_buffer(15223) := X"8CC50010";
        ram_buffer(15224) := X"00031880";
        ram_buffer(15225) := X"00A94821";
        ram_buffer(15226) := X"02031821";
        ram_buffer(15227) := X"25250080";
        ram_buffer(15228) := X"AC690018";
        ram_buffer(15229) := X"AC65001C";
        ram_buffer(15230) := X"8FA30034";
        ram_buffer(15231) := X"00000000";
        ram_buffer(15232) := X"00431021";
        ram_buffer(15233) := X"00021040";
        ram_buffer(15234) := X"24420002";
        ram_buffer(15235) := X"1000FF8A";
        ram_buffer(15236) := X"00442021";
        ram_buffer(15237) := X"8E040014";
        ram_buffer(15238) := X"8E2300EC";
        ram_buffer(15239) := X"8FA60028";
        ram_buffer(15240) := X"26730001";
        ram_buffer(15241) := X"24C60004";
        ram_buffer(15242) := X"AFA60028";
        ram_buffer(15243) := X"8FA6002C";
        ram_buffer(15244) := X"0264282A";
        ram_buffer(15245) := X"24C60004";
        ram_buffer(15246) := X"AE00000C";
        ram_buffer(15247) := X"26B50004";
        ram_buffer(15248) := X"AFA6002C";
        ram_buffer(15249) := X"14A0FEC9";
        ram_buffer(15250) := X"00009021";
        ram_buffer(15251) := X"8E020008";
        ram_buffer(15252) := X"28630002";
        ram_buffer(15253) := X"24420001";
        ram_buffer(15254) := X"AE020008";
        ram_buffer(15255) := X"8E220150";
        ram_buffer(15256) := X"14600014";
        ram_buffer(15257) := X"24030001";
        ram_buffer(15258) := X"AC430014";
        ram_buffer(15259) := X"AC40000C";
        ram_buffer(15260) := X"AC400010";
        ram_buffer(15261) := X"10000003";
        ram_buffer(15262) := X"24020001";
        ram_buffer(15263) := X"AE130010";
        ram_buffer(15264) := X"AE12000C";
        ram_buffer(15265) := X"8FBF005C";
        ram_buffer(15266) := X"8FBE0058";
        ram_buffer(15267) := X"8FB70054";
        ram_buffer(15268) := X"8FB60050";
        ram_buffer(15269) := X"8FB5004C";
        ram_buffer(15270) := X"8FB40048";
        ram_buffer(15271) := X"8FB30044";
        ram_buffer(15272) := X"8FB20040";
        ram_buffer(15273) := X"8FB1003C";
        ram_buffer(15274) := X"8FB00038";
        ram_buffer(15275) := X"03E00008";
        ram_buffer(15276) := X"27BD0060";
        ram_buffer(15277) := X"8E2400E8";
        ram_buffer(15278) := X"8C430008";
        ram_buffer(15279) := X"2484FFFF";
        ram_buffer(15280) := X"0064182B";
        ram_buffer(15281) := X"10600006";
        ram_buffer(15282) := X"00000000";
        ram_buffer(15283) := X"8E2300F0";
        ram_buffer(15284) := X"00000000";
        ram_buffer(15285) := X"8C63000C";
        ram_buffer(15286) := X"1000FFE4";
        ram_buffer(15287) := X"AC430014";
        ram_buffer(15288) := X"8E2300F0";
        ram_buffer(15289) := X"00000000";
        ram_buffer(15290) := X"8C630048";
        ram_buffer(15291) := X"1000FFDF";
        ram_buffer(15292) := X"AC430014";
        ram_buffer(15293) := X"27BDFF88";
        ram_buffer(15294) := X"8C8300E8";
        ram_buffer(15295) := X"8C820034";
        ram_buffer(15296) := X"AFB10054";
        ram_buffer(15297) := X"00808821";
        ram_buffer(15298) := X"8C840150";
        ram_buffer(15299) := X"2463FFFF";
        ram_buffer(15300) := X"AFB3005C";
        ram_buffer(15301) := X"AFBF0074";
        ram_buffer(15302) := X"AFBE0070";
        ram_buffer(15303) := X"AFB7006C";
        ram_buffer(15304) := X"AFB60068";
        ram_buffer(15305) := X"AFB50064";
        ram_buffer(15306) := X"AFB40060";
        ram_buffer(15307) := X"AFB20058";
        ram_buffer(15308) := X"AFB00050";
        ram_buffer(15309) := X"AFA50044";
        ram_buffer(15310) := X"AFA40034";
        ram_buffer(15311) := X"AFA30038";
        ram_buffer(15312) := X"8E33003C";
        ram_buffer(15313) := X"18400070";
        ram_buffer(15314) := X"24820040";
        ram_buffer(15315) := X"AFA20030";
        ram_buffer(15316) := X"8FA20044";
        ram_buffer(15317) := X"AFA0003C";
        ram_buffer(15318) := X"AFA20020";
        ram_buffer(15319) := X"3C0201FF";
        ram_buffer(15320) := X"3442FFFF";
        ram_buffer(15321) := X"AFA20048";
        ram_buffer(15322) := X"8FB00034";
        ram_buffer(15323) := X"8E67000C";
        ram_buffer(15324) := X"8E060008";
        ram_buffer(15325) := X"8FA30030";
        ram_buffer(15326) := X"00E60018";
        ram_buffer(15327) := X"8E220004";
        ram_buffer(15328) := X"8C650000";
        ram_buffer(15329) := X"24030001";
        ram_buffer(15330) := X"AFA30010";
        ram_buffer(15331) := X"8C420020";
        ram_buffer(15332) := X"00003012";
        ram_buffer(15333) := X"0040F809";
        ram_buffer(15334) := X"02202021";
        ram_buffer(15335) := X"AFA20040";
        ram_buffer(15336) := X"8FA30038";
        ram_buffer(15337) := X"8E020008";
        ram_buffer(15338) := X"8E72000C";
        ram_buffer(15339) := X"0043182B";
        ram_buffer(15340) := X"1460000A";
        ram_buffer(15341) := X"00000000";
        ram_buffer(15342) := X"8E630020";
        ram_buffer(15343) := X"00000000";
        ram_buffer(15344) := X"16400002";
        ram_buffer(15345) := X"0072001B";
        ram_buffer(15346) := X"0007000D";
        ram_buffer(15347) := X"00001810";
        ram_buffer(15348) := X"10600002";
        ram_buffer(15349) := X"00000000";
        ram_buffer(15350) := X"00609021";
        ram_buffer(15351) := X"8E75001C";
        ram_buffer(15352) := X"8E700008";
        ram_buffer(15353) := X"00000000";
        ram_buffer(15354) := X"16000002";
        ram_buffer(15355) := X"02B0001B";
        ram_buffer(15356) := X"0007000D";
        ram_buffer(15357) := X"0000A010";
        ram_buffer(15358) := X"1A800002";
        ram_buffer(15359) := X"00000000";
        ram_buffer(15360) := X"0214A023";
        ram_buffer(15361) := X"1A40002D";
        ram_buffer(15362) := X"00000000";
        ram_buffer(15363) := X"001511C0";
        ram_buffer(15364) := X"AFA20028";
        ram_buffer(15365) := X"8FB70040";
        ram_buffer(15366) := X"001411C0";
        ram_buffer(15367) := X"AFA2002C";
        ram_buffer(15368) := X"0000F021";
        ram_buffer(15369) := X"8FA20020";
        ram_buffer(15370) := X"8E240160";
        ram_buffer(15371) := X"001E18C0";
        ram_buffer(15372) := X"8EF60000";
        ram_buffer(15373) := X"8C460000";
        ram_buffer(15374) := X"AFB50018";
        ram_buffer(15375) := X"AFA00014";
        ram_buffer(15376) := X"AFA30010";
        ram_buffer(15377) := X"8C830004";
        ram_buffer(15378) := X"02C03821";
        ram_buffer(15379) := X"02602821";
        ram_buffer(15380) := X"0060F809";
        ram_buffer(15381) := X"02202021";
        ram_buffer(15382) := X"1A800012";
        ram_buffer(15383) := X"00000000";
        ram_buffer(15384) := X"8FA20028";
        ram_buffer(15385) := X"00000000";
        ram_buffer(15386) := X"02C21821";
        ram_buffer(15387) := X"8FB6002C";
        ram_buffer(15388) := X"00602021";
        ram_buffer(15389) := X"02C02821";
        ram_buffer(15390) := X"0C0264DD";
        ram_buffer(15391) := X"AFA30024";
        ram_buffer(15392) := X"8FA30024";
        ram_buffer(15393) := X"00000000";
        ram_buffer(15394) := X"00601021";
        ram_buffer(15395) := X"8464FF80";
        ram_buffer(15396) := X"00561821";
        ram_buffer(15397) := X"A4440000";
        ram_buffer(15398) := X"24420080";
        ram_buffer(15399) := X"1443FFFD";
        ram_buffer(15400) := X"00000000";
        ram_buffer(15401) := X"27DE0001";
        ram_buffer(15402) := X"165EFFDE";
        ram_buffer(15403) := X"26F70004";
        ram_buffer(15404) := X"8FA20034";
        ram_buffer(15405) := X"00000000";
        ram_buffer(15406) := X"8C420008";
        ram_buffer(15407) := X"8FA30038";
        ram_buffer(15408) := X"00000000";
        ram_buffer(15409) := X"1062001D";
        ram_buffer(15410) := X"00000000";
        ram_buffer(15411) := X"8FA3003C";
        ram_buffer(15412) := X"8E220034";
        ram_buffer(15413) := X"24630001";
        ram_buffer(15414) := X"AFA3003C";
        ram_buffer(15415) := X"0062102A";
        ram_buffer(15416) := X"8FA30030";
        ram_buffer(15417) := X"26730054";
        ram_buffer(15418) := X"24630004";
        ram_buffer(15419) := X"AFA30030";
        ram_buffer(15420) := X"8FA30020";
        ram_buffer(15421) := X"00000000";
        ram_buffer(15422) := X"24630004";
        ram_buffer(15423) := X"1440FF9A";
        ram_buffer(15424) := X"AFA30020";
        ram_buffer(15425) := X"8FA50044";
        ram_buffer(15426) := X"8FBF0074";
        ram_buffer(15427) := X"8FBE0070";
        ram_buffer(15428) := X"8FB7006C";
        ram_buffer(15429) := X"8FB60068";
        ram_buffer(15430) := X"8FB50064";
        ram_buffer(15431) := X"8FB40060";
        ram_buffer(15432) := X"8FB3005C";
        ram_buffer(15433) := X"8FB20058";
        ram_buffer(15434) := X"8FB00050";
        ram_buffer(15435) := X"02202021";
        ram_buffer(15436) := X"8FB10054";
        ram_buffer(15437) := X"08023A1E";
        ram_buffer(15438) := X"27BD0078";
        ram_buffer(15439) := X"0295A021";
        ram_buffer(15440) := X"16000002";
        ram_buffer(15441) := X"0290001B";
        ram_buffer(15442) := X"0007000D";
        ram_buffer(15443) := X"8E62000C";
        ram_buffer(15444) := X"00000000";
        ram_buffer(15445) := X"0242102A";
        ram_buffer(15446) := X"0000B812";
        ram_buffer(15447) := X"1040FFDB";
        ram_buffer(15448) := X"00124080";
        ram_buffer(15449) := X"8FA20048";
        ram_buffer(15450) := X"00000000";
        ram_buffer(15451) := X"02021021";
        ram_buffer(15452) := X"000211C0";
        ram_buffer(15453) := X"AFA20028";
        ram_buffer(15454) := X"245E0080";
        ram_buffer(15455) := X"8FA20040";
        ram_buffer(15456) := X"0014B1C0";
        ram_buffer(15457) := X"0048A021";
        ram_buffer(15458) := X"8E820000";
        ram_buffer(15459) := X"02C02821";
        ram_buffer(15460) := X"AFA20024";
        ram_buffer(15461) := X"8E95FFFC";
        ram_buffer(15462) := X"0C0264DD";
        ram_buffer(15463) := X"00402021";
        ram_buffer(15464) := X"8FA20024";
        ram_buffer(15465) := X"12E0000F";
        ram_buffer(15466) := X"00000000";
        ram_buffer(15467) := X"8FA30028";
        ram_buffer(15468) := X"00003021";
        ram_buffer(15469) := X"02A32821";
        ram_buffer(15470) := X"84A30000";
        ram_buffer(15471) := X"1A000005";
        ram_buffer(15472) := X"005E2021";
        ram_buffer(15473) := X"A4430000";
        ram_buffer(15474) := X"24420080";
        ram_buffer(15475) := X"1482FFFD";
        ram_buffer(15476) := X"00000000";
        ram_buffer(15477) := X"24C60001";
        ram_buffer(15478) := X"00801021";
        ram_buffer(15479) := X"16E6FFF6";
        ram_buffer(15480) := X"00BE2821";
        ram_buffer(15481) := X"8E62000C";
        ram_buffer(15482) := X"26520001";
        ram_buffer(15483) := X"0242102A";
        ram_buffer(15484) := X"1440FFE5";
        ram_buffer(15485) := X"26940004";
        ram_buffer(15486) := X"1000FFB4";
        ram_buffer(15487) := X"00000000";
        ram_buffer(15488) := X"27BDFF78";
        ram_buffer(15489) := X"AFBE0080";
        ram_buffer(15490) := X"8C9E0150";
        ram_buffer(15491) := X"8C860100";
        ram_buffer(15492) := X"8FC20010";
        ram_buffer(15493) := X"AFA5008C";
        ram_buffer(15494) := X"00403821";
        ram_buffer(15495) := X"AFA20024";
        ram_buffer(15496) := X"8FC20014";
        ram_buffer(15497) := X"24C5FFFF";
        ram_buffer(15498) := X"00E2182A";
        ram_buffer(15499) := X"AFB7007C";
        ram_buffer(15500) := X"AFBF0084";
        ram_buffer(15501) := X"0080B821";
        ram_buffer(15502) := X"AFB60078";
        ram_buffer(15503) := X"AFB50074";
        ram_buffer(15504) := X"AFB40070";
        ram_buffer(15505) := X"AFB3006C";
        ram_buffer(15506) := X"AFB20068";
        ram_buffer(15507) := X"AFB10064";
        ram_buffer(15508) := X"AFB00060";
        ram_buffer(15509) := X"8C8400E8";
        ram_buffer(15510) := X"10600151";
        ram_buffer(15511) := X"AFA50054";
        ram_buffer(15512) := X"8FC3000C";
        ram_buffer(15513) := X"2493FFFF";
        ram_buffer(15514) := X"AFA30048";
        ram_buffer(15515) := X"00602021";
        ram_buffer(15516) := X"000718C0";
        ram_buffer(15517) := X"AFA30050";
        ram_buffer(15518) := X"00A4182B";
        ram_buffer(15519) := X"27C40018";
        ram_buffer(15520) := X"146000E2";
        ram_buffer(15521) := X"AFA40058";
        ram_buffer(15522) := X"03C0A021";
        ram_buffer(15523) := X"8EE300EC";
        ram_buffer(15524) := X"00000000";
        ram_buffer(15525) := X"186000CD";
        ram_buffer(15526) := X"26E200F0";
        ram_buffer(15527) := X"AFA20040";
        ram_buffer(15528) := X"8FA40048";
        ram_buffer(15529) := X"8FA20054";
        ram_buffer(15530) := X"8FB1008C";
        ram_buffer(15531) := X"0082102B";
        ram_buffer(15532) := X"AFA2004C";
        ram_buffer(15533) := X"8FA20040";
        ram_buffer(15534) := X"AFA00044";
        ram_buffer(15535) := X"0000A821";
        ram_buffer(15536) := X"8C500000";
        ram_buffer(15537) := X"8FA2004C";
        ram_buffer(15538) := X"00000000";
        ram_buffer(15539) := X"10400141";
        ram_buffer(15540) := X"00000000";
        ram_buffer(15541) := X"8E160034";
        ram_buffer(15542) := X"8E020040";
        ram_buffer(15543) := X"8FA50048";
        ram_buffer(15544) := X"8E040038";
        ram_buffer(15545) := X"00A20018";
        ram_buffer(15546) := X"00001012";
        ram_buffer(15547) := X"188000AD";
        ram_buffer(15548) := X"AFA20020";
        ram_buffer(15549) := X"26C20001";
        ram_buffer(15550) := X"AFA2002C";
        ram_buffer(15551) := X"26C20002";
        ram_buffer(15552) := X"AFA20030";
        ram_buffer(15553) := X"26C20003";
        ram_buffer(15554) := X"AFA20034";
        ram_buffer(15555) := X"26C20004";
        ram_buffer(15556) := X"8FB20050";
        ram_buffer(15557) := X"0000F021";
        ram_buffer(15558) := X"AFA20038";
        ram_buffer(15559) := X"26C20005";
        ram_buffer(15560) := X"02A01821";
        ram_buffer(15561) := X"AFA2003C";
        ram_buffer(15562) := X"03C01021";
        ram_buffer(15563) := X"02C0A821";
        ram_buffer(15564) := X"0200F021";
        ram_buffer(15565) := X"0280B021";
        ram_buffer(15566) := X"00408021";
        ram_buffer(15567) := X"0240A021";
        ram_buffer(15568) := X"10000007";
        ram_buffer(15569) := X"00609021";
        ram_buffer(15570) := X"8FC30038";
        ram_buffer(15571) := X"26100001";
        ram_buffer(15572) := X"0203182A";
        ram_buffer(15573) := X"02459021";
        ram_buffer(15574) := X"1060008F";
        ram_buffer(15575) := X"26940008";
        ram_buffer(15576) := X"8EC30008";
        ram_buffer(15577) := X"00000000";
        ram_buffer(15578) := X"0073182B";
        ram_buffer(15579) := X"14600007";
        ram_buffer(15580) := X"26430006";
        ram_buffer(15581) := X"8FA20024";
        ram_buffer(15582) := X"8FC30048";
        ram_buffer(15583) := X"02022021";
        ram_buffer(15584) := X"0083182A";
        ram_buffer(15585) := X"106000AE";
        ram_buffer(15586) := X"26430006";
        ram_buffer(15587) := X"8FA20020";
        ram_buffer(15588) := X"00031880";
        ram_buffer(15589) := X"8EE40160";
        ram_buffer(15590) := X"02C31821";
        ram_buffer(15591) := X"8C670000";
        ram_buffer(15592) := X"8E260000";
        ram_buffer(15593) := X"AFB50018";
        ram_buffer(15594) := X"AFA20014";
        ram_buffer(15595) := X"AFB40010";
        ram_buffer(15596) := X"8C830004";
        ram_buffer(15597) := X"03C02821";
        ram_buffer(15598) := X"0060F809";
        ram_buffer(15599) := X"02E02021";
        ram_buffer(15600) := X"8FC50034";
        ram_buffer(15601) := X"00000000";
        ram_buffer(15602) := X"02A5182A";
        ram_buffer(15603) := X"1060FFDE";
        ram_buffer(15604) := X"02B21821";
        ram_buffer(15605) := X"00031880";
        ram_buffer(15606) := X"02C31821";
        ram_buffer(15607) := X"8C640018";
        ram_buffer(15608) := X"00B52823";
        ram_buffer(15609) := X"000529C0";
        ram_buffer(15610) := X"0C0264DD";
        ram_buffer(15611) := X"AFA30028";
        ram_buffer(15612) := X"8FC50034";
        ram_buffer(15613) := X"00000000";
        ram_buffer(15614) := X"02A5202A";
        ram_buffer(15615) := X"1080FFD2";
        ram_buffer(15616) := X"00000000";
        ram_buffer(15617) := X"8FA30028";
        ram_buffer(15618) := X"8FA2002C";
        ram_buffer(15619) := X"8C660014";
        ram_buffer(15620) := X"8C640018";
        ram_buffer(15621) := X"84C60000";
        ram_buffer(15622) := X"0045182A";
        ram_buffer(15623) := X"1060FFCA";
        ram_buffer(15624) := X"A4860000";
        ram_buffer(15625) := X"00521821";
        ram_buffer(15626) := X"00031880";
        ram_buffer(15627) := X"02C31821";
        ram_buffer(15628) := X"8C660014";
        ram_buffer(15629) := X"8FA20030";
        ram_buffer(15630) := X"8C640018";
        ram_buffer(15631) := X"84C60000";
        ram_buffer(15632) := X"0045182A";
        ram_buffer(15633) := X"1060FFC0";
        ram_buffer(15634) := X"A4860000";
        ram_buffer(15635) := X"00521821";
        ram_buffer(15636) := X"00031880";
        ram_buffer(15637) := X"02C31821";
        ram_buffer(15638) := X"8C660014";
        ram_buffer(15639) := X"8FA20034";
        ram_buffer(15640) := X"8C640018";
        ram_buffer(15641) := X"84C60000";
        ram_buffer(15642) := X"0045182A";
        ram_buffer(15643) := X"1060FFB6";
        ram_buffer(15644) := X"A4860000";
        ram_buffer(15645) := X"00521821";
        ram_buffer(15646) := X"00031880";
        ram_buffer(15647) := X"02C31821";
        ram_buffer(15648) := X"8C660014";
        ram_buffer(15649) := X"8FA20038";
        ram_buffer(15650) := X"8C640018";
        ram_buffer(15651) := X"84C60000";
        ram_buffer(15652) := X"0045182A";
        ram_buffer(15653) := X"1060FFAC";
        ram_buffer(15654) := X"A4860000";
        ram_buffer(15655) := X"00521821";
        ram_buffer(15656) := X"00031880";
        ram_buffer(15657) := X"02C31821";
        ram_buffer(15658) := X"8C660014";
        ram_buffer(15659) := X"8FA2003C";
        ram_buffer(15660) := X"8C640018";
        ram_buffer(15661) := X"84C60000";
        ram_buffer(15662) := X"0045182A";
        ram_buffer(15663) := X"1060FFA2";
        ram_buffer(15664) := X"A4860000";
        ram_buffer(15665) := X"00521821";
        ram_buffer(15666) := X"00031880";
        ram_buffer(15667) := X"02C31821";
        ram_buffer(15668) := X"8C640014";
        ram_buffer(15669) := X"8C660018";
        ram_buffer(15670) := X"84870000";
        ram_buffer(15671) := X"26A30006";
        ram_buffer(15672) := X"0065202A";
        ram_buffer(15673) := X"1080FF98";
        ram_buffer(15674) := X"A4C70000";
        ram_buffer(15675) := X"00721821";
        ram_buffer(15676) := X"00031880";
        ram_buffer(15677) := X"02C31821";
        ram_buffer(15678) := X"8C640014";
        ram_buffer(15679) := X"8C660018";
        ram_buffer(15680) := X"84870000";
        ram_buffer(15681) := X"26A30007";
        ram_buffer(15682) := X"0065202A";
        ram_buffer(15683) := X"1080FF8E";
        ram_buffer(15684) := X"A4C70000";
        ram_buffer(15685) := X"00721821";
        ram_buffer(15686) := X"00031880";
        ram_buffer(15687) := X"02C31821";
        ram_buffer(15688) := X"8C640014";
        ram_buffer(15689) := X"8C660018";
        ram_buffer(15690) := X"84870000";
        ram_buffer(15691) := X"26A30008";
        ram_buffer(15692) := X"0065202A";
        ram_buffer(15693) := X"1080FF84";
        ram_buffer(15694) := X"A4C70000";
        ram_buffer(15695) := X"00721821";
        ram_buffer(15696) := X"00031880";
        ram_buffer(15697) := X"02C31821";
        ram_buffer(15698) := X"8C640014";
        ram_buffer(15699) := X"8C660018";
        ram_buffer(15700) := X"84870000";
        ram_buffer(15701) := X"26A30009";
        ram_buffer(15702) := X"0065202A";
        ram_buffer(15703) := X"1080FF7A";
        ram_buffer(15704) := X"A4C70000";
        ram_buffer(15705) := X"00721821";
        ram_buffer(15706) := X"00031880";
        ram_buffer(15707) := X"02C31821";
        ram_buffer(15708) := X"8C640014";
        ram_buffer(15709) := X"8C630018";
        ram_buffer(15710) := X"84840000";
        ram_buffer(15711) := X"26100001";
        ram_buffer(15712) := X"A4640000";
        ram_buffer(15713) := X"8FC30038";
        ram_buffer(15714) := X"02459021";
        ram_buffer(15715) := X"0203182A";
        ram_buffer(15716) := X"1460FF73";
        ram_buffer(15717) := X"26940008";
        ram_buffer(15718) := X"8EE300EC";
        ram_buffer(15719) := X"02C0A021";
        ram_buffer(15720) := X"0240A821";
        ram_buffer(15721) := X"8FA20044";
        ram_buffer(15722) := X"26310004";
        ram_buffer(15723) := X"24420001";
        ram_buffer(15724) := X"AFA20044";
        ram_buffer(15725) := X"0043202A";
        ram_buffer(15726) := X"8FA20040";
        ram_buffer(15727) := X"00000000";
        ram_buffer(15728) := X"24420004";
        ram_buffer(15729) := X"1480FF3E";
        ram_buffer(15730) := X"AFA20040";
        ram_buffer(15731) := X"8EE20164";
        ram_buffer(15732) := X"8FA50058";
        ram_buffer(15733) := X"8C420004";
        ram_buffer(15734) := X"00000000";
        ram_buffer(15735) := X"0040F809";
        ram_buffer(15736) := X"02E02021";
        ram_buffer(15737) := X"1040005C";
        ram_buffer(15738) := X"00000000";
        ram_buffer(15739) := X"8FA20048";
        ram_buffer(15740) := X"8FA30054";
        ram_buffer(15741) := X"24420001";
        ram_buffer(15742) := X"AFA20048";
        ram_buffer(15743) := X"0062102B";
        ram_buffer(15744) := X"1040FF22";
        ram_buffer(15745) := X"0280F021";
        ram_buffer(15746) := X"8E820014";
        ram_buffer(15747) := X"8FA30024";
        ram_buffer(15748) := X"AFC0000C";
        ram_buffer(15749) := X"24630001";
        ram_buffer(15750) := X"AFA30024";
        ram_buffer(15751) := X"0062102A";
        ram_buffer(15752) := X"8FA30050";
        ram_buffer(15753) := X"AFA00048";
        ram_buffer(15754) := X"24630008";
        ram_buffer(15755) := X"1440FF16";
        ram_buffer(15756) := X"AFA30050";
        ram_buffer(15757) := X"8EE20150";
        ram_buffer(15758) := X"1000005A";
        ram_buffer(15759) := X"00000000";
        ram_buffer(15760) := X"00121880";
        ram_buffer(15761) := X"02C31821";
        ram_buffer(15762) := X"8FC50034";
        ram_buffer(15763) := X"8C640018";
        ram_buffer(15764) := X"000529C0";
        ram_buffer(15765) := X"0C0264DD";
        ram_buffer(15766) := X"AFA30028";
        ram_buffer(15767) := X"8FC50034";
        ram_buffer(15768) := X"00000000";
        ram_buffer(15769) := X"18A0FF38";
        ram_buffer(15770) := X"24020001";
        ram_buffer(15771) := X"8FA30028";
        ram_buffer(15772) := X"00000000";
        ram_buffer(15773) := X"8C640014";
        ram_buffer(15774) := X"8C660018";
        ram_buffer(15775) := X"84870000";
        ram_buffer(15776) := X"10A2FF31";
        ram_buffer(15777) := X"A4C70000";
        ram_buffer(15778) := X"84870000";
        ram_buffer(15779) := X"8C66001C";
        ram_buffer(15780) := X"24020002";
        ram_buffer(15781) := X"10A2FF2C";
        ram_buffer(15782) := X"A4C70000";
        ram_buffer(15783) := X"84870000";
        ram_buffer(15784) := X"8C660020";
        ram_buffer(15785) := X"24020003";
        ram_buffer(15786) := X"10A2FF27";
        ram_buffer(15787) := X"A4C70000";
        ram_buffer(15788) := X"84870000";
        ram_buffer(15789) := X"8C660024";
        ram_buffer(15790) := X"24020004";
        ram_buffer(15791) := X"10A2FF22";
        ram_buffer(15792) := X"A4C70000";
        ram_buffer(15793) := X"84870000";
        ram_buffer(15794) := X"8C660028";
        ram_buffer(15795) := X"24020005";
        ram_buffer(15796) := X"10A2FF1D";
        ram_buffer(15797) := X"A4C70000";
        ram_buffer(15798) := X"8C66002C";
        ram_buffer(15799) := X"84870000";
        ram_buffer(15800) := X"00000000";
        ram_buffer(15801) := X"A4C70000";
        ram_buffer(15802) := X"24060006";
        ram_buffer(15803) := X"10A6FF16";
        ram_buffer(15804) := X"00000000";
        ram_buffer(15805) := X"8C660030";
        ram_buffer(15806) := X"84870000";
        ram_buffer(15807) := X"00000000";
        ram_buffer(15808) := X"A4C70000";
        ram_buffer(15809) := X"24060007";
        ram_buffer(15810) := X"10A6FF0F";
        ram_buffer(15811) := X"00000000";
        ram_buffer(15812) := X"8C660034";
        ram_buffer(15813) := X"84870000";
        ram_buffer(15814) := X"00000000";
        ram_buffer(15815) := X"A4C70000";
        ram_buffer(15816) := X"24060008";
        ram_buffer(15817) := X"10A6FF08";
        ram_buffer(15818) := X"00000000";
        ram_buffer(15819) := X"8C660038";
        ram_buffer(15820) := X"84870000";
        ram_buffer(15821) := X"00000000";
        ram_buffer(15822) := X"A4C70000";
        ram_buffer(15823) := X"24060009";
        ram_buffer(15824) := X"10A6FF01";
        ram_buffer(15825) := X"00000000";
        ram_buffer(15826) := X"84840000";
        ram_buffer(15827) := X"8C63003C";
        ram_buffer(15828) := X"1000FEFD";
        ram_buffer(15829) := X"A4640000";
        ram_buffer(15830) := X"8FA30024";
        ram_buffer(15831) := X"00000000";
        ram_buffer(15832) := X"AE830010";
        ram_buffer(15833) := X"8FA30048";
        ram_buffer(15834) := X"00000000";
        ram_buffer(15835) := X"AE83000C";
        ram_buffer(15836) := X"8FBF0084";
        ram_buffer(15837) := X"8FBE0080";
        ram_buffer(15838) := X"8FB7007C";
        ram_buffer(15839) := X"8FB60078";
        ram_buffer(15840) := X"8FB50074";
        ram_buffer(15841) := X"8FB40070";
        ram_buffer(15842) := X"8FB3006C";
        ram_buffer(15843) := X"8FB20068";
        ram_buffer(15844) := X"8FB10064";
        ram_buffer(15845) := X"8FB00060";
        ram_buffer(15846) := X"03E00008";
        ram_buffer(15847) := X"27BD0088";
        ram_buffer(15848) := X"03C01021";
        ram_buffer(15849) := X"8FC40008";
        ram_buffer(15850) := X"8EE300EC";
        ram_buffer(15851) := X"24840001";
        ram_buffer(15852) := X"28630002";
        ram_buffer(15853) := X"1460000A";
        ram_buffer(15854) := X"AFC40008";
        ram_buffer(15855) := X"24030001";
        ram_buffer(15856) := X"AC430014";
        ram_buffer(15857) := X"AC40000C";
        ram_buffer(15858) := X"AC400010";
        ram_buffer(15859) := X"1000FFE8";
        ram_buffer(15860) := X"24020001";
        ram_buffer(15861) := X"8E160044";
        ram_buffer(15862) := X"1000FEBF";
        ram_buffer(15863) := X"00000000";
        ram_buffer(15864) := X"8EE400E8";
        ram_buffer(15865) := X"8C430008";
        ram_buffer(15866) := X"2484FFFF";
        ram_buffer(15867) := X"0064182B";
        ram_buffer(15868) := X"10600006";
        ram_buffer(15869) := X"00000000";
        ram_buffer(15870) := X"8EE300F0";
        ram_buffer(15871) := X"00000000";
        ram_buffer(15872) := X"8C63000C";
        ram_buffer(15873) := X"1000FFEF";
        ram_buffer(15874) := X"AC430014";
        ram_buffer(15875) := X"8EE300F0";
        ram_buffer(15876) := X"00000000";
        ram_buffer(15877) := X"8C630048";
        ram_buffer(15878) := X"1000FFEA";
        ram_buffer(15879) := X"AC430014";
        ram_buffer(15880) := X"8C820004";
        ram_buffer(15881) := X"27BDFFC8";
        ram_buffer(15882) := X"8C420000";
        ram_buffer(15883) := X"24060068";
        ram_buffer(15884) := X"AFB20024";
        ram_buffer(15885) := X"AFB10020";
        ram_buffer(15886) := X"AFB0001C";
        ram_buffer(15887) := X"AFBF0034";
        ram_buffer(15888) := X"AFB50030";
        ram_buffer(15889) := X"AFB4002C";
        ram_buffer(15890) := X"AFB30028";
        ram_buffer(15891) := X"00A08021";
        ram_buffer(15892) := X"24050001";
        ram_buffer(15893) := X"0040F809";
        ram_buffer(15894) := X"00809021";
        ram_buffer(15895) := X"00408821";
        ram_buffer(15896) := X"AE420150";
        ram_buffer(15897) := X"3C021009";
        ram_buffer(15898) := X"2442E6F0";
        ram_buffer(15899) := X"12000028";
        ram_buffer(15900) := X"AE220000";
        ram_buffer(15901) := X"8E420034";
        ram_buffer(15902) := X"8E50003C";
        ram_buffer(15903) := X"1840001B";
        ram_buffer(15904) := X"26310040";
        ram_buffer(15905) := X"00009821";
        ram_buffer(15906) := X"8E050008";
        ram_buffer(15907) := X"8E04001C";
        ram_buffer(15908) := X"8E420004";
        ram_buffer(15909) := X"00000000";
        ram_buffer(15910) := X"8C540014";
        ram_buffer(15911) := X"0C0264B3";
        ram_buffer(15912) := X"26730001";
        ram_buffer(15913) := X"8E05000C";
        ram_buffer(15914) := X"8E040020";
        ram_buffer(15915) := X"0C0264B3";
        ram_buffer(15916) := X"0040A821";
        ram_buffer(15917) := X"8E03000C";
        ram_buffer(15918) := X"02A03821";
        ram_buffer(15919) := X"AFA30014";
        ram_buffer(15920) := X"AFA20010";
        ram_buffer(15921) := X"00003021";
        ram_buffer(15922) := X"24050001";
        ram_buffer(15923) := X"0280F809";
        ram_buffer(15924) := X"02402021";
        ram_buffer(15925) := X"8E430034";
        ram_buffer(15926) := X"26100054";
        ram_buffer(15927) := X"0263182A";
        ram_buffer(15928) := X"AE220000";
        ram_buffer(15929) := X"1460FFE8";
        ram_buffer(15930) := X"26310004";
        ram_buffer(15931) := X"8FBF0034";
        ram_buffer(15932) := X"8FB50030";
        ram_buffer(15933) := X"8FB4002C";
        ram_buffer(15934) := X"8FB30028";
        ram_buffer(15935) := X"8FB20024";
        ram_buffer(15936) := X"8FB10020";
        ram_buffer(15937) := X"8FB0001C";
        ram_buffer(15938) := X"03E00008";
        ram_buffer(15939) := X"27BD0038";
        ram_buffer(15940) := X"8E420004";
        ram_buffer(15941) := X"24060500";
        ram_buffer(15942) := X"8C420004";
        ram_buffer(15943) := X"24050001";
        ram_buffer(15944) := X"0040F809";
        ram_buffer(15945) := X"02402021";
        ram_buffer(15946) := X"244B0080";
        ram_buffer(15947) := X"244A0100";
        ram_buffer(15948) := X"24490180";
        ram_buffer(15949) := X"24480200";
        ram_buffer(15950) := X"24470280";
        ram_buffer(15951) := X"24460300";
        ram_buffer(15952) := X"24450380";
        ram_buffer(15953) := X"24440400";
        ram_buffer(15954) := X"24430480";
        ram_buffer(15955) := X"AE220018";
        ram_buffer(15956) := X"AE2B001C";
        ram_buffer(15957) := X"AE2A0020";
        ram_buffer(15958) := X"AE290024";
        ram_buffer(15959) := X"AE280028";
        ram_buffer(15960) := X"AE27002C";
        ram_buffer(15961) := X"AE260030";
        ram_buffer(15962) := X"AE250034";
        ram_buffer(15963) := X"AE240038";
        ram_buffer(15964) := X"AE23003C";
        ram_buffer(15965) := X"1000FFDD";
        ram_buffer(15966) := X"AE200040";
        ram_buffer(15967) := X"8C830004";
        ram_buffer(15968) := X"27BDFFE8";
        ram_buffer(15969) := X"8C620000";
        ram_buffer(15970) := X"24062000";
        ram_buffer(15971) := X"AFB00010";
        ram_buffer(15972) := X"8C900158";
        ram_buffer(15973) := X"AFBF0014";
        ram_buffer(15974) := X"0040F809";
        ram_buffer(15975) := X"24050001";
        ram_buffer(15976) := X"3C040080";
        ram_buffer(15977) := X"3C0B004C";
        ram_buffer(15978) := X"AE020008";
        ram_buffer(15979) := X"00005021";
        ram_buffer(15980) := X"00004821";
        ram_buffer(15981) := X"24847FFF";
        ram_buffer(15982) := X"00004021";
        ram_buffer(15983) := X"00003821";
        ram_buffer(15984) := X"34068000";
        ram_buffer(15985) := X"00002821";
        ram_buffer(15986) := X"00001821";
        ram_buffer(15987) := X"340D9646";
        ram_buffer(15988) := X"340C8000";
        ram_buffer(15989) := X"356B8B00";
        ram_buffer(15990) := X"AC430000";
        ram_buffer(15991) := X"24634C8B";
        ram_buffer(15992) := X"AC450400";
        ram_buffer(15993) := X"AC460800";
        ram_buffer(15994) := X"AC470C00";
        ram_buffer(15995) := X"AC481000";
        ram_buffer(15996) := X"AC441400";
        ram_buffer(15997) := X"AC491800";
        ram_buffer(15998) := X"AC4A1C00";
        ram_buffer(15999) := X"00AD2821";
        ram_buffer(16000) := X"24420004";
        ram_buffer(16001) := X"24C61D2F";
        ram_buffer(16002) := X"24E7D4CD";
        ram_buffer(16003) := X"2508AB33";
        ram_buffer(16004) := X"008C2021";
        ram_buffer(16005) := X"252994D1";
        ram_buffer(16006) := X"146BFFEF";
        ram_buffer(16007) := X"254AEB2F";
        ram_buffer(16008) := X"8FBF0014";
        ram_buffer(16009) := X"8FB00010";
        ram_buffer(16010) := X"03E00008";
        ram_buffer(16011) := X"27BD0018";
        ram_buffer(16012) := X"8FAE0010";
        ram_buffer(16013) := X"8C820158";
        ram_buffer(16014) := X"25CEFFFF";
        ram_buffer(16015) := X"8C4C0008";
        ram_buffer(16016) := X"8C8F0018";
        ram_buffer(16017) := X"05C00036";
        ram_buffer(16018) := X"00073880";
        ram_buffer(16019) := X"8CC40000";
        ram_buffer(16020) := X"8CC30004";
        ram_buffer(16021) := X"8CC20008";
        ram_buffer(16022) := X"00872021";
        ram_buffer(16023) := X"8C890000";
        ram_buffer(16024) := X"24A50004";
        ram_buffer(16025) := X"00671821";
        ram_buffer(16026) := X"00471021";
        ram_buffer(16027) := X"8CA8FFFC";
        ram_buffer(16028) := X"8C6B0000";
        ram_buffer(16029) := X"8C4A0000";
        ram_buffer(16030) := X"11E00026";
        ram_buffer(16031) := X"012F6821";
        ram_buffer(16032) := X"91180001";
        ram_buffer(16033) := X"91190000";
        ram_buffer(16034) := X"91020002";
        ram_buffer(16035) := X"27180100";
        ram_buffer(16036) := X"0019C880";
        ram_buffer(16037) := X"0018C080";
        ram_buffer(16038) := X"0199C821";
        ram_buffer(16039) := X"0198C021";
        ram_buffer(16040) := X"24420200";
        ram_buffer(16041) := X"8F240000";
        ram_buffer(16042) := X"8F030000";
        ram_buffer(16043) := X"00021080";
        ram_buffer(16044) := X"01821021";
        ram_buffer(16045) := X"00831821";
        ram_buffer(16046) := X"8C440000";
        ram_buffer(16047) := X"25290001";
        ram_buffer(16048) := X"00641821";
        ram_buffer(16049) := X"00031C03";
        ram_buffer(16050) := X"A123FFFF";
        ram_buffer(16051) := X"8F240C00";
        ram_buffer(16052) := X"8F030C00";
        ram_buffer(16053) := X"25080003";
        ram_buffer(16054) := X"00831821";
        ram_buffer(16055) := X"8C440C00";
        ram_buffer(16056) := X"256B0001";
        ram_buffer(16057) := X"00641821";
        ram_buffer(16058) := X"00031C03";
        ram_buffer(16059) := X"A163FFFF";
        ram_buffer(16060) := X"8F231400";
        ram_buffer(16061) := X"8F181400";
        ram_buffer(16062) := X"8C441400";
        ram_buffer(16063) := X"00781021";
        ram_buffer(16064) := X"00441021";
        ram_buffer(16065) := X"00021403";
        ram_buffer(16066) := X"A1420000";
        ram_buffer(16067) := X"15A9FFDC";
        ram_buffer(16068) := X"254A0001";
        ram_buffer(16069) := X"25CEFFFF";
        ram_buffer(16070) := X"05C1FFCC";
        ram_buffer(16071) := X"24E70004";
        ram_buffer(16072) := X"03E00008";
        ram_buffer(16073) := X"00000000";
        ram_buffer(16074) := X"8FAD0010";
        ram_buffer(16075) := X"8C820158";
        ram_buffer(16076) := X"25ADFFFF";
        ram_buffer(16077) := X"8C4B0008";
        ram_buffer(16078) := X"8C8E0018";
        ram_buffer(16079) := X"05A00020";
        ram_buffer(16080) := X"00073880";
        ram_buffer(16081) := X"8CC20000";
        ram_buffer(16082) := X"24A50004";
        ram_buffer(16083) := X"00471021";
        ram_buffer(16084) := X"8C4A0000";
        ram_buffer(16085) := X"8CA9FFFC";
        ram_buffer(16086) := X"11C00016";
        ram_buffer(16087) := X"014E6021";
        ram_buffer(16088) := X"91220001";
        ram_buffer(16089) := X"91280000";
        ram_buffer(16090) := X"91240002";
        ram_buffer(16091) := X"24420100";
        ram_buffer(16092) := X"00021080";
        ram_buffer(16093) := X"00084080";
        ram_buffer(16094) := X"24840200";
        ram_buffer(16095) := X"01621021";
        ram_buffer(16096) := X"01684021";
        ram_buffer(16097) := X"00042080";
        ram_buffer(16098) := X"8C430000";
        ram_buffer(16099) := X"01642021";
        ram_buffer(16100) := X"8D020000";
        ram_buffer(16101) := X"8C840000";
        ram_buffer(16102) := X"00621021";
        ram_buffer(16103) := X"00441021";
        ram_buffer(16104) := X"00021403";
        ram_buffer(16105) := X"A1420000";
        ram_buffer(16106) := X"254A0001";
        ram_buffer(16107) := X"158AFFEC";
        ram_buffer(16108) := X"25290003";
        ram_buffer(16109) := X"25ADFFFF";
        ram_buffer(16110) := X"05A1FFE2";
        ram_buffer(16111) := X"24E70004";
        ram_buffer(16112) := X"03E00008";
        ram_buffer(16113) := X"00000000";
        ram_buffer(16114) := X"27BDFFF8";
        ram_buffer(16115) := X"8FB80018";
        ram_buffer(16116) := X"8C820158";
        ram_buffer(16117) := X"2718FFFF";
        ram_buffer(16118) := X"AFB10004";
        ram_buffer(16119) := X"AFB00000";
        ram_buffer(16120) := X"8C4E0008";
        ram_buffer(16121) := X"8C990018";
        ram_buffer(16122) := X"00073880";
        ram_buffer(16123) := X"0700003F";
        ram_buffer(16124) := X"240D00FF";
        ram_buffer(16125) := X"8CC90000";
        ram_buffer(16126) := X"8CC2000C";
        ram_buffer(16127) := X"01274821";
        ram_buffer(16128) := X"8CC40004";
        ram_buffer(16129) := X"8CC30008";
        ram_buffer(16130) := X"00471021";
        ram_buffer(16131) := X"8D2C0000";
        ram_buffer(16132) := X"8C490000";
        ram_buffer(16133) := X"24A50004";
        ram_buffer(16134) := X"00872021";
        ram_buffer(16135) := X"00671821";
        ram_buffer(16136) := X"8CA8FFFC";
        ram_buffer(16137) := X"8C8B0000";
        ram_buffer(16138) := X"8C6A0000";
        ram_buffer(16139) := X"1320002C";
        ram_buffer(16140) := X"01397821";
        ram_buffer(16141) := X"91100001";
        ram_buffer(16142) := X"91110000";
        ram_buffer(16143) := X"91020002";
        ram_buffer(16144) := X"01B08023";
        ram_buffer(16145) := X"91030003";
        ram_buffer(16146) := X"01B18823";
        ram_buffer(16147) := X"26100100";
        ram_buffer(16148) := X"01A21023";
        ram_buffer(16149) := X"00118880";
        ram_buffer(16150) := X"00108080";
        ram_buffer(16151) := X"A1230000";
        ram_buffer(16152) := X"01D18821";
        ram_buffer(16153) := X"01D08021";
        ram_buffer(16154) := X"24420200";
        ram_buffer(16155) := X"8E240000";
        ram_buffer(16156) := X"8E030000";
        ram_buffer(16157) := X"00021080";
        ram_buffer(16158) := X"01C21021";
        ram_buffer(16159) := X"00831821";
        ram_buffer(16160) := X"8C440000";
        ram_buffer(16161) := X"25290001";
        ram_buffer(16162) := X"00641821";
        ram_buffer(16163) := X"00031C03";
        ram_buffer(16164) := X"A1830000";
        ram_buffer(16165) := X"8E240C00";
        ram_buffer(16166) := X"8E030C00";
        ram_buffer(16167) := X"25080004";
        ram_buffer(16168) := X"00831821";
        ram_buffer(16169) := X"8C440C00";
        ram_buffer(16170) := X"258C0001";
        ram_buffer(16171) := X"00641821";
        ram_buffer(16172) := X"00031C03";
        ram_buffer(16173) := X"A1630000";
        ram_buffer(16174) := X"8E231400";
        ram_buffer(16175) := X"8E101400";
        ram_buffer(16176) := X"8C441400";
        ram_buffer(16177) := X"00701021";
        ram_buffer(16178) := X"00441021";
        ram_buffer(16179) := X"00021403";
        ram_buffer(16180) := X"A1420000";
        ram_buffer(16181) := X"256B0001";
        ram_buffer(16182) := X"15E9FFD6";
        ram_buffer(16183) := X"254A0001";
        ram_buffer(16184) := X"2718FFFF";
        ram_buffer(16185) := X"0701FFC3";
        ram_buffer(16186) := X"24E70004";
        ram_buffer(16187) := X"8FB10004";
        ram_buffer(16188) := X"8FB00000";
        ram_buffer(16189) := X"03E00008";
        ram_buffer(16190) := X"27BD0008";
        ram_buffer(16191) := X"8FAA0010";
        ram_buffer(16192) := X"8C8B0018";
        ram_buffer(16193) := X"254AFFFF";
        ram_buffer(16194) := X"8C890020";
        ram_buffer(16195) := X"05400010";
        ram_buffer(16196) := X"00073880";
        ram_buffer(16197) := X"8CC20000";
        ram_buffer(16198) := X"24A50004";
        ram_buffer(16199) := X"00471021";
        ram_buffer(16200) := X"8C420000";
        ram_buffer(16201) := X"8CA3FFFC";
        ram_buffer(16202) := X"11600006";
        ram_buffer(16203) := X"004B4021";
        ram_buffer(16204) := X"90640000";
        ram_buffer(16205) := X"24420001";
        ram_buffer(16206) := X"A044FFFF";
        ram_buffer(16207) := X"1502FFFC";
        ram_buffer(16208) := X"00691821";
        ram_buffer(16209) := X"254AFFFF";
        ram_buffer(16210) := X"0541FFF2";
        ram_buffer(16211) := X"24E70004";
        ram_buffer(16212) := X"03E00008";
        ram_buffer(16213) := X"00000000";
        ram_buffer(16214) := X"8FAD0010";
        ram_buffer(16215) := X"8C880034";
        ram_buffer(16216) := X"25ADFFFF";
        ram_buffer(16217) := X"8C8B0018";
        ram_buffer(16218) := X"05A0001B";
        ram_buffer(16219) := X"00077080";
        ram_buffer(16220) := X"01C57023";
        ram_buffer(16221) := X"240FFFFF";
        ram_buffer(16222) := X"19000014";
        ram_buffer(16223) := X"00000000";
        ram_buffer(16224) := X"00AE6021";
        ram_buffer(16225) := X"00C05021";
        ram_buffer(16226) := X"00004821";
        ram_buffer(16227) := X"8D420000";
        ram_buffer(16228) := X"8CA30000";
        ram_buffer(16229) := X"004C1021";
        ram_buffer(16230) := X"8C420000";
        ram_buffer(16231) := X"11600008";
        ram_buffer(16232) := X"00000000";
        ram_buffer(16233) := X"00691821";
        ram_buffer(16234) := X"004B3821";
        ram_buffer(16235) := X"90640000";
        ram_buffer(16236) := X"24420001";
        ram_buffer(16237) := X"A044FFFF";
        ram_buffer(16238) := X"14E2FFFC";
        ram_buffer(16239) := X"00681821";
        ram_buffer(16240) := X"25290001";
        ram_buffer(16241) := X"1509FFF1";
        ram_buffer(16242) := X"254A0004";
        ram_buffer(16243) := X"25ADFFFF";
        ram_buffer(16244) := X"15AFFFE9";
        ram_buffer(16245) := X"24A50004";
        ram_buffer(16246) := X"03E00008";
        ram_buffer(16247) := X"00000000";
        ram_buffer(16248) := X"03E00008";
        ram_buffer(16249) := X"00000000";
        ram_buffer(16250) := X"8C820004";
        ram_buffer(16251) := X"27BDFFE0";
        ram_buffer(16252) := X"8C420000";
        ram_buffer(16253) := X"2406000C";
        ram_buffer(16254) := X"AFB10018";
        ram_buffer(16255) := X"AFB00014";
        ram_buffer(16256) := X"AFBF001C";
        ram_buffer(16257) := X"00808021";
        ram_buffer(16258) := X"0040F809";
        ram_buffer(16259) := X"24050001";
        ram_buffer(16260) := X"8E030024";
        ram_buffer(16261) := X"3C041009";
        ram_buffer(16262) := X"00408821";
        ram_buffer(16263) := X"2484FDE0";
        ram_buffer(16264) := X"2C620006";
        ram_buffer(16265) := X"AE110158";
        ram_buffer(16266) := X"1040002B";
        ram_buffer(16267) := X"AE240000";
        ram_buffer(16268) := X"00032080";
        ram_buffer(16269) := X"3C03100D";
        ram_buffer(16270) := X"24638874";
        ram_buffer(16271) := X"00641821";
        ram_buffer(16272) := X"8C620000";
        ram_buffer(16273) := X"00000000";
        ram_buffer(16274) := X"00400008";
        ram_buffer(16275) := X"00000000";
        ram_buffer(16276) := X"8E030020";
        ram_buffer(16277) := X"24020004";
        ram_buffer(16278) := X"10620007";
        ram_buffer(16279) := X"00000000";
        ram_buffer(16280) := X"8E020000";
        ram_buffer(16281) := X"24040007";
        ram_buffer(16282) := X"8C430000";
        ram_buffer(16283) := X"AC440014";
        ram_buffer(16284) := X"0060F809";
        ram_buffer(16285) := X"02002021";
        ram_buffer(16286) := X"8E020038";
        ram_buffer(16287) := X"00000000";
        ram_buffer(16288) := X"2C430006";
        ram_buffer(16289) := X"10600082";
        ram_buffer(16290) := X"3C04100D";
        ram_buffer(16291) := X"00021880";
        ram_buffer(16292) := X"2484888C";
        ram_buffer(16293) := X"00831821";
        ram_buffer(16294) := X"8C630000";
        ram_buffer(16295) := X"00000000";
        ram_buffer(16296) := X"00600008";
        ram_buffer(16297) := X"00000000";
        ram_buffer(16298) := X"8E030020";
        ram_buffer(16299) := X"24020003";
        ram_buffer(16300) := X"1462FFEB";
        ram_buffer(16301) := X"00000000";
        ram_buffer(16302) := X"1000FFEF";
        ram_buffer(16303) := X"00000000";
        ram_buffer(16304) := X"8E030020";
        ram_buffer(16305) := X"24020001";
        ram_buffer(16306) := X"1462FFE5";
        ram_buffer(16307) := X"00000000";
        ram_buffer(16308) := X"1000FFE9";
        ram_buffer(16309) := X"00000000";
        ram_buffer(16310) := X"8E020020";
        ram_buffer(16311) := X"00000000";
        ram_buffer(16312) := X"1C40FFE5";
        ram_buffer(16313) := X"00000000";
        ram_buffer(16314) := X"1000FFDD";
        ram_buffer(16315) := X"00000000";
        ram_buffer(16316) := X"8E030034";
        ram_buffer(16317) := X"24020004";
        ram_buffer(16318) := X"10620007";
        ram_buffer(16319) := X"00000000";
        ram_buffer(16320) := X"8E020000";
        ram_buffer(16321) := X"24040008";
        ram_buffer(16322) := X"8C430000";
        ram_buffer(16323) := X"AC440014";
        ram_buffer(16324) := X"0060F809";
        ram_buffer(16325) := X"02002021";
        ram_buffer(16326) := X"8E020024";
        ram_buffer(16327) := X"24030004";
        ram_buffer(16328) := X"1043006C";
        ram_buffer(16329) := X"24030005";
        ram_buffer(16330) := X"1043001A";
        ram_buffer(16331) := X"3C021009";
        ram_buffer(16332) := X"8E020000";
        ram_buffer(16333) := X"8FBF001C";
        ram_buffer(16334) := X"8FB10018";
        ram_buffer(16335) := X"8C590000";
        ram_buffer(16336) := X"24030019";
        ram_buffer(16337) := X"02002021";
        ram_buffer(16338) := X"8FB00014";
        ram_buffer(16339) := X"AC430014";
        ram_buffer(16340) := X"03200008";
        ram_buffer(16341) := X"27BD0020";
        ram_buffer(16342) := X"8E030034";
        ram_buffer(16343) := X"24020004";
        ram_buffer(16344) := X"10620007";
        ram_buffer(16345) := X"00000000";
        ram_buffer(16346) := X"8E020000";
        ram_buffer(16347) := X"24040008";
        ram_buffer(16348) := X"8C430000";
        ram_buffer(16349) := X"AC440014";
        ram_buffer(16350) := X"0060F809";
        ram_buffer(16351) := X"02002021";
        ram_buffer(16352) := X"8E030024";
        ram_buffer(16353) := X"24020004";
        ram_buffer(16354) := X"1462FFE9";
        ram_buffer(16355) := X"00000000";
        ram_buffer(16356) := X"3C021009";
        ram_buffer(16357) := X"2442FD58";
        ram_buffer(16358) := X"AE220004";
        ram_buffer(16359) := X"8FBF001C";
        ram_buffer(16360) := X"8FB10018";
        ram_buffer(16361) := X"8FB00014";
        ram_buffer(16362) := X"03E00008";
        ram_buffer(16363) := X"27BD0020";
        ram_buffer(16364) := X"8E030034";
        ram_buffer(16365) := X"24020003";
        ram_buffer(16366) := X"10620007";
        ram_buffer(16367) := X"00000000";
        ram_buffer(16368) := X"8E020000";
        ram_buffer(16369) := X"24040008";
        ram_buffer(16370) := X"8C430000";
        ram_buffer(16371) := X"AC440014";
        ram_buffer(16372) := X"0060F809";
        ram_buffer(16373) := X"02002021";
        ram_buffer(16374) := X"8E020024";
        ram_buffer(16375) := X"24030002";
        ram_buffer(16376) := X"10430043";
        ram_buffer(16377) := X"24030003";
        ram_buffer(16378) := X"1443FFD1";
        ram_buffer(16379) := X"3C021009";
        ram_buffer(16380) := X"1000FFE9";
        ram_buffer(16381) := X"2442FD58";
        ram_buffer(16382) := X"8E030034";
        ram_buffer(16383) := X"24020003";
        ram_buffer(16384) := X"10620007";
        ram_buffer(16385) := X"00000000";
        ram_buffer(16386) := X"8E020000";
        ram_buffer(16387) := X"24040008";
        ram_buffer(16388) := X"8C430000";
        ram_buffer(16389) := X"AC440014";
        ram_buffer(16390) := X"0060F809";
        ram_buffer(16391) := X"02002021";
        ram_buffer(16392) := X"8E030024";
        ram_buffer(16393) := X"24020002";
        ram_buffer(16394) := X"1462FFC1";
        ram_buffer(16395) := X"3C021009";
        ram_buffer(16396) := X"1000FFD9";
        ram_buffer(16397) := X"2442FD58";
        ram_buffer(16398) := X"8E030034";
        ram_buffer(16399) := X"24020001";
        ram_buffer(16400) := X"10620007";
        ram_buffer(16401) := X"00000000";
        ram_buffer(16402) := X"8E020000";
        ram_buffer(16403) := X"24040008";
        ram_buffer(16404) := X"8C430000";
        ram_buffer(16405) := X"AC440014";
        ram_buffer(16406) := X"0060F809";
        ram_buffer(16407) := X"02002021";
        ram_buffer(16408) := X"8E020024";
        ram_buffer(16409) := X"24030001";
        ram_buffer(16410) := X"10430005";
        ram_buffer(16411) := X"24030002";
        ram_buffer(16412) := X"10430026";
        ram_buffer(16413) := X"24030003";
        ram_buffer(16414) := X"1443FFAD";
        ram_buffer(16415) := X"00000000";
        ram_buffer(16416) := X"3C021009";
        ram_buffer(16417) := X"2442FCFC";
        ram_buffer(16418) := X"1000FFC4";
        ram_buffer(16419) := X"AE220004";
        ram_buffer(16420) := X"8E030024";
        ram_buffer(16421) := X"00000000";
        ram_buffer(16422) := X"14430006";
        ram_buffer(16423) := X"00000000";
        ram_buffer(16424) := X"8E030034";
        ram_buffer(16425) := X"8E020020";
        ram_buffer(16426) := X"00000000";
        ram_buffer(16427) := X"1062FFB8";
        ram_buffer(16428) := X"00000000";
        ram_buffer(16429) := X"8E020000";
        ram_buffer(16430) := X"24040019";
        ram_buffer(16431) := X"8C430000";
        ram_buffer(16432) := X"AC440014";
        ram_buffer(16433) := X"0060F809";
        ram_buffer(16434) := X"02002021";
        ram_buffer(16435) := X"1000FFB1";
        ram_buffer(16436) := X"3C021009";
        ram_buffer(16437) := X"3C021009";
        ram_buffer(16438) := X"2442F97C";
        ram_buffer(16439) := X"AE220000";
        ram_buffer(16440) := X"3C021009";
        ram_buffer(16441) := X"2442FBC8";
        ram_buffer(16442) := X"1000FFAC";
        ram_buffer(16443) := X"AE220004";
        ram_buffer(16444) := X"3C021009";
        ram_buffer(16445) := X"2442F97C";
        ram_buffer(16446) := X"AE220000";
        ram_buffer(16447) := X"3C021009";
        ram_buffer(16448) := X"2442FA30";
        ram_buffer(16449) := X"1000FFA5";
        ram_buffer(16450) := X"AE220004";
        ram_buffer(16451) := X"3C021009";
        ram_buffer(16452) := X"2442F97C";
        ram_buffer(16453) := X"AE220000";
        ram_buffer(16454) := X"3C021009";
        ram_buffer(16455) := X"2442FB28";
        ram_buffer(16456) := X"1000FF9E";
        ram_buffer(16457) := X"AE220004";
        ram_buffer(16458) := X"03E00008";
        ram_buffer(16459) := X"00000000";
        ram_buffer(16460) := X"8C820034";
        ram_buffer(16461) := X"27BDFFC8";
        ram_buffer(16462) := X"AFB50028";
        ram_buffer(16463) := X"AFB00014";
        ram_buffer(16464) := X"AFBF0034";
        ram_buffer(16465) := X"AFB70030";
        ram_buffer(16466) := X"AFB6002C";
        ram_buffer(16467) := X"AFB40024";
        ram_buffer(16468) := X"AFB30020";
        ram_buffer(16469) := X"AFB2001C";
        ram_buffer(16470) := X"AFB10018";
        ram_buffer(16471) := X"8C95015C";
        ram_buffer(16472) := X"8C90003C";
        ram_buffer(16473) := X"1840001D";
        ram_buffer(16474) := X"0080B821";
        ram_buffer(16475) := X"8FB40048";
        ram_buffer(16476) := X"00069880";
        ram_buffer(16477) := X"00A09021";
        ram_buffer(16478) := X"00E08821";
        ram_buffer(16479) := X"26B5000C";
        ram_buffer(16480) := X"0000B021";
        ram_buffer(16481) := X"0014A080";
        ram_buffer(16482) := X"8E07000C";
        ram_buffer(16483) := X"8E230000";
        ram_buffer(16484) := X"02870018";
        ram_buffer(16485) := X"8E460000";
        ram_buffer(16486) := X"8EA20000";
        ram_buffer(16487) := X"02002821";
        ram_buffer(16488) := X"00D33021";
        ram_buffer(16489) := X"02E02021";
        ram_buffer(16490) := X"26D60001";
        ram_buffer(16491) := X"26100054";
        ram_buffer(16492) := X"26520004";
        ram_buffer(16493) := X"26310004";
        ram_buffer(16494) := X"26B50004";
        ram_buffer(16495) := X"00003812";
        ram_buffer(16496) := X"0040F809";
        ram_buffer(16497) := X"00673821";
        ram_buffer(16498) := X"8EE20034";
        ram_buffer(16499) := X"00000000";
        ram_buffer(16500) := X"02C2102A";
        ram_buffer(16501) := X"1440FFEC";
        ram_buffer(16502) := X"00000000";
        ram_buffer(16503) := X"8FBF0034";
        ram_buffer(16504) := X"8FB70030";
        ram_buffer(16505) := X"8FB6002C";
        ram_buffer(16506) := X"8FB50028";
        ram_buffer(16507) := X"8FB40024";
        ram_buffer(16508) := X"8FB30020";
        ram_buffer(16509) := X"8FB2001C";
        ram_buffer(16510) := X"8FB10018";
        ram_buffer(16511) := X"8FB00014";
        ram_buffer(16512) := X"03E00008";
        ram_buffer(16513) := X"27BD0038";
        ram_buffer(16514) := X"27BDFFB8";
        ram_buffer(16515) := X"8C8300E0";
        ram_buffer(16516) := X"AFB00020";
        ram_buffer(16517) := X"8CB00008";
        ram_buffer(16518) := X"AFB60038";
        ram_buffer(16519) := X"16000002";
        ram_buffer(16520) := X"0070001A";
        ram_buffer(16521) := X"0007000D";
        ram_buffer(16522) := X"8C9600E4";
        ram_buffer(16523) := X"8CA2000C";
        ram_buffer(16524) := X"AFB3002C";
        ram_buffer(16525) := X"AFB40030";
        ram_buffer(16526) := X"8CB4001C";
        ram_buffer(16527) := X"AFB10024";
        ram_buffer(16528) := X"0014A0C0";
        ram_buffer(16529) := X"8C880018";
        ram_buffer(16530) := X"AFB7003C";
        ram_buffer(16531) := X"AFB20028";
        ram_buffer(16532) := X"AFB50034";
        ram_buffer(16533) := X"AFBF0044";
        ram_buffer(16534) := X"AFBE0040";
        ram_buffer(16535) := X"00A0A821";
        ram_buffer(16536) := X"00C05021";
        ram_buffer(16537) := X"00008012";
        ram_buffer(16538) := X"00000000";
        ram_buffer(16539) := X"00000000";
        ram_buffer(16540) := X"14400002";
        ram_buffer(16541) := X"02C2001A";
        ram_buffer(16542) := X"0007000D";
        ram_buffer(16543) := X"00009812";
        ram_buffer(16544) := X"00000000";
        ram_buffer(16545) := X"00000000";
        ram_buffer(16546) := X"02130018";
        ram_buffer(16547) := X"00008812";
        ram_buffer(16548) := X"001197C2";
        ram_buffer(16549) := X"02519021";
        ram_buffer(16550) := X"02900018";
        ram_buffer(16551) := X"0000B812";
        ram_buffer(16552) := X"02E8B823";
        ram_buffer(16553) := X"1AE00017";
        ram_buffer(16554) := X"00129043";
        ram_buffer(16555) := X"1AC00015";
        ram_buffer(16556) := X"00000000";
        ram_buffer(16557) := X"00C01821";
        ram_buffer(16558) := X"0000F021";
        ram_buffer(16559) := X"8C640000";
        ram_buffer(16560) := X"02E03021";
        ram_buffer(16561) := X"00882021";
        ram_buffer(16562) := X"9085FFFF";
        ram_buffer(16563) := X"AFA7001C";
        ram_buffer(16564) := X"AFAA0018";
        ram_buffer(16565) := X"AFA30014";
        ram_buffer(16566) := X"0C02801D";
        ram_buffer(16567) := X"AFA80010";
        ram_buffer(16568) := X"8FA30014";
        ram_buffer(16569) := X"27DE0001";
        ram_buffer(16570) := X"8FA80010";
        ram_buffer(16571) := X"8FAA0018";
        ram_buffer(16572) := X"8FA7001C";
        ram_buffer(16573) := X"16DEFFF1";
        ram_buffer(16574) := X"24630004";
        ram_buffer(16575) := X"8EA2000C";
        ram_buffer(16576) := X"00000000";
        ram_buffer(16577) := X"18400028";
        ram_buffer(16578) := X"00000000";
        ram_buffer(16579) := X"00E06021";
        ram_buffer(16580) := X"00137080";
        ram_buffer(16581) := X"00006821";
        ram_buffer(16582) := X"8D890000";
        ram_buffer(16583) := X"1280001D";
        ram_buffer(16584) := X"014E4021";
        ram_buffer(16585) := X"01345821";
        ram_buffer(16586) := X"014E4021";
        ram_buffer(16587) := X"00003821";
        ram_buffer(16588) := X"1A60000E";
        ram_buffer(16589) := X"00001821";
        ram_buffer(16590) := X"01403021";
        ram_buffer(16591) := X"00001821";
        ram_buffer(16592) := X"8CC20000";
        ram_buffer(16593) := X"1A000006";
        ram_buffer(16594) := X"00471021";
        ram_buffer(16595) := X"00502821";
        ram_buffer(16596) := X"24420001";
        ram_buffer(16597) := X"9044FFFF";
        ram_buffer(16598) := X"1445FFFD";
        ram_buffer(16599) := X"00641821";
        ram_buffer(16600) := X"24C60004";
        ram_buffer(16601) := X"14C8FFF6";
        ram_buffer(16602) := X"00000000";
        ram_buffer(16603) := X"02431821";
        ram_buffer(16604) := X"16200002";
        ram_buffer(16605) := X"0071001A";
        ram_buffer(16606) := X"0007000D";
        ram_buffer(16607) := X"25290001";
        ram_buffer(16608) := X"00F03821";
        ram_buffer(16609) := X"00001812";
        ram_buffer(16610) := X"152BFFE9";
        ram_buffer(16611) := X"A123FFFF";
        ram_buffer(16612) := X"8EA2000C";
        ram_buffer(16613) := X"25AD0001";
        ram_buffer(16614) := X"01A2182A";
        ram_buffer(16615) := X"258C0004";
        ram_buffer(16616) := X"1460FFDD";
        ram_buffer(16617) := X"01005021";
        ram_buffer(16618) := X"8FBF0044";
        ram_buffer(16619) := X"8FBE0040";
        ram_buffer(16620) := X"8FB7003C";
        ram_buffer(16621) := X"8FB60038";
        ram_buffer(16622) := X"8FB50034";
        ram_buffer(16623) := X"8FB40030";
        ram_buffer(16624) := X"8FB3002C";
        ram_buffer(16625) := X"8FB20028";
        ram_buffer(16626) := X"8FB10024";
        ram_buffer(16627) := X"8FB00020";
        ram_buffer(16628) := X"03E00008";
        ram_buffer(16629) := X"27BD0048";
        ram_buffer(16630) := X"27BDFFC8";
        ram_buffer(16631) := X"AFB3001C";
        ram_buffer(16632) := X"8CB3001C";
        ram_buffer(16633) := X"AFB50024";
        ram_buffer(16634) := X"8C950018";
        ram_buffer(16635) := X"AFB40020";
        ram_buffer(16636) := X"0013A100";
        ram_buffer(16637) := X"0295A023";
        ram_buffer(16638) := X"AFB20018";
        ram_buffer(16639) := X"AFB10014";
        ram_buffer(16640) := X"AFB00010";
        ram_buffer(16641) := X"AFBF0034";
        ram_buffer(16642) := X"AFBE0030";
        ram_buffer(16643) := X"AFB7002C";
        ram_buffer(16644) := X"AFB60028";
        ram_buffer(16645) := X"00A08021";
        ram_buffer(16646) := X"00C08821";
        ram_buffer(16647) := X"00E09021";
        ram_buffer(16648) := X"1A80000F";
        ram_buffer(16649) := X"001398C0";
        ram_buffer(16650) := X"8C9600E4";
        ram_buffer(16651) := X"00000000";
        ram_buffer(16652) := X"1AC0000B";
        ram_buffer(16653) := X"00000000";
        ram_buffer(16654) := X"00C0F021";
        ram_buffer(16655) := X"0000B821";
        ram_buffer(16656) := X"8FC40000";
        ram_buffer(16657) := X"02803021";
        ram_buffer(16658) := X"00952021";
        ram_buffer(16659) := X"9085FFFF";
        ram_buffer(16660) := X"0C02801D";
        ram_buffer(16661) := X"26F70001";
        ram_buffer(16662) := X"16D7FFF9";
        ram_buffer(16663) := X"27DE0004";
        ram_buffer(16664) := X"8E02000C";
        ram_buffer(16665) := X"00000000";
        ram_buffer(16666) := X"1840001A";
        ram_buffer(16667) := X"00000000";
        ram_buffer(16668) := X"02403821";
        ram_buffer(16669) := X"02203021";
        ram_buffer(16670) := X"00005021";
        ram_buffer(16671) := X"8CE30000";
        ram_buffer(16672) := X"8CC40000";
        ram_buffer(16673) := X"1260000E";
        ram_buffer(16674) := X"00000000";
        ram_buffer(16675) := X"00734821";
        ram_buffer(16676) := X"00002821";
        ram_buffer(16677) := X"90820000";
        ram_buffer(16678) := X"90880001";
        ram_buffer(16679) := X"24630001";
        ram_buffer(16680) := X"00481021";
        ram_buffer(16681) := X"00451021";
        ram_buffer(16682) := X"00021043";
        ram_buffer(16683) := X"A062FFFF";
        ram_buffer(16684) := X"38A50001";
        ram_buffer(16685) := X"1469FFF7";
        ram_buffer(16686) := X"24840002";
        ram_buffer(16687) := X"8E02000C";
        ram_buffer(16688) := X"254A0001";
        ram_buffer(16689) := X"0142182A";
        ram_buffer(16690) := X"24E70004";
        ram_buffer(16691) := X"1460FFEB";
        ram_buffer(16692) := X"24C60004";
        ram_buffer(16693) := X"8FBF0034";
        ram_buffer(16694) := X"8FBE0030";
        ram_buffer(16695) := X"8FB7002C";
        ram_buffer(16696) := X"8FB60028";
        ram_buffer(16697) := X"8FB50024";
        ram_buffer(16698) := X"8FB40020";
        ram_buffer(16699) := X"8FB3001C";
        ram_buffer(16700) := X"8FB20018";
        ram_buffer(16701) := X"8FB10014";
        ram_buffer(16702) := X"8FB00010";
        ram_buffer(16703) := X"03E00008";
        ram_buffer(16704) := X"27BD0038";
        ram_buffer(16705) := X"27BDFFC8";
        ram_buffer(16706) := X"AFB20018";
        ram_buffer(16707) := X"8CB2001C";
        ram_buffer(16708) := X"AFB50024";
        ram_buffer(16709) := X"8C950018";
        ram_buffer(16710) := X"AFB40020";
        ram_buffer(16711) := X"0012A100";
        ram_buffer(16712) := X"0295A023";
        ram_buffer(16713) := X"AFB3001C";
        ram_buffer(16714) := X"AFB10014";
        ram_buffer(16715) := X"AFB00010";
        ram_buffer(16716) := X"AFBF0034";
        ram_buffer(16717) := X"AFBE0030";
        ram_buffer(16718) := X"AFB7002C";
        ram_buffer(16719) := X"AFB60028";
        ram_buffer(16720) := X"00A08021";
        ram_buffer(16721) := X"00C08821";
        ram_buffer(16722) := X"00E09821";
        ram_buffer(16723) := X"1A80000F";
        ram_buffer(16724) := X"001290C0";
        ram_buffer(16725) := X"8C9600E4";
        ram_buffer(16726) := X"00000000";
        ram_buffer(16727) := X"1AC0000B";
        ram_buffer(16728) := X"00000000";
        ram_buffer(16729) := X"00C0F021";
        ram_buffer(16730) := X"0000B821";
        ram_buffer(16731) := X"8FC40000";
        ram_buffer(16732) := X"02803021";
        ram_buffer(16733) := X"00952021";
        ram_buffer(16734) := X"9085FFFF";
        ram_buffer(16735) := X"0C02801D";
        ram_buffer(16736) := X"26F70001";
        ram_buffer(16737) := X"16D7FFF9";
        ram_buffer(16738) := X"27DE0004";
        ram_buffer(16739) := X"8E02000C";
        ram_buffer(16740) := X"00000000";
        ram_buffer(16741) := X"18400020";
        ram_buffer(16742) := X"00000000";
        ram_buffer(16743) := X"02603821";
        ram_buffer(16744) := X"02203021";
        ram_buffer(16745) := X"00006821";
        ram_buffer(16746) := X"8CE40000";
        ram_buffer(16747) := X"8CC50000";
        ram_buffer(16748) := X"8CC80004";
        ram_buffer(16749) := X"12400013";
        ram_buffer(16750) := X"00000000";
        ram_buffer(16751) := X"00926021";
        ram_buffer(16752) := X"24090001";
        ram_buffer(16753) := X"90A30000";
        ram_buffer(16754) := X"90AB0001";
        ram_buffer(16755) := X"91020000";
        ram_buffer(16756) := X"910A0001";
        ram_buffer(16757) := X"006B1821";
        ram_buffer(16758) := X"00621021";
        ram_buffer(16759) := X"004A1021";
        ram_buffer(16760) := X"00491021";
        ram_buffer(16761) := X"24840001";
        ram_buffer(16762) := X"00021083";
        ram_buffer(16763) := X"A082FFFF";
        ram_buffer(16764) := X"39290003";
        ram_buffer(16765) := X"24A50002";
        ram_buffer(16766) := X"148CFFF2";
        ram_buffer(16767) := X"25080002";
        ram_buffer(16768) := X"8E02000C";
        ram_buffer(16769) := X"25AD0001";
        ram_buffer(16770) := X"01A2182A";
        ram_buffer(16771) := X"24E70004";
        ram_buffer(16772) := X"1460FFE5";
        ram_buffer(16773) := X"24C60008";
        ram_buffer(16774) := X"8FBF0034";
        ram_buffer(16775) := X"8FBE0030";
        ram_buffer(16776) := X"8FB7002C";
        ram_buffer(16777) := X"8FB60028";
        ram_buffer(16778) := X"8FB50024";
        ram_buffer(16779) := X"8FB40020";
        ram_buffer(16780) := X"8FB3001C";
        ram_buffer(16781) := X"8FB20018";
        ram_buffer(16782) := X"8FB10014";
        ram_buffer(16783) := X"8FB00010";
        ram_buffer(16784) := X"03E00008";
        ram_buffer(16785) := X"27BD0038";
        ram_buffer(16786) := X"27BDFFB0";
        ram_buffer(16787) := X"AFB1002C";
        ram_buffer(16788) := X"8CB1001C";
        ram_buffer(16789) := X"AFB40038";
        ram_buffer(16790) := X"8C940018";
        ram_buffer(16791) := X"AFB00028";
        ram_buffer(16792) := X"00118100";
        ram_buffer(16793) := X"02148023";
        ram_buffer(16794) := X"AFB70044";
        ram_buffer(16795) := X"AFB5003C";
        ram_buffer(16796) := X"AFB20030";
        ram_buffer(16797) := X"AFBF004C";
        ram_buffer(16798) := X"AFBE0048";
        ram_buffer(16799) := X"AFB60040";
        ram_buffer(16800) := X"AFB30034";
        ram_buffer(16801) := X"AFA50054";
        ram_buffer(16802) := X"0080A821";
        ram_buffer(16803) := X"00C0B821";
        ram_buffer(16804) := X"00E09021";
        ram_buffer(16805) := X"1A000010";
        ram_buffer(16806) := X"001188C0";
        ram_buffer(16807) := X"8C9300E4";
        ram_buffer(16808) := X"00000000";
        ram_buffer(16809) := X"2A62FFFF";
        ram_buffer(16810) := X"1440000B";
        ram_buffer(16811) := X"24DEFFFC";
        ram_buffer(16812) := X"26730002";
        ram_buffer(16813) := X"0000B021";
        ram_buffer(16814) := X"8FC40000";
        ram_buffer(16815) := X"02003021";
        ram_buffer(16816) := X"00942021";
        ram_buffer(16817) := X"9085FFFF";
        ram_buffer(16818) := X"0C02801D";
        ram_buffer(16819) := X"26D60001";
        ram_buffer(16820) := X"1676FFF9";
        ram_buffer(16821) := X"27DE0004";
        ram_buffer(16822) := X"8EA200B8";
        ram_buffer(16823) := X"8FA30054";
        ram_buffer(16824) := X"00028100";
        ram_buffer(16825) := X"00023180";
        ram_buffer(16826) := X"02063021";
        ram_buffer(16827) := X"8C63000C";
        ram_buffer(16828) := X"00063023";
        ram_buffer(16829) := X"186000A7";
        ram_buffer(16830) := X"24C64000";
        ram_buffer(16831) := X"2623FFFE";
        ram_buffer(16832) := X"00111040";
        ram_buffer(16833) := X"AFA3001C";
        ram_buffer(16834) := X"2442FFFC";
        ram_buffer(16835) := X"2623FFFF";
        ram_buffer(16836) := X"AFA00010";
        ram_buffer(16837) := X"AFA30020";
        ram_buffer(16838) := X"34158000";
        ram_buffer(16839) := X"0240F021";
        ram_buffer(16840) := X"0040B021";
        ram_buffer(16841) := X"8EF3FFFC";
        ram_buffer(16842) := X"8EF10008";
        ram_buffer(16843) := X"926A0000";
        ram_buffer(16844) := X"92640001";
        ram_buffer(16845) := X"92280000";
        ram_buffer(16846) := X"8EF20000";
        ram_buffer(16847) := X"92220001";
        ram_buffer(16848) := X"008A2021";
        ram_buffer(16849) := X"8EE50004";
        ram_buffer(16850) := X"92490000";
        ram_buffer(16851) := X"00882021";
        ram_buffer(16852) := X"92470001";
        ram_buffer(16853) := X"92430002";
        ram_buffer(16854) := X"00822021";
        ram_buffer(16855) := X"90AB0000";
        ram_buffer(16856) := X"00892021";
        ram_buffer(16857) := X"90AE0001";
        ram_buffer(16858) := X"00831821";
        ram_buffer(16859) := X"00E92021";
        ram_buffer(16860) := X"008B2021";
        ram_buffer(16861) := X"008E2021";
        ram_buffer(16862) := X"00860018";
        ram_buffer(16863) := X"926D0002";
        ram_buffer(16864) := X"90A20002";
        ram_buffer(16865) := X"922C0002";
        ram_buffer(16866) := X"01AA5021";
        ram_buffer(16867) := X"006B1821";
        ram_buffer(16868) := X"00621821";
        ram_buffer(16869) := X"01481021";
        ram_buffer(16870) := X"00031840";
        ram_buffer(16871) := X"004C1021";
        ram_buffer(16872) := X"00431021";
        ram_buffer(16873) := X"8FC40000";
        ram_buffer(16874) := X"00001812";
        ram_buffer(16875) := X"8FA80020";
        ram_buffer(16876) := X"24870001";
        ram_buffer(16877) := X"00500018";
        ram_buffer(16878) := X"24A50002";
        ram_buffer(16879) := X"26520002";
        ram_buffer(16880) := X"26730002";
        ram_buffer(16881) := X"26310002";
        ram_buffer(16882) := X"AFA70014";
        ram_buffer(16883) := X"AFA50018";
        ram_buffer(16884) := X"0088A021";
        ram_buffer(16885) := X"00E0C821";
        ram_buffer(16886) := X"0220C021";
        ram_buffer(16887) := X"02607821";
        ram_buffer(16888) := X"00A07021";
        ram_buffer(16889) := X"00001012";
        ram_buffer(16890) := X"00431821";
        ram_buffer(16891) := X"00751821";
        ram_buffer(16892) := X"00031C03";
        ram_buffer(16893) := X"02406821";
        ram_buffer(16894) := X"A0830000";
        ram_buffer(16895) := X"91E70001";
        ram_buffer(16896) := X"91E30000";
        ram_buffer(16897) := X"93020000";
        ram_buffer(16898) := X"93040001";
        ram_buffer(16899) := X"00671821";
        ram_buffer(16900) := X"00621021";
        ram_buffer(16901) := X"91A7FFFF";
        ram_buffer(16902) := X"91A90002";
        ram_buffer(16903) := X"00441021";
        ram_buffer(16904) := X"91E50002";
        ram_buffer(16905) := X"91CCFFFF";
        ram_buffer(16906) := X"91E4FFFF";
        ram_buffer(16907) := X"91A80000";
        ram_buffer(16908) := X"91AB0001";
        ram_buffer(16909) := X"00473821";
        ram_buffer(16910) := X"91CA0000";
        ram_buffer(16911) := X"91C20002";
        ram_buffer(16912) := X"00E93821";
        ram_buffer(16913) := X"00852021";
        ram_buffer(16914) := X"00EC3821";
        ram_buffer(16915) := X"91C50001";
        ram_buffer(16916) := X"010B4021";
        ram_buffer(16917) := X"00E23821";
        ram_buffer(16918) := X"010A1021";
        ram_buffer(16919) := X"00451021";
        ram_buffer(16920) := X"00460018";
        ram_buffer(16921) := X"9303FFFF";
        ram_buffer(16922) := X"93090002";
        ram_buffer(16923) := X"00832021";
        ram_buffer(16924) := X"00073840";
        ram_buffer(16925) := X"00891821";
        ram_buffer(16926) := X"00671821";
        ram_buffer(16927) := X"27390001";
        ram_buffer(16928) := X"25AD0002";
        ram_buffer(16929) := X"25CE0002";
        ram_buffer(16930) := X"25EF0002";
        ram_buffer(16931) := X"27180002";
        ram_buffer(16932) := X"00001012";
        ram_buffer(16933) := X"00000000";
        ram_buffer(16934) := X"00000000";
        ram_buffer(16935) := X"00700018";
        ram_buffer(16936) := X"00001812";
        ram_buffer(16937) := X"00621021";
        ram_buffer(16938) := X"00551021";
        ram_buffer(16939) := X"00021403";
        ram_buffer(16940) := X"1734FFD2";
        ram_buffer(16941) := X"A322FFFF";
        ram_buffer(16942) := X"02769821";
        ram_buffer(16943) := X"02368821";
        ram_buffer(16944) := X"92640001";
        ram_buffer(16945) := X"92680000";
        ram_buffer(16946) := X"92220000";
        ram_buffer(16947) := X"02569021";
        ram_buffer(16948) := X"92290001";
        ram_buffer(16949) := X"01044021";
        ram_buffer(16950) := X"9247FFFF";
        ram_buffer(16951) := X"01024021";
        ram_buffer(16952) := X"8FA20018";
        ram_buffer(16953) := X"01094021";
        ram_buffer(16954) := X"00565021";
        ram_buffer(16955) := X"924B0001";
        ram_buffer(16956) := X"01073821";
        ram_buffer(16957) := X"92480000";
        ram_buffer(16958) := X"91420001";
        ram_buffer(16959) := X"914CFFFF";
        ram_buffer(16960) := X"914A0000";
        ram_buffer(16961) := X"9265FFFF";
        ram_buffer(16962) := X"00EB3821";
        ram_buffer(16963) := X"010B4021";
        ram_buffer(16964) := X"00EC3821";
        ram_buffer(16965) := X"010A5021";
        ram_buffer(16966) := X"00A42021";
        ram_buffer(16967) := X"00E22821";
        ram_buffer(16968) := X"01421021";
        ram_buffer(16969) := X"00460018";
        ram_buffer(16970) := X"9223FFFF";
        ram_buffer(16971) := X"00052840";
        ram_buffer(16972) := X"00832021";
        ram_buffer(16973) := X"00891821";
        ram_buffer(16974) := X"00651821";
        ram_buffer(16975) := X"8FA40014";
        ram_buffer(16976) := X"8FA5001C";
        ram_buffer(16977) := X"27DE0004";
        ram_buffer(16978) := X"00852021";
        ram_buffer(16979) := X"8FA50010";
        ram_buffer(16980) := X"00001012";
        ram_buffer(16981) := X"24A50001";
        ram_buffer(16982) := X"AFA50010";
        ram_buffer(16983) := X"00700018";
        ram_buffer(16984) := X"00001812";
        ram_buffer(16985) := X"00621021";
        ram_buffer(16986) := X"34038000";
        ram_buffer(16987) := X"00431021";
        ram_buffer(16988) := X"00021403";
        ram_buffer(16989) := X"A0820000";
        ram_buffer(16990) := X"8FA20054";
        ram_buffer(16991) := X"00000000";
        ram_buffer(16992) := X"8C42000C";
        ram_buffer(16993) := X"00000000";
        ram_buffer(16994) := X"00A2102A";
        ram_buffer(16995) := X"1440FF65";
        ram_buffer(16996) := X"26F70008";
        ram_buffer(16997) := X"8FBF004C";
        ram_buffer(16998) := X"8FBE0048";
        ram_buffer(16999) := X"8FB70044";
        ram_buffer(17000) := X"8FB60040";
        ram_buffer(17001) := X"8FB5003C";
        ram_buffer(17002) := X"8FB40038";
        ram_buffer(17003) := X"8FB30034";
        ram_buffer(17004) := X"8FB20030";
        ram_buffer(17005) := X"8FB1002C";
        ram_buffer(17006) := X"8FB00028";
        ram_buffer(17007) := X"03E00008";
        ram_buffer(17008) := X"27BD0050";
        ram_buffer(17009) := X"27BDFFC8";
        ram_buffer(17010) := X"AFB3001C";
        ram_buffer(17011) := X"8CB3001C";
        ram_buffer(17012) := X"AFB20018";
        ram_buffer(17013) := X"8C920018";
        ram_buffer(17014) := X"001398C0";
        ram_buffer(17015) := X"AFB60028";
        ram_buffer(17016) := X"0272B023";
        ram_buffer(17017) := X"AFB7002C";
        ram_buffer(17018) := X"AFB40020";
        ram_buffer(17019) := X"AFB00010";
        ram_buffer(17020) := X"AFBF0034";
        ram_buffer(17021) := X"AFBE0030";
        ram_buffer(17022) := X"AFB50024";
        ram_buffer(17023) := X"AFB10014";
        ram_buffer(17024) := X"00A08021";
        ram_buffer(17025) := X"0080B821";
        ram_buffer(17026) := X"00C0A021";
        ram_buffer(17027) := X"1AC00010";
        ram_buffer(17028) := X"AFA70044";
        ram_buffer(17029) := X"8C9100E4";
        ram_buffer(17030) := X"00000000";
        ram_buffer(17031) := X"2A22FFFF";
        ram_buffer(17032) := X"1440000B";
        ram_buffer(17033) := X"24D5FFFC";
        ram_buffer(17034) := X"26310002";
        ram_buffer(17035) := X"0000F021";
        ram_buffer(17036) := X"8EA40000";
        ram_buffer(17037) := X"02C03021";
        ram_buffer(17038) := X"00922021";
        ram_buffer(17039) := X"9085FFFF";
        ram_buffer(17040) := X"0C02801D";
        ram_buffer(17041) := X"27DE0001";
        ram_buffer(17042) := X"163EFFF9";
        ram_buffer(17043) := X"26B50004";
        ram_buffer(17044) := X"8EEE00B8";
        ram_buffer(17045) := X"240D0080";
        ram_buffer(17046) := X"8E02000C";
        ram_buffer(17047) := X"01AE6823";
        ram_buffer(17048) := X"000D6A40";
        ram_buffer(17049) := X"1840005B";
        ram_buffer(17050) := X"000E7180";
        ram_buffer(17051) := X"8FA70044";
        ram_buffer(17052) := X"2672FFFE";
        ram_buffer(17053) := X"02803021";
        ram_buffer(17054) := X"00008821";
        ram_buffer(17055) := X"2673FFFF";
        ram_buffer(17056) := X"340F8000";
        ram_buffer(17057) := X"34148000";
        ram_buffer(17058) := X"8CCC0004";
        ram_buffer(17059) := X"8CC9FFFC";
        ram_buffer(17060) := X"8CD80000";
        ram_buffer(17061) := X"91830000";
        ram_buffer(17062) := X"91220000";
        ram_buffer(17063) := X"93150000";
        ram_buffer(17064) := X"91240001";
        ram_buffer(17065) := X"91880001";
        ram_buffer(17066) := X"93050001";
        ram_buffer(17067) := X"00431021";
        ram_buffer(17068) := X"00555821";
        ram_buffer(17069) := X"00881821";
        ram_buffer(17070) := X"00654021";
        ram_buffer(17071) := X"004B1021";
        ram_buffer(17072) := X"00481021";
        ram_buffer(17073) := X"004E0018";
        ram_buffer(17074) := X"8CE30000";
        ram_buffer(17075) := X"27180001";
        ram_buffer(17076) := X"24790001";
        ram_buffer(17077) := X"25850001";
        ram_buffer(17078) := X"25290001";
        ram_buffer(17079) := X"01936021";
        ram_buffer(17080) := X"03205021";
        ram_buffer(17081) := X"03002021";
        ram_buffer(17082) := X"00001012";
        ram_buffer(17083) := X"00000000";
        ram_buffer(17084) := X"00000000";
        ram_buffer(17085) := X"01B50018";
        ram_buffer(17086) := X"0000A812";
        ram_buffer(17087) := X"00551021";
        ram_buffer(17088) := X"004F1021";
        ram_buffer(17089) := X"00021403";
        ram_buffer(17090) := X"10000002";
        ram_buffer(17091) := X"A0620000";
        ram_buffer(17092) := X"00604021";
        ram_buffer(17093) := X"24840001";
        ram_buffer(17094) := X"9082FFFF";
        ram_buffer(17095) := X"25290001";
        ram_buffer(17096) := X"01A20018";
        ram_buffer(17097) := X"24A50001";
        ram_buffer(17098) := X"91360000";
        ram_buffer(17099) := X"90A30000";
        ram_buffer(17100) := X"90970000";
        ram_buffer(17101) := X"0102A823";
        ram_buffer(17102) := X"02C31821";
        ram_buffer(17103) := X"02AB5821";
        ram_buffer(17104) := X"00771821";
        ram_buffer(17105) := X"0163A821";
        ram_buffer(17106) := X"254A0001";
        ram_buffer(17107) := X"01005821";
        ram_buffer(17108) := X"00001012";
        ram_buffer(17109) := X"00000000";
        ram_buffer(17110) := X"00000000";
        ram_buffer(17111) := X"02AE0018";
        ram_buffer(17112) := X"0000A812";
        ram_buffer(17113) := X"00551021";
        ram_buffer(17114) := X"004F1021";
        ram_buffer(17115) := X"00021403";
        ram_buffer(17116) := X"14ACFFE7";
        ram_buffer(17117) := X"A142FFFF";
        ram_buffer(17118) := X"0312C021";
        ram_buffer(17119) := X"93020000";
        ram_buffer(17120) := X"0332C821";
        ram_buffer(17121) := X"01A20018";
        ram_buffer(17122) := X"00622023";
        ram_buffer(17123) := X"00884021";
        ram_buffer(17124) := X"01031821";
        ram_buffer(17125) := X"26310001";
        ram_buffer(17126) := X"24E70004";
        ram_buffer(17127) := X"00001012";
        ram_buffer(17128) := X"00000000";
        ram_buffer(17129) := X"00000000";
        ram_buffer(17130) := X"006E0018";
        ram_buffer(17131) := X"00001812";
        ram_buffer(17132) := X"00431021";
        ram_buffer(17133) := X"00541021";
        ram_buffer(17134) := X"00021403";
        ram_buffer(17135) := X"A3220000";
        ram_buffer(17136) := X"8E02000C";
        ram_buffer(17137) := X"00000000";
        ram_buffer(17138) := X"0222102A";
        ram_buffer(17139) := X"1440FFAE";
        ram_buffer(17140) := X"24C60004";
        ram_buffer(17141) := X"8FBF0034";
        ram_buffer(17142) := X"8FBE0030";
        ram_buffer(17143) := X"8FB7002C";
        ram_buffer(17144) := X"8FB60028";
        ram_buffer(17145) := X"8FB50024";
        ram_buffer(17146) := X"8FB40020";
        ram_buffer(17147) := X"8FB3001C";
        ram_buffer(17148) := X"8FB20018";
        ram_buffer(17149) := X"8FB10014";
        ram_buffer(17150) := X"8FB00010";
        ram_buffer(17151) := X"03E00008";
        ram_buffer(17152) := X"27BD0038";
        ram_buffer(17153) := X"27BDFFD0";
        ram_buffer(17154) := X"8C830018";
        ram_buffer(17155) := X"8C8200E4";
        ram_buffer(17156) := X"AFB00018";
        ram_buffer(17157) := X"00E08021";
        ram_buffer(17158) := X"AFB20020";
        ram_buffer(17159) := X"AFB1001C";
        ram_buffer(17160) := X"00A09021";
        ram_buffer(17161) := X"00808821";
        ram_buffer(17162) := X"AFA30014";
        ram_buffer(17163) := X"00C02021";
        ram_buffer(17164) := X"AFA20010";
        ram_buffer(17165) := X"00003821";
        ram_buffer(17166) := X"02003021";
        ram_buffer(17167) := X"00002821";
        ram_buffer(17168) := X"AFB30024";
        ram_buffer(17169) := X"AFBF002C";
        ram_buffer(17170) := X"0C0264BB";
        ram_buffer(17171) := X"AFB40028";
        ram_buffer(17172) := X"8E52001C";
        ram_buffer(17173) := X"8E330018";
        ram_buffer(17174) := X"001290C0";
        ram_buffer(17175) := X"02539023";
        ram_buffer(17176) := X"1A40000D";
        ram_buffer(17177) := X"00000000";
        ram_buffer(17178) := X"8E3400E4";
        ram_buffer(17179) := X"00000000";
        ram_buffer(17180) := X"1A800009";
        ram_buffer(17181) := X"00008821";
        ram_buffer(17182) := X"8E040000";
        ram_buffer(17183) := X"02403021";
        ram_buffer(17184) := X"00932021";
        ram_buffer(17185) := X"9085FFFF";
        ram_buffer(17186) := X"0C02801D";
        ram_buffer(17187) := X"26310001";
        ram_buffer(17188) := X"1691FFF9";
        ram_buffer(17189) := X"26100004";
        ram_buffer(17190) := X"8FBF002C";
        ram_buffer(17191) := X"8FB40028";
        ram_buffer(17192) := X"8FB30024";
        ram_buffer(17193) := X"8FB20020";
        ram_buffer(17194) := X"8FB1001C";
        ram_buffer(17195) := X"8FB00018";
        ram_buffer(17196) := X"03E00008";
        ram_buffer(17197) := X"27BD0030";
        ram_buffer(17198) := X"8C820004";
        ram_buffer(17199) := X"27BDFFC0";
        ram_buffer(17200) := X"8C420000";
        ram_buffer(17201) := X"24060034";
        ram_buffer(17202) := X"AFB70034";
        ram_buffer(17203) := X"AFB00018";
        ram_buffer(17204) := X"AFBF003C";
        ram_buffer(17205) := X"AFBE0038";
        ram_buffer(17206) := X"AFB60030";
        ram_buffer(17207) := X"AFB5002C";
        ram_buffer(17208) := X"AFB40028";
        ram_buffer(17209) := X"AFB30024";
        ram_buffer(17210) := X"AFB20020";
        ram_buffer(17211) := X"AFB1001C";
        ram_buffer(17212) := X"24050001";
        ram_buffer(17213) := X"0040F809";
        ram_buffer(17214) := X"0080B821";
        ram_buffer(17215) := X"00408021";
        ram_buffer(17216) := X"AEE2015C";
        ram_buffer(17217) := X"3C021009";
        ram_buffer(17218) := X"24420128";
        ram_buffer(17219) := X"8EE300B4";
        ram_buffer(17220) := X"AE020000";
        ram_buffer(17221) := X"3C021009";
        ram_buffer(17222) := X"24420130";
        ram_buffer(17223) := X"AE020004";
        ram_buffer(17224) := X"1460008B";
        ram_buffer(17225) := X"AE000008";
        ram_buffer(17226) := X"8EE40034";
        ram_buffer(17227) := X"8EFE003C";
        ram_buffer(17228) := X"18800049";
        ram_buffer(17229) := X"3C021009";
        ram_buffer(17230) := X"3C111009";
        ram_buffer(17231) := X"3C141009";
        ram_buffer(17232) := X"AFA20014";
        ram_buffer(17233) := X"3C131009";
        ram_buffer(17234) := X"3C021009";
        ram_buffer(17235) := X"2615000C";
        ram_buffer(17236) := X"24120001";
        ram_buffer(17237) := X"0000B021";
        ram_buffer(17238) := X"26310208";
        ram_buffer(17239) := X"26940504";
        ram_buffer(17240) := X"267303D8";
        ram_buffer(17241) := X"10000019";
        ram_buffer(17242) := X"AFA20010";
        ram_buffer(17243) := X"1067004F";
        ram_buffer(17244) := X"00000000";
        ram_buffer(17245) := X"14400002";
        ram_buffer(17246) := X"0062001A";
        ram_buffer(17247) := X"0007000D";
        ram_buffer(17248) := X"00001810";
        ram_buffer(17249) := X"14600040";
        ram_buffer(17250) := X"00000000";
        ram_buffer(17251) := X"8EE300E4";
        ram_buffer(17252) := X"8FC2000C";
        ram_buffer(17253) := X"00000000";
        ram_buffer(17254) := X"14400002";
        ram_buffer(17255) := X"0062001A";
        ram_buffer(17256) := X"0007000D";
        ram_buffer(17257) := X"00001810";
        ram_buffer(17258) := X"14600037";
        ram_buffer(17259) := X"00000000";
        ram_buffer(17260) := X"AEB10000";
        ram_buffer(17261) := X"00009021";
        ram_buffer(17262) := X"26D60001";
        ram_buffer(17263) := X"02C4102A";
        ram_buffer(17264) := X"27DE0054";
        ram_buffer(17265) := X"1040001E";
        ram_buffer(17266) := X"26B50004";
        ram_buffer(17267) := X"8FC20008";
        ram_buffer(17268) := X"8EE300E0";
        ram_buffer(17269) := X"00000000";
        ram_buffer(17270) := X"1443FFE4";
        ram_buffer(17271) := X"00023840";
        ram_buffer(17272) := X"8FC7000C";
        ram_buffer(17273) := X"8EE800E4";
        ram_buffer(17274) := X"00000000";
        ram_buffer(17275) := X"10E80037";
        ram_buffer(17276) := X"00024840";
        ram_buffer(17277) := X"1449FFDF";
        ram_buffer(17278) := X"00000000";
        ram_buffer(17279) := X"00073840";
        ram_buffer(17280) := X"14E8FFDC";
        ram_buffer(17281) := X"00000000";
        ram_buffer(17282) := X"8EE200B8";
        ram_buffer(17283) := X"00000000";
        ram_buffer(17284) := X"1040003C";
        ram_buffer(17285) := X"00000000";
        ram_buffer(17286) := X"8FA20014";
        ram_buffer(17287) := X"26D60001";
        ram_buffer(17288) := X"24420648";
        ram_buffer(17289) := X"AEA20000";
        ram_buffer(17290) := X"24020001";
        ram_buffer(17291) := X"AE020008";
        ram_buffer(17292) := X"02C4102A";
        ram_buffer(17293) := X"27DE0054";
        ram_buffer(17294) := X"1440FFE4";
        ram_buffer(17295) := X"26B50004";
        ram_buffer(17296) := X"8EE200B8";
        ram_buffer(17297) := X"00000000";
        ram_buffer(17298) := X"10400003";
        ram_buffer(17299) := X"00000000";
        ram_buffer(17300) := X"1240002E";
        ram_buffer(17301) := X"00002821";
        ram_buffer(17302) := X"8FBF003C";
        ram_buffer(17303) := X"8FBE0038";
        ram_buffer(17304) := X"8FB70034";
        ram_buffer(17305) := X"8FB60030";
        ram_buffer(17306) := X"8FB5002C";
        ram_buffer(17307) := X"8FB40028";
        ram_buffer(17308) := X"8FB30024";
        ram_buffer(17309) := X"8FB20020";
        ram_buffer(17310) := X"8FB1001C";
        ram_buffer(17311) := X"8FB00018";
        ram_buffer(17312) := X"03E00008";
        ram_buffer(17313) := X"27BD0040";
        ram_buffer(17314) := X"8EE20000";
        ram_buffer(17315) := X"24040025";
        ram_buffer(17316) := X"8C430000";
        ram_buffer(17317) := X"AC440014";
        ram_buffer(17318) := X"0060F809";
        ram_buffer(17319) := X"02E02021";
        ram_buffer(17320) := X"8EE40034";
        ram_buffer(17321) := X"1000FFC5";
        ram_buffer(17322) := X"26D60001";
        ram_buffer(17323) := X"8FC7000C";
        ram_buffer(17324) := X"8EE800E4";
        ram_buffer(17325) := X"00000000";
        ram_buffer(17326) := X"14E8FFD0";
        ram_buffer(17327) := X"00000000";
        ram_buffer(17328) := X"AEB30000";
        ram_buffer(17329) := X"1000FFBC";
        ram_buffer(17330) := X"00009021";
        ram_buffer(17331) := X"8EE200B8";
        ram_buffer(17332) := X"00000000";
        ram_buffer(17333) := X"10400006";
        ram_buffer(17334) := X"3C021009";
        ram_buffer(17335) := X"244209C4";
        ram_buffer(17336) := X"AEA20000";
        ram_buffer(17337) := X"24020001";
        ram_buffer(17338) := X"1000FFB3";
        ram_buffer(17339) := X"AE020008";
        ram_buffer(17340) := X"8FA20010";
        ram_buffer(17341) := X"00000000";
        ram_buffer(17342) := X"24420C04";
        ram_buffer(17343) := X"1000FFAE";
        ram_buffer(17344) := X"AEA20000";
        ram_buffer(17345) := X"1000FFAC";
        ram_buffer(17346) := X"AEB40000";
        ram_buffer(17347) := X"8EE20000";
        ram_buffer(17348) := X"8FBF003C";
        ram_buffer(17349) := X"8FBE0038";
        ram_buffer(17350) := X"8FB60030";
        ram_buffer(17351) := X"8FB5002C";
        ram_buffer(17352) := X"8FB40028";
        ram_buffer(17353) := X"8FB30024";
        ram_buffer(17354) := X"8FB20020";
        ram_buffer(17355) := X"8FB1001C";
        ram_buffer(17356) := X"8FB00018";
        ram_buffer(17357) := X"8C590004";
        ram_buffer(17358) := X"24030062";
        ram_buffer(17359) := X"02E02021";
        ram_buffer(17360) := X"8FB70034";
        ram_buffer(17361) := X"AC430014";
        ram_buffer(17362) := X"03200008";
        ram_buffer(17363) := X"27BD0040";
        ram_buffer(17364) := X"8EE20000";
        ram_buffer(17365) := X"24040017";
        ram_buffer(17366) := X"8C430000";
        ram_buffer(17367) := X"AC440014";
        ram_buffer(17368) := X"0060F809";
        ram_buffer(17369) := X"02E02021";
        ram_buffer(17370) := X"1000FF6F";
        ram_buffer(17371) := X"00000000";
        ram_buffer(17372) := X"27BDFFD8";
        ram_buffer(17373) := X"AFB2001C";
        ram_buffer(17374) := X"8C9200C0";
        ram_buffer(17375) := X"AFB30020";
        ram_buffer(17376) := X"AFB10018";
        ram_buffer(17377) := X"AFB00014";
        ram_buffer(17378) := X"AFBF0024";
        ram_buffer(17379) := X"00808821";
        ram_buffer(17380) := X"8C900164";
        ram_buffer(17381) := X"1240000F";
        ram_buffer(17382) := X"00A09821";
        ram_buffer(17383) := X"8E020024";
        ram_buffer(17384) := X"00000000";
        ram_buffer(17385) := X"1440000A";
        ram_buffer(17386) := X"2442FFFF";
        ram_buffer(17387) := X"8C8600EC";
        ram_buffer(17388) := X"00000000";
        ram_buffer(17389) := X"18C00004";
        ram_buffer(17390) := X"00063080";
        ram_buffer(17391) := X"00002821";
        ram_buffer(17392) := X"0C02801D";
        ram_buffer(17393) := X"26040014";
        ram_buffer(17394) := X"02401021";
        ram_buffer(17395) := X"2442FFFF";
        ram_buffer(17396) := X"AE020024";
        ram_buffer(17397) := X"8E220108";
        ram_buffer(17398) := X"00000000";
        ram_buffer(17399) := X"18400059";
        ram_buffer(17400) := X"00021080";
        ram_buffer(17401) := X"3C0F100D";
        ram_buffer(17402) := X"3C09100D";
        ram_buffer(17403) := X"02605821";
        ram_buffer(17404) := X"262D010C";
        ram_buffer(17405) := X"02626021";
        ram_buffer(17406) := X"25EF896C";
        ram_buffer(17407) := X"25298A68";
        ram_buffer(17408) := X"8DA30000";
        ram_buffer(17409) := X"8D680000";
        ram_buffer(17410) := X"2462003C";
        ram_buffer(17411) := X"00021080";
        ram_buffer(17412) := X"02221021";
        ram_buffer(17413) := X"8C420000";
        ram_buffer(17414) := X"00035080";
        ram_buffer(17415) := X"8C440014";
        ram_buffer(17416) := X"8C430018";
        ram_buffer(17417) := X"020A5021";
        ram_buffer(17418) := X"24840012";
        ram_buffer(17419) := X"24630016";
        ram_buffer(17420) := X"850E0000";
        ram_buffer(17421) := X"8D420014";
        ram_buffer(17422) := X"00042080";
        ram_buffer(17423) := X"00031880";
        ram_buffer(17424) := X"02042021";
        ram_buffer(17425) := X"02031821";
        ram_buffer(17426) := X"01C21023";
        ram_buffer(17427) := X"8C840004";
        ram_buffer(17428) := X"8C670004";
        ram_buffer(17429) := X"04400047";
        ram_buffer(17430) := X"00000000";
        ram_buffer(17431) := X"10400005";
        ram_buffer(17432) := X"00001821";
        ram_buffer(17433) := X"00021043";
        ram_buffer(17434) := X"1440FFFE";
        ram_buffer(17435) := X"24630001";
        ram_buffer(17436) := X"00031880";
        ram_buffer(17437) := X"00831821";
        ram_buffer(17438) := X"8C620000";
        ram_buffer(17439) := X"01E02821";
        ram_buffer(17440) := X"24420001";
        ram_buffer(17441) := X"AC620000";
        ram_buffer(17442) := X"00002021";
        ram_buffer(17443) := X"8CA20000";
        ram_buffer(17444) := X"00000000";
        ram_buffer(17445) := X"00021040";
        ram_buffer(17446) := X"01021021";
        ram_buffer(17447) := X"84420000";
        ram_buffer(17448) := X"00000000";
        ram_buffer(17449) := X"1040002F";
        ram_buffer(17450) := X"28830010";
        ram_buffer(17451) := X"14600008";
        ram_buffer(17452) := X"00000000";
        ram_buffer(17453) := X"8CE603C0";
        ram_buffer(17454) := X"2484FFF0";
        ram_buffer(17455) := X"00041902";
        ram_buffer(17456) := X"24C60001";
        ram_buffer(17457) := X"00C33021";
        ram_buffer(17458) := X"3084000F";
        ram_buffer(17459) := X"ACE603C0";
        ram_buffer(17460) := X"04400026";
        ram_buffer(17461) := X"00000000";
        ram_buffer(17462) := X"00021043";
        ram_buffer(17463) := X"10400004";
        ram_buffer(17464) := X"24030001";
        ram_buffer(17465) := X"00021043";
        ram_buffer(17466) := X"1440FFFE";
        ram_buffer(17467) := X"24630001";
        ram_buffer(17468) := X"00042100";
        ram_buffer(17469) := X"00831821";
        ram_buffer(17470) := X"00031880";
        ram_buffer(17471) := X"00E31821";
        ram_buffer(17472) := X"8C620000";
        ram_buffer(17473) := X"00002021";
        ram_buffer(17474) := X"24420001";
        ram_buffer(17475) := X"AC620000";
        ram_buffer(17476) := X"24A50004";
        ram_buffer(17477) := X"1525FFDD";
        ram_buffer(17478) := X"00000000";
        ram_buffer(17479) := X"10800005";
        ram_buffer(17480) := X"00000000";
        ram_buffer(17481) := X"8CE20000";
        ram_buffer(17482) := X"00000000";
        ram_buffer(17483) := X"24420001";
        ram_buffer(17484) := X"ACE20000";
        ram_buffer(17485) := X"256B0004";
        ram_buffer(17486) := X"AD4E0014";
        ram_buffer(17487) := X"158BFFB0";
        ram_buffer(17488) := X"25AD0004";
        ram_buffer(17489) := X"8FBF0024";
        ram_buffer(17490) := X"8FB30020";
        ram_buffer(17491) := X"8FB2001C";
        ram_buffer(17492) := X"8FB10018";
        ram_buffer(17493) := X"8FB00014";
        ram_buffer(17494) := X"24020001";
        ram_buffer(17495) := X"03E00008";
        ram_buffer(17496) := X"27BD0028";
        ram_buffer(17497) := X"1000FFEA";
        ram_buffer(17498) := X"24840001";
        ram_buffer(17499) := X"1000FFDA";
        ram_buffer(17500) := X"00021023";
        ram_buffer(17501) := X"1000FFB9";
        ram_buffer(17502) := X"00021023";
        ram_buffer(17503) := X"27BDFF98";
        ram_buffer(17504) := X"AFB3004C";
        ram_buffer(17505) := X"8C930164";
        ram_buffer(17506) := X"AFB00040";
        ram_buffer(17507) := X"2662000C";
        ram_buffer(17508) := X"8C900014";
        ram_buffer(17509) := X"AFB60058";
        ram_buffer(17510) := X"24060018";
        ram_buffer(17511) := X"0080B021";
        ram_buffer(17512) := X"00402821";
        ram_buffer(17513) := X"AFB7005C";
        ram_buffer(17514) := X"AFB50054";
        ram_buffer(17515) := X"AFB40050";
        ram_buffer(17516) := X"AFB20048";
        ram_buffer(17517) := X"AFB10044";
        ram_buffer(17518) := X"AFBF0064";
        ram_buffer(17519) := X"AFBE0060";
        ram_buffer(17520) := X"AFA20038";
        ram_buffer(17521) := X"8E110000";
        ram_buffer(17522) := X"8E120004";
        ram_buffer(17523) := X"0C027F93";
        ram_buffer(17524) := X"27A40018";
        ram_buffer(17525) := X"8E740010";
        ram_buffer(17526) := X"8E75000C";
        ram_buffer(17527) := X"26970007";
        ram_buffer(17528) := X"24130018";
        ram_buffer(17529) := X"2402007F";
        ram_buffer(17530) := X"02779823";
        ram_buffer(17531) := X"02629804";
        ram_buffer(17532) := X"2AE20008";
        ram_buffer(17533) := X"1440000F";
        ram_buffer(17534) := X"02759825";
        ram_buffer(17535) := X"241E00FF";
        ram_buffer(17536) := X"00131403";
        ram_buffer(17537) := X"2652FFFF";
        ram_buffer(17538) := X"A2220000";
        ram_buffer(17539) := X"305000FF";
        ram_buffer(17540) := X"1240001E";
        ram_buffer(17541) := X"26310001";
        ram_buffer(17542) := X"121E0028";
        ram_buffer(17543) := X"00000000";
        ram_buffer(17544) := X"26F7FFF8";
        ram_buffer(17545) := X"2EE20008";
        ram_buffer(17546) := X"1040FFF5";
        ram_buffer(17547) := X"00139A00";
        ram_buffer(17548) := X"8ED00014";
        ram_buffer(17549) := X"0000A021";
        ram_buffer(17550) := X"0000A821";
        ram_buffer(17551) := X"8FA40038";
        ram_buffer(17552) := X"AE110000";
        ram_buffer(17553) := X"AE120004";
        ram_buffer(17554) := X"27A50018";
        ram_buffer(17555) := X"24060018";
        ram_buffer(17556) := X"AFB50018";
        ram_buffer(17557) := X"0C027F93";
        ram_buffer(17558) := X"AFB4001C";
        ram_buffer(17559) := X"8FBF0064";
        ram_buffer(17560) := X"8FBE0060";
        ram_buffer(17561) := X"8FB7005C";
        ram_buffer(17562) := X"8FB60058";
        ram_buffer(17563) := X"8FB50054";
        ram_buffer(17564) := X"8FB40050";
        ram_buffer(17565) := X"8FB3004C";
        ram_buffer(17566) := X"8FB20048";
        ram_buffer(17567) := X"8FB10044";
        ram_buffer(17568) := X"8FB00040";
        ram_buffer(17569) := X"03E00008";
        ram_buffer(17570) := X"27BD0068";
        ram_buffer(17571) := X"8ED20014";
        ram_buffer(17572) := X"00000000";
        ram_buffer(17573) := X"8E42000C";
        ram_buffer(17574) := X"00000000";
        ram_buffer(17575) := X"0040F809";
        ram_buffer(17576) := X"02C02021";
        ram_buffer(17577) := X"10400015";
        ram_buffer(17578) := X"00000000";
        ram_buffer(17579) := X"8E510000";
        ram_buffer(17580) := X"8E520004";
        ram_buffer(17581) := X"161EFFDA";
        ram_buffer(17582) := X"00000000";
        ram_buffer(17583) := X"2652FFFF";
        ram_buffer(17584) := X"A2200000";
        ram_buffer(17585) := X"1640FFD6";
        ram_buffer(17586) := X"26310001";
        ram_buffer(17587) := X"8ED00014";
        ram_buffer(17588) := X"00000000";
        ram_buffer(17589) := X"8E02000C";
        ram_buffer(17590) := X"00000000";
        ram_buffer(17591) := X"0040F809";
        ram_buffer(17592) := X"02C02021";
        ram_buffer(17593) := X"10400005";
        ram_buffer(17594) := X"26F7FFF8";
        ram_buffer(17595) := X"8E110000";
        ram_buffer(17596) := X"8E120004";
        ram_buffer(17597) := X"1000FFCC";
        ram_buffer(17598) := X"2EE20008";
        ram_buffer(17599) := X"8EC20000";
        ram_buffer(17600) := X"24040016";
        ram_buffer(17601) := X"8C450000";
        ram_buffer(17602) := X"AC440014";
        ram_buffer(17603) := X"00A0F809";
        ram_buffer(17604) := X"02C02021";
        ram_buffer(17605) := X"8ED00014";
        ram_buffer(17606) := X"1000FFC8";
        ram_buffer(17607) := X"00009021";
        ram_buffer(17608) := X"8C820164";
        ram_buffer(17609) := X"27BDFF68";
        ram_buffer(17610) := X"AFB00070";
        ram_buffer(17611) := X"AFA20058";
        ram_buffer(17612) := X"00408021";
        ram_buffer(17613) := X"8C820014";
        ram_buffer(17614) := X"2603000C";
        ram_buffer(17615) := X"8C480000";
        ram_buffer(17616) := X"8C470004";
        ram_buffer(17617) := X"AFB7008C";
        ram_buffer(17618) := X"AFA5009C";
        ram_buffer(17619) := X"0080B821";
        ram_buffer(17620) := X"24060018";
        ram_buffer(17621) := X"00602821";
        ram_buffer(17622) := X"27A40018";
        ram_buffer(17623) := X"AFBE0090";
        ram_buffer(17624) := X"AFB60088";
        ram_buffer(17625) := X"AFA8003C";
        ram_buffer(17626) := X"AFA70038";
        ram_buffer(17627) := X"AFBF0094";
        ram_buffer(17628) := X"AFB50084";
        ram_buffer(17629) := X"AFB40080";
        ram_buffer(17630) := X"AFB3007C";
        ram_buffer(17631) := X"AFB20078";
        ram_buffer(17632) := X"AFB10074";
        ram_buffer(17633) := X"0C027F93";
        ram_buffer(17634) := X"AFA3006C";
        ram_buffer(17635) := X"8EE200C0";
        ram_buffer(17636) := X"8E1E000C";
        ram_buffer(17637) := X"8E160010";
        ram_buffer(17638) := X"8FA70038";
        ram_buffer(17639) := X"8FA8003C";
        ram_buffer(17640) := X"10400005";
        ram_buffer(17641) := X"00000000";
        ram_buffer(17642) := X"8E020024";
        ram_buffer(17643) := X"00000000";
        ram_buffer(17644) := X"10400208";
        ram_buffer(17645) := X"26C90007";
        ram_buffer(17646) := X"8EE20108";
        ram_buffer(17647) := X"00000000";
        ram_buffer(17648) := X"18400097";
        ram_buffer(17649) := X"26E2010C";
        ram_buffer(17650) := X"AFA20054";
        ram_buffer(17651) := X"8FA2009C";
        ram_buffer(17652) := X"AFA0005C";
        ram_buffer(17653) := X"AFA20050";
        ram_buffer(17654) := X"3C02100D";
        ram_buffer(17655) := X"AFA20068";
        ram_buffer(17656) := X"3C02100D";
        ram_buffer(17657) := X"24428A64";
        ram_buffer(17658) := X"24120001";
        ram_buffer(17659) := X"AFA20064";
        ram_buffer(17660) := X"8FA20054";
        ram_buffer(17661) := X"27A60010";
        ram_buffer(17662) := X"8C430000";
        ram_buffer(17663) := X"8FA20050";
        ram_buffer(17664) := X"00000000";
        ram_buffer(17665) := X"8C420000";
        ram_buffer(17666) := X"00000000";
        ram_buffer(17667) := X"00402821";
        ram_buffer(17668) := X"AFA2004C";
        ram_buffer(17669) := X"2462003C";
        ram_buffer(17670) := X"00021080";
        ram_buffer(17671) := X"24630004";
        ram_buffer(17672) := X"02E21021";
        ram_buffer(17673) := X"8C420000";
        ram_buffer(17674) := X"00602021";
        ram_buffer(17675) := X"00042080";
        ram_buffer(17676) := X"AFA30060";
        ram_buffer(17677) := X"00C42021";
        ram_buffer(17678) := X"8C430014";
        ram_buffer(17679) := X"8C420018";
        ram_buffer(17680) := X"84B00000";
        ram_buffer(17681) := X"8C840000";
        ram_buffer(17682) := X"8FA50058";
        ram_buffer(17683) := X"2463000A";
        ram_buffer(17684) := X"2442000E";
        ram_buffer(17685) := X"02042023";
        ram_buffer(17686) := X"00031880";
        ram_buffer(17687) := X"00021080";
        ram_buffer(17688) := X"00A31821";
        ram_buffer(17689) := X"00A21021";
        ram_buffer(17690) := X"00802821";
        ram_buffer(17691) := X"AFA40038";
        ram_buffer(17692) := X"8C510004";
        ram_buffer(17693) := X"8C640004";
        ram_buffer(17694) := X"04A00188";
        ram_buffer(17695) := X"00000000";
        ram_buffer(17696) := X"10A000B2";
        ram_buffer(17697) := X"00A01021";
        ram_buffer(17698) := X"00008021";
        ram_buffer(17699) := X"00021043";
        ram_buffer(17700) := X"1440FFFE";
        ram_buffer(17701) := X"26100001";
        ram_buffer(17702) := X"00902821";
        ram_buffer(17703) := X"00101080";
        ram_buffer(17704) := X"80B30400";
        ram_buffer(17705) := X"00822021";
        ram_buffer(17706) := X"8C940000";
        ram_buffer(17707) := X"126000AF";
        ram_buffer(17708) := X"00000000";
        ram_buffer(17709) := X"02721004";
        ram_buffer(17710) := X"02D3B021";
        ram_buffer(17711) := X"2442FFFF";
        ram_buffer(17712) := X"24040018";
        ram_buffer(17713) := X"00962023";
        ram_buffer(17714) := X"00541024";
        ram_buffer(17715) := X"00821004";
        ram_buffer(17716) := X"2AC40008";
        ram_buffer(17717) := X"1480000D";
        ram_buffer(17718) := X"03C2F025";
        ram_buffer(17719) := X"241500FF";
        ram_buffer(17720) := X"001E1403";
        ram_buffer(17721) := X"24E7FFFF";
        ram_buffer(17722) := X"A1020000";
        ram_buffer(17723) := X"10E000B7";
        ram_buffer(17724) := X"305300FF";
        ram_buffer(17725) := X"127500C1";
        ram_buffer(17726) := X"25080001";
        ram_buffer(17727) := X"26D6FFF8";
        ram_buffer(17728) := X"2AC20008";
        ram_buffer(17729) := X"1040FFF6";
        ram_buffer(17730) := X"001EF200";
        ram_buffer(17731) := X"16000167";
        ram_buffer(17732) := X"02121004";
        ram_buffer(17733) := X"8FA20068";
        ram_buffer(17734) := X"00008021";
        ram_buffer(17735) := X"24428968";
        ram_buffer(17736) := X"AFA20044";
        ram_buffer(17737) := X"241400FF";
        ram_buffer(17738) := X"8C420004";
        ram_buffer(17739) := X"8FA3004C";
        ram_buffer(17740) := X"00021040";
        ram_buffer(17741) := X"00621021";
        ram_buffer(17742) := X"84420000";
        ram_buffer(17743) := X"00000000";
        ram_buffer(17744) := X"14400065";
        ram_buffer(17745) := X"AFA20048";
        ram_buffer(17746) := X"26100001";
        ram_buffer(17747) := X"8FA20044";
        ram_buffer(17748) := X"8FA30064";
        ram_buffer(17749) := X"24420004";
        ram_buffer(17750) := X"1443FFF3";
        ram_buffer(17751) := X"AFA20044";
        ram_buffer(17752) := X"1200001C";
        ram_buffer(17753) := X"00000000";
        ram_buffer(17754) := X"82300400";
        ram_buffer(17755) := X"8E310000";
        ram_buffer(17756) := X"120001FE";
        ram_buffer(17757) := X"24050027";
        ram_buffer(17758) := X"02121004";
        ram_buffer(17759) := X"02D0B021";
        ram_buffer(17760) := X"2442FFFF";
        ram_buffer(17761) := X"24030018";
        ram_buffer(17762) := X"00761823";
        ram_buffer(17763) := X"00511024";
        ram_buffer(17764) := X"00621004";
        ram_buffer(17765) := X"2AC30008";
        ram_buffer(17766) := X"1460000E";
        ram_buffer(17767) := X"03C2F025";
        ram_buffer(17768) := X"241000FF";
        ram_buffer(17769) := X"001E1403";
        ram_buffer(17770) := X"24E7FFFF";
        ram_buffer(17771) := X"A1020000";
        ram_buffer(17772) := X"10E001C6";
        ram_buffer(17773) := X"305100FF";
        ram_buffer(17774) := X"25080001";
        ram_buffer(17775) := X"123001B3";
        ram_buffer(17776) := X"00000000";
        ram_buffer(17777) := X"26D6FFF8";
        ram_buffer(17778) := X"2AC20008";
        ram_buffer(17779) := X"1040FFF5";
        ram_buffer(17780) := X"001EF200";
        ram_buffer(17781) := X"8FA50050";
        ram_buffer(17782) := X"8FA20060";
        ram_buffer(17783) := X"8CA40000";
        ram_buffer(17784) := X"00021080";
        ram_buffer(17785) := X"84840000";
        ram_buffer(17786) := X"27A90010";
        ram_buffer(17787) := X"01221021";
        ram_buffer(17788) := X"8FA6005C";
        ram_buffer(17789) := X"AC440000";
        ram_buffer(17790) := X"8FA20054";
        ram_buffer(17791) := X"8EE30108";
        ram_buffer(17792) := X"24C60001";
        ram_buffer(17793) := X"24420004";
        ram_buffer(17794) := X"AFA20054";
        ram_buffer(17795) := X"00C3182A";
        ram_buffer(17796) := X"24A20004";
        ram_buffer(17797) := X"AFA6005C";
        ram_buffer(17798) := X"1460FF75";
        ram_buffer(17799) := X"AFA20050";
        ram_buffer(17800) := X"8EE20014";
        ram_buffer(17801) := X"8FA4006C";
        ram_buffer(17802) := X"24060018";
        ram_buffer(17803) := X"AC480000";
        ram_buffer(17804) := X"AC470004";
        ram_buffer(17805) := X"27A50018";
        ram_buffer(17806) := X"AFBE0018";
        ram_buffer(17807) := X"0C027F93";
        ram_buffer(17808) := X"AFB6001C";
        ram_buffer(17809) := X"8EE400C0";
        ram_buffer(17810) := X"00000000";
        ram_buffer(17811) := X"10800071";
        ram_buffer(17812) := X"24020001";
        ram_buffer(17813) := X"8FA50058";
        ram_buffer(17814) := X"00000000";
        ram_buffer(17815) := X"8CA20024";
        ram_buffer(17816) := X"00000000";
        ram_buffer(17817) := X"14400006";
        ram_buffer(17818) := X"00000000";
        ram_buffer(17819) := X"8CA30028";
        ram_buffer(17820) := X"00801021";
        ram_buffer(17821) := X"24630001";
        ram_buffer(17822) := X"30630007";
        ram_buffer(17823) := X"ACA30028";
        ram_buffer(17824) := X"8FA30058";
        ram_buffer(17825) := X"2442FFFF";
        ram_buffer(17826) := X"AC620024";
        ram_buffer(17827) := X"10000061";
        ram_buffer(17828) := X"24020001";
        ram_buffer(17829) := X"8EF30014";
        ram_buffer(17830) := X"00000000";
        ram_buffer(17831) := X"8E62000C";
        ram_buffer(17832) := X"00000000";
        ram_buffer(17833) := X"0040F809";
        ram_buffer(17834) := X"02E02021";
        ram_buffer(17835) := X"10400059";
        ram_buffer(17836) := X"00001021";
        ram_buffer(17837) := X"8E680000";
        ram_buffer(17838) := X"8E670004";
        ram_buffer(17839) := X"12B4001E";
        ram_buffer(17840) := X"00000000";
        ram_buffer(17841) := X"26D6FFF8";
        ram_buffer(17842) := X"2AC20008";
        ram_buffer(17843) := X"10400013";
        ram_buffer(17844) := X"001EF200";
        ram_buffer(17845) := X"2610FFF0";
        ram_buffer(17846) := X"2A020010";
        ram_buffer(17847) := X"14400073";
        ram_buffer(17848) := X"00000000";
        ram_buffer(17849) := X"822304F0";
        ram_buffer(17850) := X"8E3503C0";
        ram_buffer(17851) := X"10600055";
        ram_buffer(17852) := X"00000000";
        ram_buffer(17853) := X"00721004";
        ram_buffer(17854) := X"02C3B021";
        ram_buffer(17855) := X"2442FFFF";
        ram_buffer(17856) := X"24030018";
        ram_buffer(17857) := X"00761823";
        ram_buffer(17858) := X"00551024";
        ram_buffer(17859) := X"00621004";
        ram_buffer(17860) := X"2AC30008";
        ram_buffer(17861) := X"1460FFEF";
        ram_buffer(17862) := X"03C2F025";
        ram_buffer(17863) := X"001E1403";
        ram_buffer(17864) := X"24E7FFFF";
        ram_buffer(17865) := X"A1020000";
        ram_buffer(17866) := X"10E0FFDA";
        ram_buffer(17867) := X"305500FF";
        ram_buffer(17868) := X"16B4FFE4";
        ram_buffer(17869) := X"25080001";
        ram_buffer(17870) := X"24E7FFFF";
        ram_buffer(17871) := X"10E00017";
        ram_buffer(17872) := X"A1000000";
        ram_buffer(17873) := X"1000FFDF";
        ram_buffer(17874) := X"25080001";
        ram_buffer(17875) := X"00008021";
        ram_buffer(17876) := X"00902821";
        ram_buffer(17877) := X"00101080";
        ram_buffer(17878) := X"80B30400";
        ram_buffer(17879) := X"00822021";
        ram_buffer(17880) := X"8C940000";
        ram_buffer(17881) := X"1660FF53";
        ram_buffer(17882) := X"00000000";
        ram_buffer(17883) := X"8EE20000";
        ram_buffer(17884) := X"24030027";
        ram_buffer(17885) := X"8C450000";
        ram_buffer(17886) := X"02E02021";
        ram_buffer(17887) := X"AC430014";
        ram_buffer(17888) := X"AFA80040";
        ram_buffer(17889) := X"00A0F809";
        ram_buffer(17890) := X"AFA7003C";
        ram_buffer(17891) := X"8FA80040";
        ram_buffer(17892) := X"8FA7003C";
        ram_buffer(17893) := X"1000FF48";
        ram_buffer(17894) := X"02721004";
        ram_buffer(17895) := X"8EF50014";
        ram_buffer(17896) := X"00000000";
        ram_buffer(17897) := X"8EA2000C";
        ram_buffer(17898) := X"00000000";
        ram_buffer(17899) := X"0040F809";
        ram_buffer(17900) := X"02E02021";
        ram_buffer(17901) := X"10400016";
        ram_buffer(17902) := X"26D6FFF8";
        ram_buffer(17903) := X"8EA80000";
        ram_buffer(17904) := X"8EA70004";
        ram_buffer(17905) := X"1000FFC1";
        ram_buffer(17906) := X"2AC20008";
        ram_buffer(17907) := X"8EF40014";
        ram_buffer(17908) := X"00000000";
        ram_buffer(17909) := X"8E82000C";
        ram_buffer(17910) := X"00000000";
        ram_buffer(17911) := X"0040F809";
        ram_buffer(17912) := X"02E02021";
        ram_buffer(17913) := X"1040000A";
        ram_buffer(17914) := X"00000000";
        ram_buffer(17915) := X"8E880000";
        ram_buffer(17916) := X"8E870004";
        ram_buffer(17917) := X"1675FF41";
        ram_buffer(17918) := X"00000000";
        ram_buffer(17919) := X"24E7FFFF";
        ram_buffer(17920) := X"10E0001E";
        ram_buffer(17921) := X"A1000000";
        ram_buffer(17922) := X"1000FF3C";
        ram_buffer(17923) := X"25080001";
        ram_buffer(17924) := X"00001021";
        ram_buffer(17925) := X"8FBF0094";
        ram_buffer(17926) := X"8FBE0090";
        ram_buffer(17927) := X"8FB7008C";
        ram_buffer(17928) := X"8FB60088";
        ram_buffer(17929) := X"8FB50084";
        ram_buffer(17930) := X"8FB40080";
        ram_buffer(17931) := X"8FB3007C";
        ram_buffer(17932) := X"8FB20078";
        ram_buffer(17933) := X"8FB10074";
        ram_buffer(17934) := X"8FB00070";
        ram_buffer(17935) := X"03E00008";
        ram_buffer(17936) := X"27BD0098";
        ram_buffer(17937) := X"8EE20000";
        ram_buffer(17938) := X"AFA30038";
        ram_buffer(17939) := X"8C4C0000";
        ram_buffer(17940) := X"24030027";
        ram_buffer(17941) := X"AC430014";
        ram_buffer(17942) := X"02E02021";
        ram_buffer(17943) := X"AFA80040";
        ram_buffer(17944) := X"0180F809";
        ram_buffer(17945) := X"AFA7003C";
        ram_buffer(17946) := X"8FA80040";
        ram_buffer(17947) := X"8FA7003C";
        ram_buffer(17948) := X"8FA30038";
        ram_buffer(17949) := X"1000FFA0";
        ram_buffer(17950) := X"00721004";
        ram_buffer(17951) := X"8EF30014";
        ram_buffer(17952) := X"00000000";
        ram_buffer(17953) := X"8E62000C";
        ram_buffer(17954) := X"00000000";
        ram_buffer(17955) := X"0040F809";
        ram_buffer(17956) := X"02E02021";
        ram_buffer(17957) := X"1040FFDE";
        ram_buffer(17958) := X"26D6FFF8";
        ram_buffer(17959) := X"8E680000";
        ram_buffer(17960) := X"8E670004";
        ram_buffer(17961) := X"1000FF17";
        ram_buffer(17962) := X"2AC20008";
        ram_buffer(17963) := X"8FA20048";
        ram_buffer(17964) := X"00000000";
        ram_buffer(17965) := X"044000C3";
        ram_buffer(17966) := X"00401821";
        ram_buffer(17967) := X"00021043";
        ram_buffer(17968) := X"10400004";
        ram_buffer(17969) := X"24150001";
        ram_buffer(17970) := X"00021043";
        ram_buffer(17971) := X"1440FFFE";
        ram_buffer(17972) := X"26B50001";
        ram_buffer(17973) := X"00101100";
        ram_buffer(17974) := X"00551021";
        ram_buffer(17975) := X"02222021";
        ram_buffer(17976) := X"80900400";
        ram_buffer(17977) := X"00021080";
        ram_buffer(17978) := X"02221021";
        ram_buffer(17979) := X"8C4C0000";
        ram_buffer(17980) := X"120000A6";
        ram_buffer(17981) := X"24030027";
        ram_buffer(17982) := X"02121004";
        ram_buffer(17983) := X"0216B021";
        ram_buffer(17984) := X"2442FFFF";
        ram_buffer(17985) := X"24030018";
        ram_buffer(17986) := X"00762023";
        ram_buffer(17987) := X"004C1024";
        ram_buffer(17988) := X"00821004";
        ram_buffer(17989) := X"2AC40008";
        ram_buffer(17990) := X"1480000C";
        ram_buffer(17991) := X"005EF025";
        ram_buffer(17992) := X"001E1403";
        ram_buffer(17993) := X"24E7FFFF";
        ram_buffer(17994) := X"A1020000";
        ram_buffer(17995) := X"10E0001F";
        ram_buffer(17996) := X"305000FF";
        ram_buffer(17997) := X"1214002B";
        ram_buffer(17998) := X"25080001";
        ram_buffer(17999) := X"26D6FFF8";
        ram_buffer(18000) := X"2AC20008";
        ram_buffer(18001) := X"1040FFF6";
        ram_buffer(18002) := X"001EF200";
        ram_buffer(18003) := X"02B21004";
        ram_buffer(18004) := X"8FA30048";
        ram_buffer(18005) := X"2442FFFF";
        ram_buffer(18006) := X"02B6B021";
        ram_buffer(18007) := X"0043A824";
        ram_buffer(18008) := X"24020018";
        ram_buffer(18009) := X"00561023";
        ram_buffer(18010) := X"00551004";
        ram_buffer(18011) := X"2AC30008";
        ram_buffer(18012) := X"1460000C";
        ram_buffer(18013) := X"005EF025";
        ram_buffer(18014) := X"001E1403";
        ram_buffer(18015) := X"24E7FFFF";
        ram_buffer(18016) := X"A1020000";
        ram_buffer(18017) := X"10E0001C";
        ram_buffer(18018) := X"305000FF";
        ram_buffer(18019) := X"12140026";
        ram_buffer(18020) := X"25080001";
        ram_buffer(18021) := X"26D6FFF8";
        ram_buffer(18022) := X"2AC20008";
        ram_buffer(18023) := X"1040FFF6";
        ram_buffer(18024) := X"001EF200";
        ram_buffer(18025) := X"1000FEE9";
        ram_buffer(18026) := X"00008021";
        ram_buffer(18027) := X"8EE50014";
        ram_buffer(18028) := X"02E02021";
        ram_buffer(18029) := X"8CA2000C";
        ram_buffer(18030) := X"00000000";
        ram_buffer(18031) := X"0040F809";
        ram_buffer(18032) := X"AFA50038";
        ram_buffer(18033) := X"1040FF92";
        ram_buffer(18034) := X"00000000";
        ram_buffer(18035) := X"8FA50038";
        ram_buffer(18036) := X"00000000";
        ram_buffer(18037) := X"8CA80000";
        ram_buffer(18038) := X"8CA70004";
        ram_buffer(18039) := X"1614FFD7";
        ram_buffer(18040) := X"00000000";
        ram_buffer(18041) := X"24E7FFFF";
        ram_buffer(18042) := X"10E00014";
        ram_buffer(18043) := X"A1000000";
        ram_buffer(18044) := X"1000FFD2";
        ram_buffer(18045) := X"25080001";
        ram_buffer(18046) := X"8EF50014";
        ram_buffer(18047) := X"00000000";
        ram_buffer(18048) := X"8EA2000C";
        ram_buffer(18049) := X"00000000";
        ram_buffer(18050) := X"0040F809";
        ram_buffer(18051) := X"02E02021";
        ram_buffer(18052) := X"1040FF7F";
        ram_buffer(18053) := X"00000000";
        ram_buffer(18054) := X"8EA80000";
        ram_buffer(18055) := X"8EA70004";
        ram_buffer(18056) := X"1614FFDC";
        ram_buffer(18057) := X"00000000";
        ram_buffer(18058) := X"24E7FFFF";
        ram_buffer(18059) := X"10E0000F";
        ram_buffer(18060) := X"A1000000";
        ram_buffer(18061) := X"1000FFD7";
        ram_buffer(18062) := X"25080001";
        ram_buffer(18063) := X"8EF00014";
        ram_buffer(18064) := X"00000000";
        ram_buffer(18065) := X"8E02000C";
        ram_buffer(18066) := X"00000000";
        ram_buffer(18067) := X"0040F809";
        ram_buffer(18068) := X"02E02021";
        ram_buffer(18069) := X"1040FF6E";
        ram_buffer(18070) := X"26D6FFF8";
        ram_buffer(18071) := X"8E080000";
        ram_buffer(18072) := X"8E070004";
        ram_buffer(18073) := X"1000FFB7";
        ram_buffer(18074) := X"2AC20008";
        ram_buffer(18075) := X"8EF00014";
        ram_buffer(18076) := X"00000000";
        ram_buffer(18077) := X"8E02000C";
        ram_buffer(18078) := X"00000000";
        ram_buffer(18079) := X"0040F809";
        ram_buffer(18080) := X"02E02021";
        ram_buffer(18081) := X"1040FF62";
        ram_buffer(18082) := X"26D6FFF8";
        ram_buffer(18083) := X"8E080000";
        ram_buffer(18084) := X"8E070004";
        ram_buffer(18085) := X"1000FFC1";
        ram_buffer(18086) := X"2AC20008";
        ram_buffer(18087) := X"24A3FFFF";
        ram_buffer(18088) := X"00051023";
        ram_buffer(18089) := X"1000FE78";
        ram_buffer(18090) := X"AFA30038";
        ram_buffer(18091) := X"8FA30038";
        ram_buffer(18092) := X"2442FFFF";
        ram_buffer(18093) := X"02D0B021";
        ram_buffer(18094) := X"00438024";
        ram_buffer(18095) := X"24020018";
        ram_buffer(18096) := X"00561023";
        ram_buffer(18097) := X"00501004";
        ram_buffer(18098) := X"2AC30008";
        ram_buffer(18099) := X"1460FE91";
        ram_buffer(18100) := X"03C2F025";
        ram_buffer(18101) := X"001E1403";
        ram_buffer(18102) := X"24E7FFFF";
        ram_buffer(18103) := X"241300FF";
        ram_buffer(18104) := X"A1020000";
        ram_buffer(18105) := X"10E0000C";
        ram_buffer(18106) := X"305000FF";
        ram_buffer(18107) := X"12130016";
        ram_buffer(18108) := X"25080001";
        ram_buffer(18109) := X"26D6FFF8";
        ram_buffer(18110) := X"2AC20008";
        ram_buffer(18111) := X"1440FE85";
        ram_buffer(18112) := X"001EF200";
        ram_buffer(18113) := X"001E1403";
        ram_buffer(18114) := X"24E7FFFF";
        ram_buffer(18115) := X"A1020000";
        ram_buffer(18116) := X"14E0FFF6";
        ram_buffer(18117) := X"305000FF";
        ram_buffer(18118) := X"8EF40014";
        ram_buffer(18119) := X"00000000";
        ram_buffer(18120) := X"8E82000C";
        ram_buffer(18121) := X"00000000";
        ram_buffer(18122) := X"0040F809";
        ram_buffer(18123) := X"02E02021";
        ram_buffer(18124) := X"1040FF37";
        ram_buffer(18125) := X"00000000";
        ram_buffer(18126) := X"8E880000";
        ram_buffer(18127) := X"8E870004";
        ram_buffer(18128) := X"1613FFEC";
        ram_buffer(18129) := X"00000000";
        ram_buffer(18130) := X"24E7FFFF";
        ram_buffer(18131) := X"10E00003";
        ram_buffer(18132) := X"A1000000";
        ram_buffer(18133) := X"1000FFE7";
        ram_buffer(18134) := X"25080001";
        ram_buffer(18135) := X"8EF00014";
        ram_buffer(18136) := X"00000000";
        ram_buffer(18137) := X"8E02000C";
        ram_buffer(18138) := X"00000000";
        ram_buffer(18139) := X"0040F809";
        ram_buffer(18140) := X"02E02021";
        ram_buffer(18141) := X"1040FF26";
        ram_buffer(18142) := X"26D6FFF8";
        ram_buffer(18143) := X"8E080000";
        ram_buffer(18144) := X"8E070004";
        ram_buffer(18145) := X"1000FFDD";
        ram_buffer(18146) := X"2AC20008";
        ram_buffer(18147) := X"8EE50000";
        ram_buffer(18148) := X"00000000";
        ram_buffer(18149) := X"8CA20000";
        ram_buffer(18150) := X"02E02021";
        ram_buffer(18151) := X"ACA30014";
        ram_buffer(18152) := X"AFA80040";
        ram_buffer(18153) := X"AFA7003C";
        ram_buffer(18154) := X"0040F809";
        ram_buffer(18155) := X"AFAC0038";
        ram_buffer(18156) := X"8FA80040";
        ram_buffer(18157) := X"8FA7003C";
        ram_buffer(18158) := X"8FAC0038";
        ram_buffer(18159) := X"1000FF4F";
        ram_buffer(18160) := X"02121004";
        ram_buffer(18161) := X"2463FFFF";
        ram_buffer(18162) := X"00021023";
        ram_buffer(18163) := X"1000FF3B";
        ram_buffer(18164) := X"AFA30048";
        ram_buffer(18165) := X"24130018";
        ram_buffer(18166) := X"2402007F";
        ram_buffer(18167) := X"02699823";
        ram_buffer(18168) := X"8FA30058";
        ram_buffer(18169) := X"02629804";
        ram_buffer(18170) := X"29220008";
        ram_buffer(18171) := X"8C710028";
        ram_buffer(18172) := X"1440000E";
        ram_buffer(18173) := X"027E9825";
        ram_buffer(18174) := X"01208021";
        ram_buffer(18175) := X"241200FF";
        ram_buffer(18176) := X"00131403";
        ram_buffer(18177) := X"24E7FFFF";
        ram_buffer(18178) := X"A1020000";
        ram_buffer(18179) := X"10E0003B";
        ram_buffer(18180) := X"305400FF";
        ram_buffer(18181) := X"12920045";
        ram_buffer(18182) := X"25080001";
        ram_buffer(18183) := X"2610FFF8";
        ram_buffer(18184) := X"2E020008";
        ram_buffer(18185) := X"1040FFF6";
        ram_buffer(18186) := X"00139A00";
        ram_buffer(18187) := X"2403FFFF";
        ram_buffer(18188) := X"24E7FFFF";
        ram_buffer(18189) := X"25020001";
        ram_buffer(18190) := X"10E00058";
        ram_buffer(18191) := X"A1030000";
        ram_buffer(18192) := X"2631FFD0";
        ram_buffer(18193) := X"24E7FFFF";
        ram_buffer(18194) := X"24480001";
        ram_buffer(18195) := X"10E00062";
        ram_buffer(18196) := X"A0510000";
        ram_buffer(18197) := X"8EE600EC";
        ram_buffer(18198) := X"00000000";
        ram_buffer(18199) := X"18C0005B";
        ram_buffer(18200) := X"00063080";
        ram_buffer(18201) := X"00002821";
        ram_buffer(18202) := X"27A40020";
        ram_buffer(18203) := X"AFA8003C";
        ram_buffer(18204) := X"AFA70038";
        ram_buffer(18205) := X"0C02801D";
        ram_buffer(18206) := X"0000B021";
        ram_buffer(18207) := X"8FA70038";
        ram_buffer(18208) := X"8FA8003C";
        ram_buffer(18209) := X"1000FDCC";
        ram_buffer(18210) := X"0000F021";
        ram_buffer(18211) := X"24E7FFFF";
        ram_buffer(18212) := X"A1000000";
        ram_buffer(18213) := X"14E0FE4B";
        ram_buffer(18214) := X"25080001";
        ram_buffer(18215) := X"8EF10014";
        ram_buffer(18216) := X"00000000";
        ram_buffer(18217) := X"8E22000C";
        ram_buffer(18218) := X"00000000";
        ram_buffer(18219) := X"0040F809";
        ram_buffer(18220) := X"02E02021";
        ram_buffer(18221) := X"1040FED6";
        ram_buffer(18222) := X"26D6FFF8";
        ram_buffer(18223) := X"8E280000";
        ram_buffer(18224) := X"8E270004";
        ram_buffer(18225) := X"1000FE41";
        ram_buffer(18226) := X"2AC20008";
        ram_buffer(18227) := X"8EF30014";
        ram_buffer(18228) := X"00000000";
        ram_buffer(18229) := X"8E62000C";
        ram_buffer(18230) := X"00000000";
        ram_buffer(18231) := X"0040F809";
        ram_buffer(18232) := X"02E02021";
        ram_buffer(18233) := X"1040FECA";
        ram_buffer(18234) := X"00000000";
        ram_buffer(18235) := X"8E680000";
        ram_buffer(18236) := X"8E670004";
        ram_buffer(18237) := X"1000FE31";
        ram_buffer(18238) := X"00000000";
        ram_buffer(18239) := X"8EF50014";
        ram_buffer(18240) := X"00000000";
        ram_buffer(18241) := X"8EA2000C";
        ram_buffer(18242) := X"00000000";
        ram_buffer(18243) := X"0040F809";
        ram_buffer(18244) := X"02E02021";
        ram_buffer(18245) := X"1040FEBE";
        ram_buffer(18246) := X"00000000";
        ram_buffer(18247) := X"8EA80000";
        ram_buffer(18248) := X"8EA70004";
        ram_buffer(18249) := X"1692FFBD";
        ram_buffer(18250) := X"00000000";
        ram_buffer(18251) := X"24E7FFFF";
        ram_buffer(18252) := X"A1000000";
        ram_buffer(18253) := X"14E0FFB9";
        ram_buffer(18254) := X"25080001";
        ram_buffer(18255) := X"8EF40014";
        ram_buffer(18256) := X"00000000";
        ram_buffer(18257) := X"8E82000C";
        ram_buffer(18258) := X"00000000";
        ram_buffer(18259) := X"0040F809";
        ram_buffer(18260) := X"02E02021";
        ram_buffer(18261) := X"1040FEAE";
        ram_buffer(18262) := X"2610FFF8";
        ram_buffer(18263) := X"8E880000";
        ram_buffer(18264) := X"8E870004";
        ram_buffer(18265) := X"1000FFAF";
        ram_buffer(18266) := X"2E020008";
        ram_buffer(18267) := X"8EE30000";
        ram_buffer(18268) := X"00000000";
        ram_buffer(18269) := X"8C620000";
        ram_buffer(18270) := X"02E02021";
        ram_buffer(18271) := X"AC650014";
        ram_buffer(18272) := X"AFA8003C";
        ram_buffer(18273) := X"0040F809";
        ram_buffer(18274) := X"AFA70038";
        ram_buffer(18275) := X"8FA8003C";
        ram_buffer(18276) := X"8FA70038";
        ram_buffer(18277) := X"1000FDF9";
        ram_buffer(18278) := X"02121004";
        ram_buffer(18279) := X"8EF00014";
        ram_buffer(18280) := X"00000000";
        ram_buffer(18281) := X"8E02000C";
        ram_buffer(18282) := X"00000000";
        ram_buffer(18283) := X"0040F809";
        ram_buffer(18284) := X"02E02021";
        ram_buffer(18285) := X"1040FE96";
        ram_buffer(18286) := X"2631FFD0";
        ram_buffer(18287) := X"8E020000";
        ram_buffer(18288) := X"8E070004";
        ram_buffer(18289) := X"1000FFA0";
        ram_buffer(18290) := X"24E7FFFF";
        ram_buffer(18291) := X"0000B021";
        ram_buffer(18292) := X"1000FD79";
        ram_buffer(18293) := X"0000F021";
        ram_buffer(18294) := X"8EF00014";
        ram_buffer(18295) := X"00000000";
        ram_buffer(18296) := X"8E02000C";
        ram_buffer(18297) := X"00000000";
        ram_buffer(18298) := X"0040F809";
        ram_buffer(18299) := X"02E02021";
        ram_buffer(18300) := X"1040FE88";
        ram_buffer(18301) := X"00001021";
        ram_buffer(18302) := X"8E080000";
        ram_buffer(18303) := X"8E070004";
        ram_buffer(18304) := X"1000FF94";
        ram_buffer(18305) := X"00000000";
        ram_buffer(18306) := X"27BDFAC8";
        ram_buffer(18307) := X"AFB1051C";
        ram_buffer(18308) := X"8CD10000";
        ram_buffer(18309) := X"AFB00518";
        ram_buffer(18310) := X"AFBF0534";
        ram_buffer(18311) := X"AFB60530";
        ram_buffer(18312) := X"AFB5052C";
        ram_buffer(18313) := X"AFB40528";
        ram_buffer(18314) := X"AFB30524";
        ram_buffer(18315) := X"AFB20520";
        ram_buffer(18316) := X"1220004E";
        ram_buffer(18317) := X"00A08021";
        ram_buffer(18318) := X"26150001";
        ram_buffer(18319) := X"24120001";
        ram_buffer(18320) := X"0000A021";
        ram_buffer(18321) := X"24160011";
        ram_buffer(18322) := X"92B30000";
        ram_buffer(18323) := X"27A20414";
        ram_buffer(18324) := X"00542021";
        ram_buffer(18325) := X"02603021";
        ram_buffer(18326) := X"12600003";
        ram_buffer(18327) := X"02402821";
        ram_buffer(18328) := X"0C02801D";
        ram_buffer(18329) := X"0293A021";
        ram_buffer(18330) := X"26520001";
        ram_buffer(18331) := X"1656FFF6";
        ram_buffer(18332) := X"26B50001";
        ram_buffer(18333) := X"27A20010";
        ram_buffer(18334) := X"00541021";
        ram_buffer(18335) := X"A0400404";
        ram_buffer(18336) := X"83A50414";
        ram_buffer(18337) := X"00000000";
        ram_buffer(18338) := X"10A00014";
        ram_buffer(18339) := X"00A03821";
        ram_buffer(18340) := X"00002021";
        ram_buffer(18341) := X"00003021";
        ram_buffer(18342) := X"27A80414";
        ram_buffer(18343) := X"14A70030";
        ram_buffer(18344) := X"00061880";
        ram_buffer(18345) := X"24C20001";
        ram_buffer(18346) := X"27A50010";
        ram_buffer(18347) := X"00A31821";
        ram_buffer(18348) := X"01021021";
        ram_buffer(18349) := X"80450000";
        ram_buffer(18350) := X"AC640000";
        ram_buffer(18351) := X"00483023";
        ram_buffer(18352) := X"24840001";
        ram_buffer(18353) := X"24630004";
        ram_buffer(18354) := X"10A7FFFA";
        ram_buffer(18355) := X"24420001";
        ram_buffer(18356) := X"00042040";
        ram_buffer(18357) := X"14A0FFF1";
        ram_buffer(18358) := X"24E70001";
        ram_buffer(18359) := X"24060100";
        ram_buffer(18360) := X"00002821";
        ram_buffer(18361) := X"0C02801D";
        ram_buffer(18362) := X"26240400";
        ram_buffer(18363) := X"12800012";
        ram_buffer(18364) := X"26940011";
        ram_buffer(18365) := X"26030011";
        ram_buffer(18366) := X"27A40010";
        ram_buffer(18367) := X"27A50414";
        ram_buffer(18368) := X"02148021";
        ram_buffer(18369) := X"90620000";
        ram_buffer(18370) := X"8C860000";
        ram_buffer(18371) := X"00021080";
        ram_buffer(18372) := X"02221021";
        ram_buffer(18373) := X"AC460000";
        ram_buffer(18374) := X"90620000";
        ram_buffer(18375) := X"90A60000";
        ram_buffer(18376) := X"02221021";
        ram_buffer(18377) := X"24630001";
        ram_buffer(18378) := X"A0460400";
        ram_buffer(18379) := X"24840004";
        ram_buffer(18380) := X"1470FFF4";
        ram_buffer(18381) := X"24A50001";
        ram_buffer(18382) := X"8FBF0534";
        ram_buffer(18383) := X"8FB60530";
        ram_buffer(18384) := X"8FB5052C";
        ram_buffer(18385) := X"8FB40528";
        ram_buffer(18386) := X"8FB30524";
        ram_buffer(18387) := X"8FB20520";
        ram_buffer(18388) := X"8FB1051C";
        ram_buffer(18389) := X"8FB00518";
        ram_buffer(18390) := X"03E00008";
        ram_buffer(18391) := X"27BD0538";
        ram_buffer(18392) := X"00042040";
        ram_buffer(18393) := X"1000FFCD";
        ram_buffer(18394) := X"24E70001";
        ram_buffer(18395) := X"8C820004";
        ram_buffer(18396) := X"00C09021";
        ram_buffer(18397) := X"8C420000";
        ram_buffer(18398) := X"24060500";
        ram_buffer(18399) := X"0040F809";
        ram_buffer(18400) := X"24050001";
        ram_buffer(18401) := X"AE420000";
        ram_buffer(18402) := X"1000FFAB";
        ram_buffer(18403) := X"00408821";
        ram_buffer(18404) := X"27BDFFC8";
        ram_buffer(18405) := X"AFBE0030";
        ram_buffer(18406) := X"AFB60028";
        ram_buffer(18407) := X"AFB20018";
        ram_buffer(18408) := X"AFBF0034";
        ram_buffer(18409) := X"AFB7002C";
        ram_buffer(18410) := X"AFB50024";
        ram_buffer(18411) := X"AFB40020";
        ram_buffer(18412) := X"AFB3001C";
        ram_buffer(18413) := X"AFB10014";
        ram_buffer(18414) := X"AFB00010";
        ram_buffer(18415) := X"0080F021";
        ram_buffer(18416) := X"8C920164";
        ram_buffer(18417) := X"14A0007F";
        ram_buffer(18418) := X"00A0B021";
        ram_buffer(18419) := X"3C031009";
        ram_buffer(18420) := X"3C021009";
        ram_buffer(18421) := X"2463117C";
        ram_buffer(18422) := X"24421320";
        ram_buffer(18423) := X"8FC400EC";
        ram_buffer(18424) := X"AE430008";
        ram_buffer(18425) := X"18800037";
        ram_buffer(18426) := X"AE420004";
        ram_buffer(18427) := X"27D500F0";
        ram_buffer(18428) := X"26540014";
        ram_buffer(18429) := X"00009821";
        ram_buffer(18430) := X"24170031";
        ram_buffer(18431) := X"8EA20000";
        ram_buffer(18432) := X"00000000";
        ram_buffer(18433) := X"8C510014";
        ram_buffer(18434) := X"8C500018";
        ram_buffer(18435) := X"2E220004";
        ram_buffer(18436) := X"10400061";
        ram_buffer(18437) := X"00000000";
        ram_buffer(18438) := X"26220014";
        ram_buffer(18439) := X"00021080";
        ram_buffer(18440) := X"03C21021";
        ram_buffer(18441) := X"8C420000";
        ram_buffer(18442) := X"00000000";
        ram_buffer(18443) := X"10400058";
        ram_buffer(18444) := X"00000000";
        ram_buffer(18445) := X"2E020004";
        ram_buffer(18446) := X"10400035";
        ram_buffer(18447) := X"26020018";
        ram_buffer(18448) := X"00021080";
        ram_buffer(18449) := X"03C21021";
        ram_buffer(18450) := X"8C420000";
        ram_buffer(18451) := X"00000000";
        ram_buffer(18452) := X"1040002D";
        ram_buffer(18453) := X"00000000";
        ram_buffer(18454) := X"12C00038";
        ram_buffer(18455) := X"26220014";
        ram_buffer(18456) := X"00118880";
        ram_buffer(18457) := X"02518821";
        ram_buffer(18458) := X"8E24004C";
        ram_buffer(18459) := X"00000000";
        ram_buffer(18460) := X"10800062";
        ram_buffer(18461) := X"24060404";
        ram_buffer(18462) := X"00108080";
        ram_buffer(18463) := X"24060404";
        ram_buffer(18464) := X"00002821";
        ram_buffer(18465) := X"0C02801D";
        ram_buffer(18466) := X"02508021";
        ram_buffer(18467) := X"8E04005C";
        ram_buffer(18468) := X"00000000";
        ram_buffer(18469) := X"10800050";
        ram_buffer(18470) := X"24060404";
        ram_buffer(18471) := X"24060404";
        ram_buffer(18472) := X"0C02801D";
        ram_buffer(18473) := X"00002821";
        ram_buffer(18474) := X"AE800000";
        ram_buffer(18475) := X"8FC200EC";
        ram_buffer(18476) := X"26730001";
        ram_buffer(18477) := X"0262102A";
        ram_buffer(18478) := X"26B50004";
        ram_buffer(18479) := X"1440FFCF";
        ram_buffer(18480) := X"26940004";
        ram_buffer(18481) := X"8FC200C0";
        ram_buffer(18482) := X"8FBF0034";
        ram_buffer(18483) := X"AE40000C";
        ram_buffer(18484) := X"AE400010";
        ram_buffer(18485) := X"AE420024";
        ram_buffer(18486) := X"AE400028";
        ram_buffer(18487) := X"8FBE0030";
        ram_buffer(18488) := X"8FB7002C";
        ram_buffer(18489) := X"8FB60028";
        ram_buffer(18490) := X"8FB50024";
        ram_buffer(18491) := X"8FB40020";
        ram_buffer(18492) := X"8FB3001C";
        ram_buffer(18493) := X"8FB20018";
        ram_buffer(18494) := X"8FB10014";
        ram_buffer(18495) := X"8FB00010";
        ram_buffer(18496) := X"03E00008";
        ram_buffer(18497) := X"27BD0038";
        ram_buffer(18498) := X"16C0FFD5";
        ram_buffer(18499) := X"00000000";
        ram_buffer(18500) := X"8FC20000";
        ram_buffer(18501) := X"00000000";
        ram_buffer(18502) := X"AC500018";
        ram_buffer(18503) := X"8FC30000";
        ram_buffer(18504) := X"AC570014";
        ram_buffer(18505) := X"8C620000";
        ram_buffer(18506) := X"00000000";
        ram_buffer(18507) := X"0040F809";
        ram_buffer(18508) := X"03C02021";
        ram_buffer(18509) := X"16C0FFCA";
        ram_buffer(18510) := X"26220014";
        ram_buffer(18511) := X"2626000A";
        ram_buffer(18512) := X"00021080";
        ram_buffer(18513) := X"03C21021";
        ram_buffer(18514) := X"00063080";
        ram_buffer(18515) := X"8C450000";
        ram_buffer(18516) := X"02463021";
        ram_buffer(18517) := X"03C02021";
        ram_buffer(18518) := X"0C024782";
        ram_buffer(18519) := X"24C60004";
        ram_buffer(18520) := X"26020018";
        ram_buffer(18521) := X"2606000E";
        ram_buffer(18522) := X"00021080";
        ram_buffer(18523) := X"03C21021";
        ram_buffer(18524) := X"00063080";
        ram_buffer(18525) := X"02463021";
        ram_buffer(18526) := X"8C450000";
        ram_buffer(18527) := X"24C60004";
        ram_buffer(18528) := X"0C024782";
        ram_buffer(18529) := X"03C02021";
        ram_buffer(18530) := X"1000FFC8";
        ram_buffer(18531) := X"AE800000";
        ram_buffer(18532) := X"16C0FFA8";
        ram_buffer(18533) := X"00000000";
        ram_buffer(18534) := X"8FC20000";
        ram_buffer(18535) := X"00000000";
        ram_buffer(18536) := X"AC510018";
        ram_buffer(18537) := X"8FC30000";
        ram_buffer(18538) := X"AC570014";
        ram_buffer(18539) := X"8C620000";
        ram_buffer(18540) := X"00000000";
        ram_buffer(18541) := X"0040F809";
        ram_buffer(18542) := X"03C02021";
        ram_buffer(18543) := X"1000FF9E";
        ram_buffer(18544) := X"2E020004";
        ram_buffer(18545) := X"3C031009";
        ram_buffer(18546) := X"3C021009";
        ram_buffer(18547) := X"24632714";
        ram_buffer(18548) := X"1000FF82";
        ram_buffer(18549) := X"24420F70";
        ram_buffer(18550) := X"8FC20004";
        ram_buffer(18551) := X"03C02021";
        ram_buffer(18552) := X"8C420000";
        ram_buffer(18553) := X"00000000";
        ram_buffer(18554) := X"0040F809";
        ram_buffer(18555) := X"24050001";
        ram_buffer(18556) := X"AE02005C";
        ram_buffer(18557) := X"1000FFA9";
        ram_buffer(18558) := X"00402021";
        ram_buffer(18559) := X"8FC20004";
        ram_buffer(18560) := X"03C02021";
        ram_buffer(18561) := X"8C420000";
        ram_buffer(18562) := X"00000000";
        ram_buffer(18563) := X"0040F809";
        ram_buffer(18564) := X"24050001";
        ram_buffer(18565) := X"AE22004C";
        ram_buffer(18566) := X"1000FF97";
        ram_buffer(18567) := X"00402021";
        ram_buffer(18568) := X"27BDF7A0";
        ram_buffer(18569) := X"AFB30850";
        ram_buffer(18570) := X"AFB2084C";
        ram_buffer(18571) := X"AFB10848";
        ram_buffer(18572) := X"AFB00844";
        ram_buffer(18573) := X"27B10818";
        ram_buffer(18574) := X"00C09021";
        ram_buffer(18575) := X"00809821";
        ram_buffer(18576) := X"24060404";
        ram_buffer(18577) := X"27A40414";
        ram_buffer(18578) := X"00A08021";
        ram_buffer(18579) := X"00002821";
        ram_buffer(18580) := X"AFBF085C";
        ram_buffer(18581) := X"AFB50858";
        ram_buffer(18582) := X"AFB40854";
        ram_buffer(18583) := X"AFA00818";
        ram_buffer(18584) := X"AE200004";
        ram_buffer(18585) := X"AE200008";
        ram_buffer(18586) := X"AE20000C";
        ram_buffer(18587) := X"AE200010";
        ram_buffer(18588) := X"AE200014";
        ram_buffer(18589) := X"AE200018";
        ram_buffer(18590) := X"AE20001C";
        ram_buffer(18591) := X"0C02801D";
        ram_buffer(18592) := X"A2200020";
        ram_buffer(18593) := X"24060404";
        ram_buffer(18594) := X"240500FF";
        ram_buffer(18595) := X"0C02801D";
        ram_buffer(18596) := X"27A40010";
        ram_buffer(18597) := X"24020001";
        ram_buffer(18598) := X"3C0A3B9A";
        ram_buffer(18599) := X"AE420400";
        ram_buffer(18600) := X"354ACA00";
        ram_buffer(18601) := X"24060101";
        ram_buffer(18602) := X"02402021";
        ram_buffer(18603) := X"02402821";
        ram_buffer(18604) := X"01404021";
        ram_buffer(18605) := X"00001021";
        ram_buffer(18606) := X"2409FFFF";
        ram_buffer(18607) := X"8CA30000";
        ram_buffer(18608) := X"24A50004";
        ram_buffer(18609) := X"10600005";
        ram_buffer(18610) := X"0103382A";
        ram_buffer(18611) := X"14E00003";
        ram_buffer(18612) := X"00000000";
        ram_buffer(18613) := X"00404821";
        ram_buffer(18614) := X"00604021";
        ram_buffer(18615) := X"24420001";
        ram_buffer(18616) := X"1446FFF6";
        ram_buffer(18617) := X"00000000";
        ram_buffer(18618) := X"01403821";
        ram_buffer(18619) := X"00001021";
        ram_buffer(18620) := X"2408FFFF";
        ram_buffer(18621) := X"8C830000";
        ram_buffer(18622) := X"24840004";
        ram_buffer(18623) := X"10600007";
        ram_buffer(18624) := X"00E3282A";
        ram_buffer(18625) := X"14A00005";
        ram_buffer(18626) := X"00000000";
        ram_buffer(18627) := X"11220003";
        ram_buffer(18628) := X"00000000";
        ram_buffer(18629) := X"00404021";
        ram_buffer(18630) := X"00603821";
        ram_buffer(18631) := X"24420001";
        ram_buffer(18632) := X"1446FFF4";
        ram_buffer(18633) := X"00000000";
        ram_buffer(18634) := X"0500002E";
        ram_buffer(18635) := X"00094880";
        ram_buffer(18636) := X"00083880";
        ram_buffer(18637) := X"27A20010";
        ram_buffer(18638) := X"00491021";
        ram_buffer(18639) := X"02496021";
        ram_buffer(18640) := X"02475821";
        ram_buffer(18641) := X"8D850000";
        ram_buffer(18642) := X"8D6D0000";
        ram_buffer(18643) := X"8C440404";
        ram_buffer(18644) := X"8C430000";
        ram_buffer(18645) := X"00AD2821";
        ram_buffer(18646) := X"24840001";
        ram_buffer(18647) := X"AD850000";
        ram_buffer(18648) := X"AC440404";
        ram_buffer(18649) := X"0460001D";
        ram_buffer(18650) := X"AD600000";
        ram_buffer(18651) := X"00031080";
        ram_buffer(18652) := X"27A30010";
        ram_buffer(18653) := X"00622021";
        ram_buffer(18654) := X"8C850404";
        ram_buffer(18655) := X"8C830000";
        ram_buffer(18656) := X"24A50001";
        ram_buffer(18657) := X"0461FFF9";
        ram_buffer(18658) := X"AC850404";
        ram_buffer(18659) := X"27A40010";
        ram_buffer(18660) := X"27A30010";
        ram_buffer(18661) := X"00671821";
        ram_buffer(18662) := X"00821021";
        ram_buffer(18663) := X"AC480000";
        ram_buffer(18664) := X"8C640404";
        ram_buffer(18665) := X"8C620000";
        ram_buffer(18666) := X"24840001";
        ram_buffer(18667) := X"0440FFBE";
        ram_buffer(18668) := X"AC640404";
        ram_buffer(18669) := X"00021080";
        ram_buffer(18670) := X"27A30010";
        ram_buffer(18671) := X"00621821";
        ram_buffer(18672) := X"8C640404";
        ram_buffer(18673) := X"8C620000";
        ram_buffer(18674) := X"24840001";
        ram_buffer(18675) := X"0441FFF9";
        ram_buffer(18676) := X"AC640404";
        ram_buffer(18677) := X"1000FFB5";
        ram_buffer(18678) := X"02402021";
        ram_buffer(18679) := X"1000FFEB";
        ram_buffer(18680) := X"01201021";
        ram_buffer(18681) := X"27B40414";
        ram_buffer(18682) := X"24150026";
        ram_buffer(18683) := X"8E920000";
        ram_buffer(18684) := X"26940004";
        ram_buffer(18685) := X"12400009";
        ram_buffer(18686) := X"2A420021";
        ram_buffer(18687) := X"1040009D";
        ram_buffer(18688) := X"02602021";
        ram_buffer(18689) := X"27A20010";
        ram_buffer(18690) := X"00529021";
        ram_buffer(18691) := X"92420808";
        ram_buffer(18692) := X"00000000";
        ram_buffer(18693) := X"24420001";
        ram_buffer(18694) := X"A2420808";
        ram_buffer(18695) := X"1634FFF3";
        ram_buffer(18696) := X"24080001";
        ram_buffer(18697) := X"27A50835";
        ram_buffer(18698) := X"27A90825";
        ram_buffer(18699) := X"01114023";
        ram_buffer(18700) := X"90A60003";
        ram_buffer(18701) := X"00000000";
        ram_buffer(18702) := X"10C00021";
        ram_buffer(18703) := X"00000000";
        ram_buffer(18704) := X"01053821";
        ram_buffer(18705) := X"90A20001";
        ram_buffer(18706) := X"00000000";
        ram_buffer(18707) := X"14400091";
        ram_buffer(18708) := X"00A01021";
        ram_buffer(18709) := X"00E01821";
        ram_buffer(18710) := X"2442FFFF";
        ram_buffer(18711) := X"90440001";
        ram_buffer(18712) := X"00000000";
        ram_buffer(18713) := X"1080FFFC";
        ram_buffer(18714) := X"2463FFFF";
        ram_buffer(18715) := X"90A40002";
        ram_buffer(18716) := X"24C6FFFE";
        ram_buffer(18717) := X"24840001";
        ram_buffer(18718) := X"A0A40002";
        ram_buffer(18719) := X"24620001";
        ram_buffer(18720) := X"27A40010";
        ram_buffer(18721) := X"A0A60003";
        ram_buffer(18722) := X"00821021";
        ram_buffer(18723) := X"90440808";
        ram_buffer(18724) := X"27A60010";
        ram_buffer(18725) := X"24840002";
        ram_buffer(18726) := X"00C31821";
        ram_buffer(18727) := X"A0440808";
        ram_buffer(18728) := X"90620808";
        ram_buffer(18729) := X"00000000";
        ram_buffer(18730) := X"2442FFFF";
        ram_buffer(18731) := X"A0620808";
        ram_buffer(18732) := X"90A60003";
        ram_buffer(18733) := X"00000000";
        ram_buffer(18734) := X"14C0FFE2";
        ram_buffer(18735) := X"00000000";
        ram_buffer(18736) := X"24A5FFFF";
        ram_buffer(18737) := X"14A9FFDA";
        ram_buffer(18738) := X"00000000";
        ram_buffer(18739) := X"93A30828";
        ram_buffer(18740) := X"00000000";
        ram_buffer(18741) := X"1460003F";
        ram_buffer(18742) := X"24020010";
        ram_buffer(18743) := X"93A30827";
        ram_buffer(18744) := X"00000000";
        ram_buffer(18745) := X"1460006D";
        ram_buffer(18746) := X"00000000";
        ram_buffer(18747) := X"93A30826";
        ram_buffer(18748) := X"00000000";
        ram_buffer(18749) := X"14600085";
        ram_buffer(18750) := X"00000000";
        ram_buffer(18751) := X"93A30825";
        ram_buffer(18752) := X"00000000";
        ram_buffer(18753) := X"1460007F";
        ram_buffer(18754) := X"00000000";
        ram_buffer(18755) := X"93A30824";
        ram_buffer(18756) := X"00000000";
        ram_buffer(18757) := X"14600079";
        ram_buffer(18758) := X"00000000";
        ram_buffer(18759) := X"93A30823";
        ram_buffer(18760) := X"00000000";
        ram_buffer(18761) := X"14600073";
        ram_buffer(18762) := X"00000000";
        ram_buffer(18763) := X"93A30822";
        ram_buffer(18764) := X"00000000";
        ram_buffer(18765) := X"1460006D";
        ram_buffer(18766) := X"00000000";
        ram_buffer(18767) := X"93A30821";
        ram_buffer(18768) := X"00000000";
        ram_buffer(18769) := X"14600067";
        ram_buffer(18770) := X"00000000";
        ram_buffer(18771) := X"93A30820";
        ram_buffer(18772) := X"00000000";
        ram_buffer(18773) := X"14600061";
        ram_buffer(18774) := X"00000000";
        ram_buffer(18775) := X"93A3081F";
        ram_buffer(18776) := X"00000000";
        ram_buffer(18777) := X"1460005B";
        ram_buffer(18778) := X"00000000";
        ram_buffer(18779) := X"93A3081E";
        ram_buffer(18780) := X"00000000";
        ram_buffer(18781) := X"14600055";
        ram_buffer(18782) := X"00000000";
        ram_buffer(18783) := X"93A3081D";
        ram_buffer(18784) := X"00000000";
        ram_buffer(18785) := X"1460004F";
        ram_buffer(18786) := X"00000000";
        ram_buffer(18787) := X"93A3081C";
        ram_buffer(18788) := X"00000000";
        ram_buffer(18789) := X"14600049";
        ram_buffer(18790) := X"00000000";
        ram_buffer(18791) := X"93A3081B";
        ram_buffer(18792) := X"00000000";
        ram_buffer(18793) := X"14600043";
        ram_buffer(18794) := X"00000000";
        ram_buffer(18795) := X"93A3081A";
        ram_buffer(18796) := X"00000000";
        ram_buffer(18797) := X"1460003D";
        ram_buffer(18798) := X"00000000";
        ram_buffer(18799) := X"93A30819";
        ram_buffer(18800) := X"00000000";
        ram_buffer(18801) := X"14600037";
        ram_buffer(18802) := X"00000000";
        ram_buffer(18803) := X"93A30818";
        ram_buffer(18804) := X"00001021";
        ram_buffer(18805) := X"27A40010";
        ram_buffer(18806) := X"00821021";
        ram_buffer(18807) := X"2463FFFF";
        ram_buffer(18808) := X"24060011";
        ram_buffer(18809) := X"02202821";
        ram_buffer(18810) := X"02002021";
        ram_buffer(18811) := X"0C027F93";
        ram_buffer(18812) := X"A0430808";
        ram_buffer(18813) := X"24050001";
        ram_buffer(18814) := X"00003821";
        ram_buffer(18815) := X"24060100";
        ram_buffer(18816) := X"24080021";
        ram_buffer(18817) := X"27A30414";
        ram_buffer(18818) := X"10000004";
        ram_buffer(18819) := X"00001021";
        ram_buffer(18820) := X"24420001";
        ram_buffer(18821) := X"1046000A";
        ram_buffer(18822) := X"00000000";
        ram_buffer(18823) := X"8C640000";
        ram_buffer(18824) := X"00000000";
        ram_buffer(18825) := X"1485FFFA";
        ram_buffer(18826) := X"24630004";
        ram_buffer(18827) := X"02072021";
        ram_buffer(18828) := X"A0820011";
        ram_buffer(18829) := X"24420001";
        ram_buffer(18830) := X"1446FFF8";
        ram_buffer(18831) := X"24E70001";
        ram_buffer(18832) := X"24A50001";
        ram_buffer(18833) := X"14A8FFEF";
        ram_buffer(18834) := X"00000000";
        ram_buffer(18835) := X"8FBF085C";
        ram_buffer(18836) := X"AE000114";
        ram_buffer(18837) := X"8FB50858";
        ram_buffer(18838) := X"8FB40854";
        ram_buffer(18839) := X"8FB30850";
        ram_buffer(18840) := X"8FB2084C";
        ram_buffer(18841) := X"8FB10848";
        ram_buffer(18842) := X"8FB00844";
        ram_buffer(18843) := X"03E00008";
        ram_buffer(18844) := X"27BD0860";
        ram_buffer(18845) := X"8E620000";
        ram_buffer(18846) := X"00000000";
        ram_buffer(18847) := X"8C430000";
        ram_buffer(18848) := X"00000000";
        ram_buffer(18849) := X"0060F809";
        ram_buffer(18850) := X"AC550014";
        ram_buffer(18851) := X"1000FF5E";
        ram_buffer(18852) := X"27A20010";
        ram_buffer(18853) := X"1000FF75";
        ram_buffer(18854) := X"00E01821";
        ram_buffer(18855) := X"1000FFCD";
        ram_buffer(18856) := X"2402000F";
        ram_buffer(18857) := X"1000FFCB";
        ram_buffer(18858) := X"24020001";
        ram_buffer(18859) := X"1000FFC9";
        ram_buffer(18860) := X"24020002";
        ram_buffer(18861) := X"1000FFC7";
        ram_buffer(18862) := X"24020003";
        ram_buffer(18863) := X"1000FFC5";
        ram_buffer(18864) := X"24020004";
        ram_buffer(18865) := X"1000FFC3";
        ram_buffer(18866) := X"24020005";
        ram_buffer(18867) := X"1000FFC1";
        ram_buffer(18868) := X"24020006";
        ram_buffer(18869) := X"1000FFBF";
        ram_buffer(18870) := X"24020007";
        ram_buffer(18871) := X"1000FFBD";
        ram_buffer(18872) := X"24020008";
        ram_buffer(18873) := X"1000FFBB";
        ram_buffer(18874) := X"24020009";
        ram_buffer(18875) := X"1000FFB9";
        ram_buffer(18876) := X"2402000A";
        ram_buffer(18877) := X"1000FFB7";
        ram_buffer(18878) := X"2402000B";
        ram_buffer(18879) := X"1000FFB5";
        ram_buffer(18880) := X"2402000C";
        ram_buffer(18881) := X"1000FFB3";
        ram_buffer(18882) := X"2402000D";
        ram_buffer(18883) := X"1000FFB1";
        ram_buffer(18884) := X"2402000E";
        ram_buffer(18885) := X"8C8200EC";
        ram_buffer(18886) := X"27BDFFA0";
        ram_buffer(18887) := X"AFB20040";
        ram_buffer(18888) := X"AFBF005C";
        ram_buffer(18889) := X"AFBE0058";
        ram_buffer(18890) := X"AFB70054";
        ram_buffer(18891) := X"AFB60050";
        ram_buffer(18892) := X"AFB5004C";
        ram_buffer(18893) := X"AFB40048";
        ram_buffer(18894) := X"AFB30044";
        ram_buffer(18895) := X"AFB1003C";
        ram_buffer(18896) := X"AFB00038";
        ram_buffer(18897) := X"8C920164";
        ram_buffer(18898) := X"AFA00020";
        ram_buffer(18899) := X"AFA00024";
        ram_buffer(18900) := X"AFA00028";
        ram_buffer(18901) := X"AFA0002C";
        ram_buffer(18902) := X"AFA00010";
        ram_buffer(18903) := X"AFA00014";
        ram_buffer(18904) := X"AFA00018";
        ram_buffer(18905) := X"18400039";
        ram_buffer(18906) := X"AFA0001C";
        ram_buffer(18907) := X"0080A021";
        ram_buffer(18908) := X"249E00F0";
        ram_buffer(18909) := X"0000B821";
        ram_buffer(18910) := X"24130001";
        ram_buffer(18911) := X"8FC20000";
        ram_buffer(18912) := X"26F70001";
        ram_buffer(18913) := X"8C510014";
        ram_buffer(18914) := X"8C500018";
        ram_buffer(18915) := X"0011B080";
        ram_buffer(18916) := X"27A20010";
        ram_buffer(18917) := X"00561021";
        ram_buffer(18918) := X"8C420010";
        ram_buffer(18919) := X"0010A880";
        ram_buffer(18920) := X"02963021";
        ram_buffer(18921) := X"02951821";
        ram_buffer(18922) := X"14400010";
        ram_buffer(18923) := X"27DE0004";
        ram_buffer(18924) := X"8CC50050";
        ram_buffer(18925) := X"00000000";
        ram_buffer(18926) := X"10A00030";
        ram_buffer(18927) := X"02802021";
        ram_buffer(18928) := X"26310012";
        ram_buffer(18929) := X"00118880";
        ram_buffer(18930) := X"02518821";
        ram_buffer(18931) := X"8E260004";
        ram_buffer(18932) := X"02802021";
        ram_buffer(18933) := X"0C024888";
        ram_buffer(18934) := X"AFA30030";
        ram_buffer(18935) := X"27A20010";
        ram_buffer(18936) := X"0056B021";
        ram_buffer(18937) := X"8FA30030";
        ram_buffer(18938) := X"AED30010";
        ram_buffer(18939) := X"27A20010";
        ram_buffer(18940) := X"00551021";
        ram_buffer(18941) := X"8C420000";
        ram_buffer(18942) := X"00000000";
        ram_buffer(18943) := X"1440000E";
        ram_buffer(18944) := X"00000000";
        ram_buffer(18945) := X"8C650060";
        ram_buffer(18946) := X"00000000";
        ram_buffer(18947) := X"10A00024";
        ram_buffer(18948) := X"02802021";
        ram_buffer(18949) := X"26100016";
        ram_buffer(18950) := X"00108080";
        ram_buffer(18951) := X"02508021";
        ram_buffer(18952) := X"8E060004";
        ram_buffer(18953) := X"0C024888";
        ram_buffer(18954) := X"02802021";
        ram_buffer(18955) := X"27A20010";
        ram_buffer(18956) := X"0055A821";
        ram_buffer(18957) := X"AEB30000";
        ram_buffer(18958) := X"8E8200EC";
        ram_buffer(18959) := X"00000000";
        ram_buffer(18960) := X"02E2102A";
        ram_buffer(18961) := X"1440FFCD";
        ram_buffer(18962) := X"00000000";
        ram_buffer(18963) := X"8FBF005C";
        ram_buffer(18964) := X"8FBE0058";
        ram_buffer(18965) := X"8FB70054";
        ram_buffer(18966) := X"8FB60050";
        ram_buffer(18967) := X"8FB5004C";
        ram_buffer(18968) := X"8FB40048";
        ram_buffer(18969) := X"8FB30044";
        ram_buffer(18970) := X"8FB20040";
        ram_buffer(18971) := X"8FB1003C";
        ram_buffer(18972) := X"8FB00038";
        ram_buffer(18973) := X"03E00008";
        ram_buffer(18974) := X"27BD0060";
        ram_buffer(18975) := X"AFA30034";
        ram_buffer(18976) := X"0C0264A0";
        ram_buffer(18977) := X"AFA60030";
        ram_buffer(18978) := X"8FA60030";
        ram_buffer(18979) := X"00000000";
        ram_buffer(18980) := X"ACC20050";
        ram_buffer(18981) := X"8FA30034";
        ram_buffer(18982) := X"1000FFC9";
        ram_buffer(18983) := X"00402821";
        ram_buffer(18984) := X"0C0264A0";
        ram_buffer(18985) := X"AFA30030";
        ram_buffer(18986) := X"8FA30030";
        ram_buffer(18987) := X"00402821";
        ram_buffer(18988) := X"1000FFD8";
        ram_buffer(18989) := X"AC620060";
        ram_buffer(18990) := X"8C820004";
        ram_buffer(18991) := X"27BDFFE0";
        ram_buffer(18992) := X"8C420000";
        ram_buffer(18993) := X"2406006C";
        ram_buffer(18994) := X"AFBF001C";
        ram_buffer(18995) := X"AFB10018";
        ram_buffer(18996) := X"AFB00014";
        ram_buffer(18997) := X"24050001";
        ram_buffer(18998) := X"0040F809";
        ram_buffer(18999) := X"00808821";
        ram_buffer(19000) := X"00408021";
        ram_buffer(19001) := X"AE220164";
        ram_buffer(19002) := X"3C021009";
        ram_buffer(19003) := X"24421F90";
        ram_buffer(19004) := X"2604003C";
        ram_buffer(19005) := X"24060010";
        ram_buffer(19006) := X"AE020000";
        ram_buffer(19007) := X"0C02801D";
        ram_buffer(19008) := X"00002821";
        ram_buffer(19009) := X"2604002C";
        ram_buffer(19010) := X"24060010";
        ram_buffer(19011) := X"0C02801D";
        ram_buffer(19012) := X"00002821";
        ram_buffer(19013) := X"2604005C";
        ram_buffer(19014) := X"24060010";
        ram_buffer(19015) := X"0C02801D";
        ram_buffer(19016) := X"00002821";
        ram_buffer(19017) := X"8FBF001C";
        ram_buffer(19018) := X"8FB10018";
        ram_buffer(19019) := X"2604004C";
        ram_buffer(19020) := X"8FB00014";
        ram_buffer(19021) := X"24060010";
        ram_buffer(19022) := X"00002821";
        ram_buffer(19023) := X"0802801D";
        ram_buffer(19024) := X"27BD0020";
        ram_buffer(19025) := X"27BDFFC8";
        ram_buffer(19026) := X"8C82013C";
        ram_buffer(19027) := X"AFB50024";
        ram_buffer(19028) := X"8C950164";
        ram_buffer(19029) := X"AFB40020";
        ram_buffer(19030) := X"AFB20018";
        ram_buffer(19031) := X"AFB10014";
        ram_buffer(19032) := X"AFBF0034";
        ram_buffer(19033) := X"AFBE0030";
        ram_buffer(19034) := X"AFB7002C";
        ram_buffer(19035) := X"AFB60028";
        ram_buffer(19036) := X"AFB3001C";
        ram_buffer(19037) := X"AFB00010";
        ram_buffer(19038) := X"0080A021";
        ram_buffer(19039) := X"AEA40020";
        ram_buffer(19040) := X"AEA5000C";
        ram_buffer(19041) := X"8C920134";
        ram_buffer(19042) := X"14400048";
        ram_buffer(19043) := X"00A08821";
        ram_buffer(19044) := X"1640005B";
        ram_buffer(19045) := X"3C021009";
        ram_buffer(19046) := X"3C021009";
        ram_buffer(19047) := X"244247B8";
        ram_buffer(19048) := X"AEA20004";
        ram_buffer(19049) := X"16200048";
        ram_buffer(19050) := X"3C021009";
        ram_buffer(19051) := X"3C021009";
        ram_buffer(19052) := X"24422E08";
        ram_buffer(19053) := X"8E8300EC";
        ram_buffer(19054) := X"00000000";
        ram_buffer(19055) := X"18600028";
        ram_buffer(19056) := X"AEA20008";
        ram_buffer(19057) := X"269E00F0";
        ram_buffer(19058) := X"26B70024";
        ram_buffer(19059) := X"0000B021";
        ram_buffer(19060) := X"24130031";
        ram_buffer(19061) := X"8FC20000";
        ram_buffer(19062) := X"1640004C";
        ram_buffer(19063) := X"AEE00000";
        ram_buffer(19064) := X"8E83013C";
        ram_buffer(19065) := X"00000000";
        ram_buffer(19066) := X"14600017";
        ram_buffer(19067) := X"00000000";
        ram_buffer(19068) := X"8C500014";
        ram_buffer(19069) := X"00000000";
        ram_buffer(19070) := X"2E020004";
        ram_buffer(19071) := X"1040006D";
        ram_buffer(19072) := X"26020014";
        ram_buffer(19073) := X"00021080";
        ram_buffer(19074) := X"02821021";
        ram_buffer(19075) := X"8C420000";
        ram_buffer(19076) := X"00000000";
        ram_buffer(19077) := X"10400065";
        ram_buffer(19078) := X"00000000";
        ram_buffer(19079) := X"16200049";
        ram_buffer(19080) := X"26020014";
        ram_buffer(19081) := X"26060012";
        ram_buffer(19082) := X"00021080";
        ram_buffer(19083) := X"00063080";
        ram_buffer(19084) := X"02821021";
        ram_buffer(19085) := X"02A63021";
        ram_buffer(19086) := X"8C450000";
        ram_buffer(19087) := X"24C60004";
        ram_buffer(19088) := X"0C024782";
        ram_buffer(19089) := X"02802021";
        ram_buffer(19090) := X"8E8200EC";
        ram_buffer(19091) := X"26D60001";
        ram_buffer(19092) := X"02C2102A";
        ram_buffer(19093) := X"27DE0004";
        ram_buffer(19094) := X"1440FFDE";
        ram_buffer(19095) := X"26F70004";
        ram_buffer(19096) := X"8E8200C0";
        ram_buffer(19097) := X"8FBF0034";
        ram_buffer(19098) := X"AEA00038";
        ram_buffer(19099) := X"AEA0003C";
        ram_buffer(19100) := X"AEA00018";
        ram_buffer(19101) := X"AEA0001C";
        ram_buffer(19102) := X"AEA20044";
        ram_buffer(19103) := X"AEA00048";
        ram_buffer(19104) := X"8FBE0030";
        ram_buffer(19105) := X"8FB7002C";
        ram_buffer(19106) := X"8FB60028";
        ram_buffer(19107) := X"8FB50024";
        ram_buffer(19108) := X"8FB40020";
        ram_buffer(19109) := X"8FB3001C";
        ram_buffer(19110) := X"8FB20018";
        ram_buffer(19111) := X"8FB10014";
        ram_buffer(19112) := X"8FB00010";
        ram_buffer(19113) := X"03E00008";
        ram_buffer(19114) := X"27BD0038";
        ram_buffer(19115) := X"16400008";
        ram_buffer(19116) := X"3C021009";
        ram_buffer(19117) := X"3C021009";
        ram_buffer(19118) := X"24424D30";
        ram_buffer(19119) := X"1220FFBB";
        ram_buffer(19120) := X"AEA20004";
        ram_buffer(19121) := X"3C021009";
        ram_buffer(19122) := X"1000FFBA";
        ram_buffer(19123) := X"244237F0";
        ram_buffer(19124) := X"8EA30040";
        ram_buffer(19125) := X"24424FF0";
        ram_buffer(19126) := X"1460FFB2";
        ram_buffer(19127) := X"AEA20004";
        ram_buffer(19128) := X"8C820004";
        ram_buffer(19129) := X"240603E8";
        ram_buffer(19130) := X"8C420000";
        ram_buffer(19131) := X"00000000";
        ram_buffer(19132) := X"0040F809";
        ram_buffer(19133) := X"24050001";
        ram_buffer(19134) := X"1000FFAA";
        ram_buffer(19135) := X"AEA20040";
        ram_buffer(19136) := X"24426428";
        ram_buffer(19137) := X"1000FFA7";
        ram_buffer(19138) := X"AEA20004";
        ram_buffer(19139) := X"8C500018";
        ram_buffer(19140) := X"00000000";
        ram_buffer(19141) := X"2E020004";
        ram_buffer(19142) := X"10400017";
        ram_buffer(19143) := X"AEB00034";
        ram_buffer(19144) := X"26020018";
        ram_buffer(19145) := X"00021080";
        ram_buffer(19146) := X"02821021";
        ram_buffer(19147) := X"8C420000";
        ram_buffer(19148) := X"00000000";
        ram_buffer(19149) := X"1040000E";
        ram_buffer(19150) := X"00000000";
        ram_buffer(19151) := X"1220FFB9";
        ram_buffer(19152) := X"26020018";
        ram_buffer(19153) := X"00108080";
        ram_buffer(19154) := X"02B08021";
        ram_buffer(19155) := X"8E04005C";
        ram_buffer(19156) := X"00000000";
        ram_buffer(19157) := X"10800022";
        ram_buffer(19158) := X"24060404";
        ram_buffer(19159) := X"24060404";
        ram_buffer(19160) := X"0C02801D";
        ram_buffer(19161) := X"00002821";
        ram_buffer(19162) := X"1000FFB7";
        ram_buffer(19163) := X"00000000";
        ram_buffer(19164) := X"1620FFF4";
        ram_buffer(19165) := X"00000000";
        ram_buffer(19166) := X"8E820000";
        ram_buffer(19167) := X"00000000";
        ram_buffer(19168) := X"AC500018";
        ram_buffer(19169) := X"8E830000";
        ram_buffer(19170) := X"AC530014";
        ram_buffer(19171) := X"8C620000";
        ram_buffer(19172) := X"00000000";
        ram_buffer(19173) := X"0040F809";
        ram_buffer(19174) := X"02802021";
        ram_buffer(19175) := X"1620FFE9";
        ram_buffer(19176) := X"26020018";
        ram_buffer(19177) := X"1000FFA0";
        ram_buffer(19178) := X"26060012";
        ram_buffer(19179) := X"1620FFE5";
        ram_buffer(19180) := X"00000000";
        ram_buffer(19181) := X"8E820000";
        ram_buffer(19182) := X"00000000";
        ram_buffer(19183) := X"AC500018";
        ram_buffer(19184) := X"8E830000";
        ram_buffer(19185) := X"AC530014";
        ram_buffer(19186) := X"8C620000";
        ram_buffer(19187) := X"00000000";
        ram_buffer(19188) := X"0040F809";
        ram_buffer(19189) := X"02802021";
        ram_buffer(19190) := X"1000FF90";
        ram_buffer(19191) := X"00000000";
        ram_buffer(19192) := X"8E820004";
        ram_buffer(19193) := X"02802021";
        ram_buffer(19194) := X"8C420000";
        ram_buffer(19195) := X"00000000";
        ram_buffer(19196) := X"0040F809";
        ram_buffer(19197) := X"24050001";
        ram_buffer(19198) := X"AE02005C";
        ram_buffer(19199) := X"1000FFD7";
        ram_buffer(19200) := X"00402021";
        ram_buffer(19201) := X"8C82000C";
        ram_buffer(19202) := X"27BDFFC8";
        ram_buffer(19203) := X"AFB00010";
        ram_buffer(19204) := X"AFBF0034";
        ram_buffer(19205) := X"AFBE0030";
        ram_buffer(19206) := X"AFB7002C";
        ram_buffer(19207) := X"AFB60028";
        ram_buffer(19208) := X"AFB50024";
        ram_buffer(19209) := X"AFB40020";
        ram_buffer(19210) := X"AFB3001C";
        ram_buffer(19211) := X"AFB20018";
        ram_buffer(19212) := X"AFB10014";
        ram_buffer(19213) := X"00808021";
        ram_buffer(19214) := X"1040000E";
        ram_buffer(19215) := X"AC800038";
        ram_buffer(19216) := X"8FBF0034";
        ram_buffer(19217) := X"AE00003C";
        ram_buffer(19218) := X"8FBE0030";
        ram_buffer(19219) := X"8FB7002C";
        ram_buffer(19220) := X"8FB60028";
        ram_buffer(19221) := X"8FB50024";
        ram_buffer(19222) := X"8FB40020";
        ram_buffer(19223) := X"8FB3001C";
        ram_buffer(19224) := X"8FB20018";
        ram_buffer(19225) := X"8FB10014";
        ram_buffer(19226) := X"8FB00010";
        ram_buffer(19227) := X"03E00008";
        ram_buffer(19228) := X"27BD0038";
        ram_buffer(19229) := X"8C83003C";
        ram_buffer(19230) := X"00000000";
        ram_buffer(19231) := X"1060FFF0";
        ram_buffer(19232) := X"241200FF";
        ram_buffer(19233) := X"8C950040";
        ram_buffer(19234) := X"8C94001C";
        ram_buffer(19235) := X"26B30001";
        ram_buffer(19236) := X"02A3A821";
        ram_buffer(19237) := X"1440001F";
        ram_buffer(19238) := X"26970001";
        ram_buffer(19239) := X"9262FFFF";
        ram_buffer(19240) := X"24030018";
        ram_buffer(19241) := X"0077F023";
        ram_buffer(19242) := X"30420001";
        ram_buffer(19243) := X"8E040018";
        ram_buffer(19244) := X"03C21004";
        ram_buffer(19245) := X"2AE30008";
        ram_buffer(19246) := X"14600013";
        ram_buffer(19247) := X"0044F025";
        ram_buffer(19248) := X"8E030010";
        ram_buffer(19249) := X"001E1403";
        ram_buffer(19250) := X"24640001";
        ram_buffer(19251) := X"AE040010";
        ram_buffer(19252) := X"A0620000";
        ram_buffer(19253) := X"8E030014";
        ram_buffer(19254) := X"26F7FFF8";
        ram_buffer(19255) := X"2463FFFF";
        ram_buffer(19256) := X"AE030014";
        ram_buffer(19257) := X"10600010";
        ram_buffer(19258) := X"305100FF";
        ram_buffer(19259) := X"12320025";
        ram_buffer(19260) := X"00000000";
        ram_buffer(19261) := X"2AE20008";
        ram_buffer(19262) := X"1040FFF1";
        ram_buffer(19263) := X"001EF200";
        ram_buffer(19264) := X"2694FFF9";
        ram_buffer(19265) := X"32970007";
        ram_buffer(19266) := X"AE1E0018";
        ram_buffer(19267) := X"AE17001C";
        ram_buffer(19268) := X"02E0A021";
        ram_buffer(19269) := X"12B3FFCA";
        ram_buffer(19270) := X"26730001";
        ram_buffer(19271) := X"8E02000C";
        ram_buffer(19272) := X"1000FFDC";
        ram_buffer(19273) := X"00000000";
        ram_buffer(19274) := X"8E040020";
        ram_buffer(19275) := X"00000000";
        ram_buffer(19276) := X"8C960014";
        ram_buffer(19277) := X"00000000";
        ram_buffer(19278) := X"8EC2000C";
        ram_buffer(19279) := X"00000000";
        ram_buffer(19280) := X"0040F809";
        ram_buffer(19281) := X"00000000";
        ram_buffer(19282) := X"14400009";
        ram_buffer(19283) := X"24030016";
        ram_buffer(19284) := X"8E040020";
        ram_buffer(19285) := X"00000000";
        ram_buffer(19286) := X"8C820000";
        ram_buffer(19287) := X"00000000";
        ram_buffer(19288) := X"8C460000";
        ram_buffer(19289) := X"00000000";
        ram_buffer(19290) := X"00C0F809";
        ram_buffer(19291) := X"AC430014";
        ram_buffer(19292) := X"8EC40000";
        ram_buffer(19293) := X"8EC20004";
        ram_buffer(19294) := X"AE040010";
        ram_buffer(19295) := X"1632FFDD";
        ram_buffer(19296) := X"AE020014";
        ram_buffer(19297) := X"8E020010";
        ram_buffer(19298) := X"00000000";
        ram_buffer(19299) := X"24430001";
        ram_buffer(19300) := X"AE030010";
        ram_buffer(19301) := X"A0400000";
        ram_buffer(19302) := X"8E020014";
        ram_buffer(19303) := X"00000000";
        ram_buffer(19304) := X"2442FFFF";
        ram_buffer(19305) := X"1440FFD3";
        ram_buffer(19306) := X"AE020014";
        ram_buffer(19307) := X"8E040020";
        ram_buffer(19308) := X"00000000";
        ram_buffer(19309) := X"8C910014";
        ram_buffer(19310) := X"00000000";
        ram_buffer(19311) := X"8E22000C";
        ram_buffer(19312) := X"00000000";
        ram_buffer(19313) := X"0040F809";
        ram_buffer(19314) := X"00000000";
        ram_buffer(19315) := X"14400009";
        ram_buffer(19316) := X"24050016";
        ram_buffer(19317) := X"8E040020";
        ram_buffer(19318) := X"00000000";
        ram_buffer(19319) := X"8C820000";
        ram_buffer(19320) := X"00000000";
        ram_buffer(19321) := X"8C430000";
        ram_buffer(19322) := X"00000000";
        ram_buffer(19323) := X"0060F809";
        ram_buffer(19324) := X"AC450014";
        ram_buffer(19325) := X"8E230000";
        ram_buffer(19326) := X"8E220004";
        ram_buffer(19327) := X"AE030010";
        ram_buffer(19328) := X"1000FFBC";
        ram_buffer(19329) := X"AE020014";
        ram_buffer(19330) := X"27BDFFC8";
        ram_buffer(19331) := X"8C820014";
        ram_buffer(19332) := X"AFB00010";
        ram_buffer(19333) := X"8C900164";
        ram_buffer(19334) := X"AFB20018";
        ram_buffer(19335) := X"8C430004";
        ram_buffer(19336) := X"00809021";
        ram_buffer(19337) := X"8C440000";
        ram_buffer(19338) := X"8E020038";
        ram_buffer(19339) := X"AFBF0034";
        ram_buffer(19340) := X"AFBE0030";
        ram_buffer(19341) := X"AFB7002C";
        ram_buffer(19342) := X"AFB60028";
        ram_buffer(19343) := X"AFB50024";
        ram_buffer(19344) := X"AFB40020";
        ram_buffer(19345) := X"AFB3001C";
        ram_buffer(19346) := X"AFB10014";
        ram_buffer(19347) := X"AE040010";
        ram_buffer(19348) := X"1040001A";
        ram_buffer(19349) := X"AE030014";
        ram_buffer(19350) := X"00021043";
        ram_buffer(19351) := X"10400159";
        ram_buffer(19352) := X"00000000";
        ram_buffer(19353) := X"0000B821";
        ram_buffer(19354) := X"00021043";
        ram_buffer(19355) := X"1440FFFE";
        ram_buffer(19356) := X"26F70001";
        ram_buffer(19357) := X"00171900";
        ram_buffer(19358) := X"8E04000C";
        ram_buffer(19359) := X"8E020034";
        ram_buffer(19360) := X"10800070";
        ram_buffer(19361) := X"00032080";
        ram_buffer(19362) := X"24420016";
        ram_buffer(19363) := X"00021080";
        ram_buffer(19364) := X"02021021";
        ram_buffer(19365) := X"8C420004";
        ram_buffer(19366) := X"00031880";
        ram_buffer(19367) := X"00431821";
        ram_buffer(19368) := X"8C620000";
        ram_buffer(19369) := X"00000000";
        ram_buffer(19370) := X"24420001";
        ram_buffer(19371) := X"AC620000";
        ram_buffer(19372) := X"0C024B01";
        ram_buffer(19373) := X"02002021";
        ram_buffer(19374) := X"8E040010";
        ram_buffer(19375) := X"8E02000C";
        ram_buffer(19376) := X"00000000";
        ram_buffer(19377) := X"144000B1";
        ram_buffer(19378) := X"24140018";
        ram_buffer(19379) := X"8E17001C";
        ram_buffer(19380) := X"00000000";
        ram_buffer(19381) := X"26F70007";
        ram_buffer(19382) := X"0297A023";
        ram_buffer(19383) := X"8E050018";
        ram_buffer(19384) := X"2402007F";
        ram_buffer(19385) := X"02821004";
        ram_buffer(19386) := X"2AE30008";
        ram_buffer(19387) := X"146000A7";
        ram_buffer(19388) := X"0045A025";
        ram_buffer(19389) := X"24130016";
        ram_buffer(19390) := X"241600FF";
        ram_buffer(19391) := X"00141C03";
        ram_buffer(19392) := X"24820001";
        ram_buffer(19393) := X"AE020010";
        ram_buffer(19394) := X"A0830000";
        ram_buffer(19395) := X"8E020014";
        ram_buffer(19396) := X"307100FF";
        ram_buffer(19397) := X"2442FFFF";
        ram_buffer(19398) := X"10400019";
        ram_buffer(19399) := X"AE020014";
        ram_buffer(19400) := X"8E040010";
        ram_buffer(19401) := X"1236002D";
        ram_buffer(19402) := X"00000000";
        ram_buffer(19403) := X"26F7FFF8";
        ram_buffer(19404) := X"2AE30008";
        ram_buffer(19405) := X"1060FFF1";
        ram_buffer(19406) := X"0014A200";
        ram_buffer(19407) := X"8E430014";
        ram_buffer(19408) := X"8FBF0034";
        ram_buffer(19409) := X"AE000018";
        ram_buffer(19410) := X"AE00001C";
        ram_buffer(19411) := X"8FBE0030";
        ram_buffer(19412) := X"8FB7002C";
        ram_buffer(19413) := X"8FB60028";
        ram_buffer(19414) := X"8FB50024";
        ram_buffer(19415) := X"8FB40020";
        ram_buffer(19416) := X"8FB3001C";
        ram_buffer(19417) := X"8FB20018";
        ram_buffer(19418) := X"8FB10014";
        ram_buffer(19419) := X"8FB00010";
        ram_buffer(19420) := X"AC640000";
        ram_buffer(19421) := X"AC620004";
        ram_buffer(19422) := X"03E00008";
        ram_buffer(19423) := X"27BD0038";
        ram_buffer(19424) := X"8E040020";
        ram_buffer(19425) := X"00000000";
        ram_buffer(19426) := X"8C950014";
        ram_buffer(19427) := X"00000000";
        ram_buffer(19428) := X"8EA2000C";
        ram_buffer(19429) := X"00000000";
        ram_buffer(19430) := X"0040F809";
        ram_buffer(19431) := X"00000000";
        ram_buffer(19432) := X"14400009";
        ram_buffer(19433) := X"00000000";
        ram_buffer(19434) := X"8E040020";
        ram_buffer(19435) := X"00000000";
        ram_buffer(19436) := X"8C820000";
        ram_buffer(19437) := X"00000000";
        ram_buffer(19438) := X"8C430000";
        ram_buffer(19439) := X"00000000";
        ram_buffer(19440) := X"0060F809";
        ram_buffer(19441) := X"AC530014";
        ram_buffer(19442) := X"8EA40000";
        ram_buffer(19443) := X"8EA20004";
        ram_buffer(19444) := X"AE040010";
        ram_buffer(19445) := X"1636FFD5";
        ram_buffer(19446) := X"AE020014";
        ram_buffer(19447) := X"24820001";
        ram_buffer(19448) := X"AE020010";
        ram_buffer(19449) := X"A0800000";
        ram_buffer(19450) := X"8E020014";
        ram_buffer(19451) := X"00000000";
        ram_buffer(19452) := X"2442FFFF";
        ram_buffer(19453) := X"10400004";
        ram_buffer(19454) := X"AE020014";
        ram_buffer(19455) := X"8E040010";
        ram_buffer(19456) := X"1000FFCB";
        ram_buffer(19457) := X"26F7FFF8";
        ram_buffer(19458) := X"8E040020";
        ram_buffer(19459) := X"00000000";
        ram_buffer(19460) := X"8C910014";
        ram_buffer(19461) := X"00000000";
        ram_buffer(19462) := X"8E22000C";
        ram_buffer(19463) := X"00000000";
        ram_buffer(19464) := X"0040F809";
        ram_buffer(19465) := X"00000000";
        ram_buffer(19466) := X"1040005B";
        ram_buffer(19467) := X"00000000";
        ram_buffer(19468) := X"8E240000";
        ram_buffer(19469) := X"8E220004";
        ram_buffer(19470) := X"AE040010";
        ram_buffer(19471) := X"1000FFBB";
        ram_buffer(19472) := X"AE020014";
        ram_buffer(19473) := X"24420012";
        ram_buffer(19474) := X"00021080";
        ram_buffer(19475) := X"02021021";
        ram_buffer(19476) := X"8C420004";
        ram_buffer(19477) := X"00000000";
        ram_buffer(19478) := X"00431821";
        ram_buffer(19479) := X"80710400";
        ram_buffer(19480) := X"00441021";
        ram_buffer(19481) := X"8C550000";
        ram_buffer(19482) := X"8E13001C";
        ram_buffer(19483) := X"122000C7";
        ram_buffer(19484) := X"24020001";
        ram_buffer(19485) := X"02221004";
        ram_buffer(19486) := X"2442FFFF";
        ram_buffer(19487) := X"00551824";
        ram_buffer(19488) := X"02338821";
        ram_buffer(19489) := X"24020018";
        ram_buffer(19490) := X"00511023";
        ram_buffer(19491) := X"8E150018";
        ram_buffer(19492) := X"00431004";
        ram_buffer(19493) := X"2A230008";
        ram_buffer(19494) := X"0055A825";
        ram_buffer(19495) := X"0220B021";
        ram_buffer(19496) := X"14600012";
        ram_buffer(19497) := X"241400FF";
        ram_buffer(19498) := X"8E030010";
        ram_buffer(19499) := X"00151403";
        ram_buffer(19500) := X"24640001";
        ram_buffer(19501) := X"AE040010";
        ram_buffer(19502) := X"A0620000";
        ram_buffer(19503) := X"8E030014";
        ram_buffer(19504) := X"26D6FFF8";
        ram_buffer(19505) := X"2463FFFF";
        ram_buffer(19506) := X"AE030014";
        ram_buffer(19507) := X"1060003F";
        ram_buffer(19508) := X"305300FF";
        ram_buffer(19509) := X"12740054";
        ram_buffer(19510) := X"00000000";
        ram_buffer(19511) := X"2AC20008";
        ram_buffer(19512) := X"1040FFF1";
        ram_buffer(19513) := X"0015AA00";
        ram_buffer(19514) := X"32310007";
        ram_buffer(19515) := X"AE150018";
        ram_buffer(19516) := X"12E0FF6F";
        ram_buffer(19517) := X"AE11001C";
        ram_buffer(19518) := X"8E03000C";
        ram_buffer(19519) := X"8E040038";
        ram_buffer(19520) := X"1460FF6B";
        ram_buffer(19521) := X"24020001";
        ram_buffer(19522) := X"02E21004";
        ram_buffer(19523) := X"02378821";
        ram_buffer(19524) := X"2442FFFF";
        ram_buffer(19525) := X"24030018";
        ram_buffer(19526) := X"00711823";
        ram_buffer(19527) := X"00441024";
        ram_buffer(19528) := X"00621004";
        ram_buffer(19529) := X"2A230008";
        ram_buffer(19530) := X"14600015";
        ram_buffer(19531) := X"0055A825";
        ram_buffer(19532) := X"0220B821";
        ram_buffer(19533) := X"24140016";
        ram_buffer(19534) := X"241E00FF";
        ram_buffer(19535) := X"8E030010";
        ram_buffer(19536) := X"00151403";
        ram_buffer(19537) := X"24640001";
        ram_buffer(19538) := X"AE040010";
        ram_buffer(19539) := X"A0620000";
        ram_buffer(19540) := X"8E030014";
        ram_buffer(19541) := X"26F7FFF8";
        ram_buffer(19542) := X"2463FFFF";
        ram_buffer(19543) := X"AE030014";
        ram_buffer(19544) := X"10600052";
        ram_buffer(19545) := X"305300FF";
        ram_buffer(19546) := X"127E0067";
        ram_buffer(19547) := X"00000000";
        ram_buffer(19548) := X"2AE20008";
        ram_buffer(19549) := X"1040FFF1";
        ram_buffer(19550) := X"0015AA00";
        ram_buffer(19551) := X"32310007";
        ram_buffer(19552) := X"AE150018";
        ram_buffer(19553) := X"1000FF4A";
        ram_buffer(19554) := X"AE11001C";
        ram_buffer(19555) := X"8E020014";
        ram_buffer(19556) := X"1000FF6A";
        ram_buffer(19557) := X"00000000";
        ram_buffer(19558) := X"8E040020";
        ram_buffer(19559) := X"00000000";
        ram_buffer(19560) := X"8C820000";
        ram_buffer(19561) := X"00000000";
        ram_buffer(19562) := X"8C430000";
        ram_buffer(19563) := X"00000000";
        ram_buffer(19564) := X"0060F809";
        ram_buffer(19565) := X"AC530014";
        ram_buffer(19566) := X"8E240000";
        ram_buffer(19567) := X"8E220004";
        ram_buffer(19568) := X"AE040010";
        ram_buffer(19569) := X"1000FF59";
        ram_buffer(19570) := X"AE020014";
        ram_buffer(19571) := X"8E040020";
        ram_buffer(19572) := X"00000000";
        ram_buffer(19573) := X"8C9E0014";
        ram_buffer(19574) := X"00000000";
        ram_buffer(19575) := X"8FC2000C";
        ram_buffer(19576) := X"00000000";
        ram_buffer(19577) := X"0040F809";
        ram_buffer(19578) := X"00000000";
        ram_buffer(19579) := X"14400009";
        ram_buffer(19580) := X"24050016";
        ram_buffer(19581) := X"8E040020";
        ram_buffer(19582) := X"00000000";
        ram_buffer(19583) := X"8C820000";
        ram_buffer(19584) := X"00000000";
        ram_buffer(19585) := X"8C430000";
        ram_buffer(19586) := X"00000000";
        ram_buffer(19587) := X"0060F809";
        ram_buffer(19588) := X"AC450014";
        ram_buffer(19589) := X"8FC30000";
        ram_buffer(19590) := X"8FC20004";
        ram_buffer(19591) := X"AE030010";
        ram_buffer(19592) := X"1674FFAE";
        ram_buffer(19593) := X"AE020014";
        ram_buffer(19594) := X"8E020010";
        ram_buffer(19595) := X"00000000";
        ram_buffer(19596) := X"24430001";
        ram_buffer(19597) := X"AE030010";
        ram_buffer(19598) := X"A0400000";
        ram_buffer(19599) := X"8E020014";
        ram_buffer(19600) := X"00000000";
        ram_buffer(19601) := X"2442FFFF";
        ram_buffer(19602) := X"1440FFA4";
        ram_buffer(19603) := X"AE020014";
        ram_buffer(19604) := X"8E040020";
        ram_buffer(19605) := X"00000000";
        ram_buffer(19606) := X"8C930014";
        ram_buffer(19607) := X"00000000";
        ram_buffer(19608) := X"8E62000C";
        ram_buffer(19609) := X"00000000";
        ram_buffer(19610) := X"0040F809";
        ram_buffer(19611) := X"00000000";
        ram_buffer(19612) := X"14400009";
        ram_buffer(19613) := X"24050016";
        ram_buffer(19614) := X"8E040020";
        ram_buffer(19615) := X"00000000";
        ram_buffer(19616) := X"8C820000";
        ram_buffer(19617) := X"00000000";
        ram_buffer(19618) := X"8C430000";
        ram_buffer(19619) := X"00000000";
        ram_buffer(19620) := X"0060F809";
        ram_buffer(19621) := X"AC450014";
        ram_buffer(19622) := X"8E630000";
        ram_buffer(19623) := X"8E620004";
        ram_buffer(19624) := X"AE030010";
        ram_buffer(19625) := X"1000FF8D";
        ram_buffer(19626) := X"AE020014";
        ram_buffer(19627) := X"8E040020";
        ram_buffer(19628) := X"00000000";
        ram_buffer(19629) := X"8C960014";
        ram_buffer(19630) := X"00000000";
        ram_buffer(19631) := X"8EC2000C";
        ram_buffer(19632) := X"00000000";
        ram_buffer(19633) := X"0040F809";
        ram_buffer(19634) := X"00000000";
        ram_buffer(19635) := X"14400009";
        ram_buffer(19636) := X"00000000";
        ram_buffer(19637) := X"8E040020";
        ram_buffer(19638) := X"00000000";
        ram_buffer(19639) := X"8C820000";
        ram_buffer(19640) := X"00000000";
        ram_buffer(19641) := X"8C430000";
        ram_buffer(19642) := X"00000000";
        ram_buffer(19643) := X"0060F809";
        ram_buffer(19644) := X"AC540014";
        ram_buffer(19645) := X"8EC30000";
        ram_buffer(19646) := X"8EC20004";
        ram_buffer(19647) := X"AE030010";
        ram_buffer(19648) := X"167EFF9B";
        ram_buffer(19649) := X"AE020014";
        ram_buffer(19650) := X"8E020010";
        ram_buffer(19651) := X"00000000";
        ram_buffer(19652) := X"24430001";
        ram_buffer(19653) := X"AE030010";
        ram_buffer(19654) := X"A0400000";
        ram_buffer(19655) := X"8E020014";
        ram_buffer(19656) := X"00000000";
        ram_buffer(19657) := X"2442FFFF";
        ram_buffer(19658) := X"1440FF91";
        ram_buffer(19659) := X"AE020014";
        ram_buffer(19660) := X"8E040020";
        ram_buffer(19661) := X"00000000";
        ram_buffer(19662) := X"8C930014";
        ram_buffer(19663) := X"00000000";
        ram_buffer(19664) := X"8E62000C";
        ram_buffer(19665) := X"00000000";
        ram_buffer(19666) := X"0040F809";
        ram_buffer(19667) := X"00000000";
        ram_buffer(19668) := X"14400009";
        ram_buffer(19669) := X"00000000";
        ram_buffer(19670) := X"8E040020";
        ram_buffer(19671) := X"00000000";
        ram_buffer(19672) := X"8C820000";
        ram_buffer(19673) := X"00000000";
        ram_buffer(19674) := X"8C430000";
        ram_buffer(19675) := X"00000000";
        ram_buffer(19676) := X"0060F809";
        ram_buffer(19677) := X"AC540014";
        ram_buffer(19678) := X"8E630000";
        ram_buffer(19679) := X"8E620004";
        ram_buffer(19680) := X"AE030010";
        ram_buffer(19681) := X"1000FF7A";
        ram_buffer(19682) := X"AE020014";
        ram_buffer(19683) := X"8E040020";
        ram_buffer(19684) := X"24050027";
        ram_buffer(19685) := X"8C820000";
        ram_buffer(19686) := X"00000000";
        ram_buffer(19687) := X"8C430000";
        ram_buffer(19688) := X"00000000";
        ram_buffer(19689) := X"0060F809";
        ram_buffer(19690) := X"AC450014";
        ram_buffer(19691) := X"8E02000C";
        ram_buffer(19692) := X"00000000";
        ram_buffer(19693) := X"1440FEBE";
        ram_buffer(19694) := X"24020001";
        ram_buffer(19695) := X"1000FF2E";
        ram_buffer(19696) := X"02221004";
        ram_buffer(19697) := X"00001821";
        ram_buffer(19698) := X"1000FEAB";
        ram_buffer(19699) := X"0000B821";
        ram_buffer(19700) := X"8C820038";
        ram_buffer(19701) := X"00000000";
        ram_buffer(19702) := X"10400082";
        ram_buffer(19703) := X"00000000";
        ram_buffer(19704) := X"27BDFFC8";
        ram_buffer(19705) := X"00021043";
        ram_buffer(19706) := X"AFBF0034";
        ram_buffer(19707) := X"AFBE0030";
        ram_buffer(19708) := X"AFB7002C";
        ram_buffer(19709) := X"AFB60028";
        ram_buffer(19710) := X"AFB50024";
        ram_buffer(19711) := X"AFB40020";
        ram_buffer(19712) := X"AFB3001C";
        ram_buffer(19713) := X"AFB20018";
        ram_buffer(19714) := X"AFB10014";
        ram_buffer(19715) := X"104000F5";
        ram_buffer(19716) := X"AFB00010";
        ram_buffer(19717) := X"00008821";
        ram_buffer(19718) := X"00021043";
        ram_buffer(19719) := X"1440FFFE";
        ram_buffer(19720) := X"26310001";
        ram_buffer(19721) := X"00111900";
        ram_buffer(19722) := X"00808021";
        ram_buffer(19723) := X"8C84000C";
        ram_buffer(19724) := X"8E020034";
        ram_buffer(19725) := X"10800018";
        ram_buffer(19726) := X"00032080";
        ram_buffer(19727) := X"24420016";
        ram_buffer(19728) := X"00021080";
        ram_buffer(19729) := X"02021021";
        ram_buffer(19730) := X"8C420004";
        ram_buffer(19731) := X"00031880";
        ram_buffer(19732) := X"00431821";
        ram_buffer(19733) := X"8C620000";
        ram_buffer(19734) := X"00000000";
        ram_buffer(19735) := X"24420001";
        ram_buffer(19736) := X"AC620000";
        ram_buffer(19737) := X"8FBF0034";
        ram_buffer(19738) := X"8FBE0030";
        ram_buffer(19739) := X"8FB7002C";
        ram_buffer(19740) := X"8FB60028";
        ram_buffer(19741) := X"8FB50024";
        ram_buffer(19742) := X"8FB40020";
        ram_buffer(19743) := X"8FB3001C";
        ram_buffer(19744) := X"8FB20018";
        ram_buffer(19745) := X"8FB10014";
        ram_buffer(19746) := X"02002021";
        ram_buffer(19747) := X"8FB00010";
        ram_buffer(19748) := X"08024B01";
        ram_buffer(19749) := X"27BD0038";
        ram_buffer(19750) := X"24420012";
        ram_buffer(19751) := X"00021080";
        ram_buffer(19752) := X"02021021";
        ram_buffer(19753) := X"8C420004";
        ram_buffer(19754) := X"00000000";
        ram_buffer(19755) := X"00431821";
        ram_buffer(19756) := X"80720400";
        ram_buffer(19757) := X"00441021";
        ram_buffer(19758) := X"8C550000";
        ram_buffer(19759) := X"8E13001C";
        ram_buffer(19760) := X"124000BA";
        ram_buffer(19761) := X"24020001";
        ram_buffer(19762) := X"02421004";
        ram_buffer(19763) := X"2442FFFF";
        ram_buffer(19764) := X"00551824";
        ram_buffer(19765) := X"02539821";
        ram_buffer(19766) := X"24020018";
        ram_buffer(19767) := X"00531023";
        ram_buffer(19768) := X"8E150018";
        ram_buffer(19769) := X"00431004";
        ram_buffer(19770) := X"2A630008";
        ram_buffer(19771) := X"0055A825";
        ram_buffer(19772) := X"14600014";
        ram_buffer(19773) := X"0260B021";
        ram_buffer(19774) := X"24140016";
        ram_buffer(19775) := X"241E00FF";
        ram_buffer(19776) := X"8E030010";
        ram_buffer(19777) := X"00151403";
        ram_buffer(19778) := X"24640001";
        ram_buffer(19779) := X"AE040010";
        ram_buffer(19780) := X"A0620000";
        ram_buffer(19781) := X"8E030014";
        ram_buffer(19782) := X"26D6FFF8";
        ram_buffer(19783) := X"2463FFFF";
        ram_buffer(19784) := X"AE030014";
        ram_buffer(19785) := X"10600031";
        ram_buffer(19786) := X"305200FF";
        ram_buffer(19787) := X"125E0046";
        ram_buffer(19788) := X"00000000";
        ram_buffer(19789) := X"2AC20008";
        ram_buffer(19790) := X"1040FFF1";
        ram_buffer(19791) := X"0015AA00";
        ram_buffer(19792) := X"32730007";
        ram_buffer(19793) := X"AE150018";
        ram_buffer(19794) := X"1220FFC6";
        ram_buffer(19795) := X"AE13001C";
        ram_buffer(19796) := X"8E03000C";
        ram_buffer(19797) := X"8E040038";
        ram_buffer(19798) := X"1460FFC2";
        ram_buffer(19799) := X"24020001";
        ram_buffer(19800) := X"02221004";
        ram_buffer(19801) := X"2442FFFF";
        ram_buffer(19802) := X"02338821";
        ram_buffer(19803) := X"24030018";
        ram_buffer(19804) := X"00711823";
        ram_buffer(19805) := X"00441024";
        ram_buffer(19806) := X"00621004";
        ram_buffer(19807) := X"2A230008";
        ram_buffer(19808) := X"14600015";
        ram_buffer(19809) := X"02A2A825";
        ram_buffer(19810) := X"0220B021";
        ram_buffer(19811) := X"24130016";
        ram_buffer(19812) := X"241700FF";
        ram_buffer(19813) := X"8E030010";
        ram_buffer(19814) := X"00151403";
        ram_buffer(19815) := X"24640001";
        ram_buffer(19816) := X"AE040010";
        ram_buffer(19817) := X"A0620000";
        ram_buffer(19818) := X"8E030014";
        ram_buffer(19819) := X"26D6FFF8";
        ram_buffer(19820) := X"2463FFFF";
        ram_buffer(19821) := X"AE030014";
        ram_buffer(19822) := X"10600044";
        ram_buffer(19823) := X"305200FF";
        ram_buffer(19824) := X"12570059";
        ram_buffer(19825) := X"00000000";
        ram_buffer(19826) := X"2AC20008";
        ram_buffer(19827) := X"1040FFF1";
        ram_buffer(19828) := X"0015AA00";
        ram_buffer(19829) := X"32310007";
        ram_buffer(19830) := X"AE150018";
        ram_buffer(19831) := X"1000FFA1";
        ram_buffer(19832) := X"AE11001C";
        ram_buffer(19833) := X"03E00008";
        ram_buffer(19834) := X"00000000";
        ram_buffer(19835) := X"8E040020";
        ram_buffer(19836) := X"00000000";
        ram_buffer(19837) := X"8C970014";
        ram_buffer(19838) := X"00000000";
        ram_buffer(19839) := X"8EE2000C";
        ram_buffer(19840) := X"00000000";
        ram_buffer(19841) := X"0040F809";
        ram_buffer(19842) := X"00000000";
        ram_buffer(19843) := X"14400009";
        ram_buffer(19844) := X"00000000";
        ram_buffer(19845) := X"8E040020";
        ram_buffer(19846) := X"00000000";
        ram_buffer(19847) := X"8C820000";
        ram_buffer(19848) := X"00000000";
        ram_buffer(19849) := X"8C430000";
        ram_buffer(19850) := X"00000000";
        ram_buffer(19851) := X"0060F809";
        ram_buffer(19852) := X"AC540014";
        ram_buffer(19853) := X"8EE30000";
        ram_buffer(19854) := X"8EE20004";
        ram_buffer(19855) := X"AE030010";
        ram_buffer(19856) := X"165EFFBC";
        ram_buffer(19857) := X"AE020014";
        ram_buffer(19858) := X"8E020010";
        ram_buffer(19859) := X"00000000";
        ram_buffer(19860) := X"24430001";
        ram_buffer(19861) := X"AE030010";
        ram_buffer(19862) := X"A0400000";
        ram_buffer(19863) := X"8E020014";
        ram_buffer(19864) := X"00000000";
        ram_buffer(19865) := X"2442FFFF";
        ram_buffer(19866) := X"1440FFB2";
        ram_buffer(19867) := X"AE020014";
        ram_buffer(19868) := X"8E040020";
        ram_buffer(19869) := X"00000000";
        ram_buffer(19870) := X"8C920014";
        ram_buffer(19871) := X"00000000";
        ram_buffer(19872) := X"8E42000C";
        ram_buffer(19873) := X"00000000";
        ram_buffer(19874) := X"0040F809";
        ram_buffer(19875) := X"00000000";
        ram_buffer(19876) := X"14400009";
        ram_buffer(19877) := X"00000000";
        ram_buffer(19878) := X"8E040020";
        ram_buffer(19879) := X"00000000";
        ram_buffer(19880) := X"8C820000";
        ram_buffer(19881) := X"00000000";
        ram_buffer(19882) := X"8C430000";
        ram_buffer(19883) := X"00000000";
        ram_buffer(19884) := X"0060F809";
        ram_buffer(19885) := X"AC540014";
        ram_buffer(19886) := X"8E430000";
        ram_buffer(19887) := X"8E420004";
        ram_buffer(19888) := X"AE030010";
        ram_buffer(19889) := X"1000FF9B";
        ram_buffer(19890) := X"AE020014";
        ram_buffer(19891) := X"8E040020";
        ram_buffer(19892) := X"00000000";
        ram_buffer(19893) := X"8C940014";
        ram_buffer(19894) := X"00000000";
        ram_buffer(19895) := X"8E82000C";
        ram_buffer(19896) := X"00000000";
        ram_buffer(19897) := X"0040F809";
        ram_buffer(19898) := X"00000000";
        ram_buffer(19899) := X"14400009";
        ram_buffer(19900) := X"00000000";
        ram_buffer(19901) := X"8E040020";
        ram_buffer(19902) := X"00000000";
        ram_buffer(19903) := X"8C820000";
        ram_buffer(19904) := X"00000000";
        ram_buffer(19905) := X"8C430000";
        ram_buffer(19906) := X"00000000";
        ram_buffer(19907) := X"0060F809";
        ram_buffer(19908) := X"AC530014";
        ram_buffer(19909) := X"8E830000";
        ram_buffer(19910) := X"8E820004";
        ram_buffer(19911) := X"AE030010";
        ram_buffer(19912) := X"1657FFA9";
        ram_buffer(19913) := X"AE020014";
        ram_buffer(19914) := X"8E020010";
        ram_buffer(19915) := X"00000000";
        ram_buffer(19916) := X"24430001";
        ram_buffer(19917) := X"AE030010";
        ram_buffer(19918) := X"A0400000";
        ram_buffer(19919) := X"8E020014";
        ram_buffer(19920) := X"00000000";
        ram_buffer(19921) := X"2442FFFF";
        ram_buffer(19922) := X"1440FF9F";
        ram_buffer(19923) := X"AE020014";
        ram_buffer(19924) := X"8E040020";
        ram_buffer(19925) := X"00000000";
        ram_buffer(19926) := X"8C920014";
        ram_buffer(19927) := X"00000000";
        ram_buffer(19928) := X"8E42000C";
        ram_buffer(19929) := X"00000000";
        ram_buffer(19930) := X"0040F809";
        ram_buffer(19931) := X"00000000";
        ram_buffer(19932) := X"14400009";
        ram_buffer(19933) := X"00000000";
        ram_buffer(19934) := X"8E040020";
        ram_buffer(19935) := X"00000000";
        ram_buffer(19936) := X"8C820000";
        ram_buffer(19937) := X"00000000";
        ram_buffer(19938) := X"8C430000";
        ram_buffer(19939) := X"00000000";
        ram_buffer(19940) := X"0060F809";
        ram_buffer(19941) := X"AC530014";
        ram_buffer(19942) := X"8E430000";
        ram_buffer(19943) := X"8E420004";
        ram_buffer(19944) := X"AE030010";
        ram_buffer(19945) := X"1000FF88";
        ram_buffer(19946) := X"AE020014";
        ram_buffer(19947) := X"8E040020";
        ram_buffer(19948) := X"24050027";
        ram_buffer(19949) := X"8C820000";
        ram_buffer(19950) := X"00000000";
        ram_buffer(19951) := X"8C430000";
        ram_buffer(19952) := X"00000000";
        ram_buffer(19953) := X"0060F809";
        ram_buffer(19954) := X"AC450014";
        ram_buffer(19955) := X"8E02000C";
        ram_buffer(19956) := X"00000000";
        ram_buffer(19957) := X"1440FF23";
        ram_buffer(19958) := X"24020001";
        ram_buffer(19959) := X"1000FF3B";
        ram_buffer(19960) := X"02421004";
        ram_buffer(19961) := X"00001821";
        ram_buffer(19962) := X"1000FF0F";
        ram_buffer(19963) := X"00008821";
        ram_buffer(19964) := X"27BDFFB8";
        ram_buffer(19965) := X"AFB00020";
        ram_buffer(19966) := X"8C900164";
        ram_buffer(19967) := X"AFB20028";
        ram_buffer(19968) := X"8E020038";
        ram_buffer(19969) := X"AFBF0044";
        ram_buffer(19970) := X"AFBE0040";
        ram_buffer(19971) := X"AFB7003C";
        ram_buffer(19972) := X"AFB60038";
        ram_buffer(19973) := X"AFB50034";
        ram_buffer(19974) := X"AFB40030";
        ram_buffer(19975) := X"AFB3002C";
        ram_buffer(19976) := X"AFB10024";
        ram_buffer(19977) := X"10400019";
        ram_buffer(19978) := X"00809021";
        ram_buffer(19979) := X"00021043";
        ram_buffer(19980) := X"104001F0";
        ram_buffer(19981) := X"00001821";
        ram_buffer(19982) := X"00008821";
        ram_buffer(19983) := X"00021043";
        ram_buffer(19984) := X"1440FFFE";
        ram_buffer(19985) := X"26310001";
        ram_buffer(19986) := X"00111900";
        ram_buffer(19987) := X"8E04000C";
        ram_buffer(19988) := X"8E020034";
        ram_buffer(19989) := X"108000CE";
        ram_buffer(19990) := X"00032080";
        ram_buffer(19991) := X"24420016";
        ram_buffer(19992) := X"00021080";
        ram_buffer(19993) := X"02021021";
        ram_buffer(19994) := X"8C420004";
        ram_buffer(19995) := X"00031880";
        ram_buffer(19996) := X"00431821";
        ram_buffer(19997) := X"8C620000";
        ram_buffer(19998) := X"00000000";
        ram_buffer(19999) := X"24420001";
        ram_buffer(20000) := X"AC620000";
        ram_buffer(20001) := X"0C024B01";
        ram_buffer(20002) := X"02002021";
        ram_buffer(20003) := X"8E4200EC";
        ram_buffer(20004) := X"8E430134";
        ram_buffer(20005) := X"AFA00010";
        ram_buffer(20006) := X"AFA00014";
        ram_buffer(20007) := X"AFA00018";
        ram_buffer(20008) := X"18400031";
        ram_buffer(20009) := X"AFA0001C";
        ram_buffer(20010) := X"1060003B";
        ram_buffer(20011) := X"27B30010";
        ram_buffer(20012) := X"8E4300F0";
        ram_buffer(20013) := X"00000000";
        ram_buffer(20014) := X"8C710018";
        ram_buffer(20015) := X"00000000";
        ram_buffer(20016) := X"0011A080";
        ram_buffer(20017) := X"02741821";
        ram_buffer(20018) := X"8C630000";
        ram_buffer(20019) := X"00000000";
        ram_buffer(20020) := X"1060018F";
        ram_buffer(20021) := X"28430002";
        ram_buffer(20022) := X"14600023";
        ram_buffer(20023) := X"00000000";
        ram_buffer(20024) := X"8E4300F4";
        ram_buffer(20025) := X"00000000";
        ram_buffer(20026) := X"8C710018";
        ram_buffer(20027) := X"00000000";
        ram_buffer(20028) := X"0011A080";
        ram_buffer(20029) := X"02741821";
        ram_buffer(20030) := X"8C630000";
        ram_buffer(20031) := X"00000000";
        ram_buffer(20032) := X"106001A9";
        ram_buffer(20033) := X"28430003";
        ram_buffer(20034) := X"14600017";
        ram_buffer(20035) := X"00000000";
        ram_buffer(20036) := X"8E4300F8";
        ram_buffer(20037) := X"00000000";
        ram_buffer(20038) := X"8C710018";
        ram_buffer(20039) := X"00000000";
        ram_buffer(20040) := X"0011A080";
        ram_buffer(20041) := X"02741821";
        ram_buffer(20042) := X"8C630000";
        ram_buffer(20043) := X"00000000";
        ram_buffer(20044) := X"1060018A";
        ram_buffer(20045) := X"28420004";
        ram_buffer(20046) := X"1440000B";
        ram_buffer(20047) := X"00000000";
        ram_buffer(20048) := X"8E4200FC";
        ram_buffer(20049) := X"00000000";
        ram_buffer(20050) := X"8C510018";
        ram_buffer(20051) := X"00000000";
        ram_buffer(20052) := X"00111080";
        ram_buffer(20053) := X"02629821";
        ram_buffer(20054) := X"8E620000";
        ram_buffer(20055) := X"00000000";
        ram_buffer(20056) := X"10400119";
        ram_buffer(20057) := X"26330018";
        ram_buffer(20058) := X"8FBF0044";
        ram_buffer(20059) := X"8FBE0040";
        ram_buffer(20060) := X"8FB7003C";
        ram_buffer(20061) := X"8FB60038";
        ram_buffer(20062) := X"8FB50034";
        ram_buffer(20063) := X"8FB40030";
        ram_buffer(20064) := X"8FB3002C";
        ram_buffer(20065) := X"8FB20028";
        ram_buffer(20066) := X"8FB10024";
        ram_buffer(20067) := X"8FB00020";
        ram_buffer(20068) := X"03E00008";
        ram_buffer(20069) := X"27BD0048";
        ram_buffer(20070) := X"8E43013C";
        ram_buffer(20071) := X"8E4400F0";
        ram_buffer(20072) := X"146000CD";
        ram_buffer(20073) := X"24030001";
        ram_buffer(20074) := X"8C910014";
        ram_buffer(20075) := X"27B30010";
        ram_buffer(20076) := X"0011A880";
        ram_buffer(20077) := X"02751821";
        ram_buffer(20078) := X"8C630000";
        ram_buffer(20079) := X"00000000";
        ram_buffer(20080) := X"1460018E";
        ram_buffer(20081) := X"26340014";
        ram_buffer(20082) := X"0014A080";
        ram_buffer(20083) := X"0254A021";
        ram_buffer(20084) := X"8E850000";
        ram_buffer(20085) := X"00000000";
        ram_buffer(20086) := X"10A0019F";
        ram_buffer(20087) := X"00000000";
        ram_buffer(20088) := X"26230016";
        ram_buffer(20089) := X"00031880";
        ram_buffer(20090) := X"02031821";
        ram_buffer(20091) := X"8C660004";
        ram_buffer(20092) := X"0C024888";
        ram_buffer(20093) := X"02402021";
        ram_buffer(20094) := X"8E4200EC";
        ram_buffer(20095) := X"0275A821";
        ram_buffer(20096) := X"24040001";
        ram_buffer(20097) := X"28430002";
        ram_buffer(20098) := X"1460FFD7";
        ram_buffer(20099) := X"AEA40000";
        ram_buffer(20100) := X"8E43013C";
        ram_buffer(20101) := X"8E4400F4";
        ram_buffer(20102) := X"1460001A";
        ram_buffer(20103) := X"28430003";
        ram_buffer(20104) := X"8C910014";
        ram_buffer(20105) := X"00000000";
        ram_buffer(20106) := X"0011A880";
        ram_buffer(20107) := X"02751821";
        ram_buffer(20108) := X"8C630000";
        ram_buffer(20109) := X"00000000";
        ram_buffer(20110) := X"1460017C";
        ram_buffer(20111) := X"26340014";
        ram_buffer(20112) := X"0014A080";
        ram_buffer(20113) := X"0254A021";
        ram_buffer(20114) := X"8E850000";
        ram_buffer(20115) := X"00000000";
        ram_buffer(20116) := X"10A0018B";
        ram_buffer(20117) := X"00000000";
        ram_buffer(20118) := X"26230016";
        ram_buffer(20119) := X"00031880";
        ram_buffer(20120) := X"02031821";
        ram_buffer(20121) := X"8C660004";
        ram_buffer(20122) := X"0C024888";
        ram_buffer(20123) := X"02402021";
        ram_buffer(20124) := X"02759821";
        ram_buffer(20125) := X"24030001";
        ram_buffer(20126) := X"8E4200EC";
        ram_buffer(20127) := X"AE630000";
        ram_buffer(20128) := X"28430003";
        ram_buffer(20129) := X"1460FFB8";
        ram_buffer(20130) := X"00000000";
        ram_buffer(20131) := X"8E43013C";
        ram_buffer(20132) := X"8E4400F8";
        ram_buffer(20133) := X"1460FFB4";
        ram_buffer(20134) := X"27B30010";
        ram_buffer(20135) := X"8C910014";
        ram_buffer(20136) := X"00000000";
        ram_buffer(20137) := X"0011A880";
        ram_buffer(20138) := X"02751821";
        ram_buffer(20139) := X"8C630000";
        ram_buffer(20140) := X"00000000";
        ram_buffer(20141) := X"14600157";
        ram_buffer(20142) := X"26340014";
        ram_buffer(20143) := X"0014A080";
        ram_buffer(20144) := X"0254A021";
        ram_buffer(20145) := X"8E850000";
        ram_buffer(20146) := X"00000000";
        ram_buffer(20147) := X"10A00167";
        ram_buffer(20148) := X"00000000";
        ram_buffer(20149) := X"26230016";
        ram_buffer(20150) := X"00031880";
        ram_buffer(20151) := X"02031821";
        ram_buffer(20152) := X"8C660004";
        ram_buffer(20153) := X"0C024888";
        ram_buffer(20154) := X"02402021";
        ram_buffer(20155) := X"8E4200EC";
        ram_buffer(20156) := X"0275A821";
        ram_buffer(20157) := X"24030001";
        ram_buffer(20158) := X"28420004";
        ram_buffer(20159) := X"1440FF9A";
        ram_buffer(20160) := X"AEA30000";
        ram_buffer(20161) := X"8E42013C";
        ram_buffer(20162) := X"8E4300FC";
        ram_buffer(20163) := X"1440FF96";
        ram_buffer(20164) := X"00000000";
        ram_buffer(20165) := X"8C710014";
        ram_buffer(20166) := X"00000000";
        ram_buffer(20167) := X"00111080";
        ram_buffer(20168) := X"02629821";
        ram_buffer(20169) := X"8E620000";
        ram_buffer(20170) := X"00000000";
        ram_buffer(20171) := X"1440FF8E";
        ram_buffer(20172) := X"26330014";
        ram_buffer(20173) := X"00139880";
        ram_buffer(20174) := X"02539821";
        ram_buffer(20175) := X"8E650000";
        ram_buffer(20176) := X"00000000";
        ram_buffer(20177) := X"10A000A7";
        ram_buffer(20178) := X"00000000";
        ram_buffer(20179) := X"26310016";
        ram_buffer(20180) := X"00118880";
        ram_buffer(20181) := X"02118021";
        ram_buffer(20182) := X"8E060004";
        ram_buffer(20183) := X"8FBF0044";
        ram_buffer(20184) := X"8FBE0040";
        ram_buffer(20185) := X"8FB7003C";
        ram_buffer(20186) := X"8FB60038";
        ram_buffer(20187) := X"8FB50034";
        ram_buffer(20188) := X"8FB40030";
        ram_buffer(20189) := X"8FB3002C";
        ram_buffer(20190) := X"8FB10024";
        ram_buffer(20191) := X"8FB00020";
        ram_buffer(20192) := X"02402021";
        ram_buffer(20193) := X"8FB20028";
        ram_buffer(20194) := X"08024888";
        ram_buffer(20195) := X"27BD0048";
        ram_buffer(20196) := X"24420012";
        ram_buffer(20197) := X"00021080";
        ram_buffer(20198) := X"02021021";
        ram_buffer(20199) := X"8C420004";
        ram_buffer(20200) := X"00000000";
        ram_buffer(20201) := X"00431821";
        ram_buffer(20202) := X"80730400";
        ram_buffer(20203) := X"00441021";
        ram_buffer(20204) := X"8C560000";
        ram_buffer(20205) := X"8E14001C";
        ram_buffer(20206) := X"126000C7";
        ram_buffer(20207) := X"24020001";
        ram_buffer(20208) := X"02621004";
        ram_buffer(20209) := X"2442FFFF";
        ram_buffer(20210) := X"00561824";
        ram_buffer(20211) := X"0274A021";
        ram_buffer(20212) := X"24020018";
        ram_buffer(20213) := X"00541023";
        ram_buffer(20214) := X"8E160018";
        ram_buffer(20215) := X"00431004";
        ram_buffer(20216) := X"2A830008";
        ram_buffer(20217) := X"0056B025";
        ram_buffer(20218) := X"0280B821";
        ram_buffer(20219) := X"14600012";
        ram_buffer(20220) := X"241500FF";
        ram_buffer(20221) := X"8E030010";
        ram_buffer(20222) := X"00161403";
        ram_buffer(20223) := X"24640001";
        ram_buffer(20224) := X"AE040010";
        ram_buffer(20225) := X"A0620000";
        ram_buffer(20226) := X"8E030014";
        ram_buffer(20227) := X"26F7FFF8";
        ram_buffer(20228) := X"2463FFFF";
        ram_buffer(20229) := X"AE030014";
        ram_buffer(20230) := X"10600033";
        ram_buffer(20231) := X"305300FF";
        ram_buffer(20232) := X"12750048";
        ram_buffer(20233) := X"00000000";
        ram_buffer(20234) := X"2AE20008";
        ram_buffer(20235) := X"1040FFF1";
        ram_buffer(20236) := X"0016B200";
        ram_buffer(20237) := X"32940007";
        ram_buffer(20238) := X"AE160018";
        ram_buffer(20239) := X"1220FF11";
        ram_buffer(20240) := X"AE14001C";
        ram_buffer(20241) := X"8E03000C";
        ram_buffer(20242) := X"8E040038";
        ram_buffer(20243) := X"1460FF0D";
        ram_buffer(20244) := X"24020001";
        ram_buffer(20245) := X"02221004";
        ram_buffer(20246) := X"2442FFFF";
        ram_buffer(20247) := X"02348821";
        ram_buffer(20248) := X"24030018";
        ram_buffer(20249) := X"00711823";
        ram_buffer(20250) := X"00441024";
        ram_buffer(20251) := X"00621004";
        ram_buffer(20252) := X"2A230008";
        ram_buffer(20253) := X"14600015";
        ram_buffer(20254) := X"0056B025";
        ram_buffer(20255) := X"0220B821";
        ram_buffer(20256) := X"24140016";
        ram_buffer(20257) := X"241E00FF";
        ram_buffer(20258) := X"8E030010";
        ram_buffer(20259) := X"00161403";
        ram_buffer(20260) := X"24640001";
        ram_buffer(20261) := X"AE040010";
        ram_buffer(20262) := X"A0620000";
        ram_buffer(20263) := X"8E030014";
        ram_buffer(20264) := X"26F7FFF8";
        ram_buffer(20265) := X"2463FFFF";
        ram_buffer(20266) := X"AE030014";
        ram_buffer(20267) := X"10600052";
        ram_buffer(20268) := X"305300FF";
        ram_buffer(20269) := X"127E0067";
        ram_buffer(20270) := X"00000000";
        ram_buffer(20271) := X"2AE20008";
        ram_buffer(20272) := X"1040FFF1";
        ram_buffer(20273) := X"0016B200";
        ram_buffer(20274) := X"32310007";
        ram_buffer(20275) := X"AE160018";
        ram_buffer(20276) := X"1000FEEC";
        ram_buffer(20277) := X"AE11001C";
        ram_buffer(20278) := X"1443FF6A";
        ram_buffer(20279) := X"28430003";
        ram_buffer(20280) := X"1000FF21";
        ram_buffer(20281) := X"00000000";
        ram_buffer(20282) := X"8E040020";
        ram_buffer(20283) := X"00000000";
        ram_buffer(20284) := X"8C9E0014";
        ram_buffer(20285) := X"00000000";
        ram_buffer(20286) := X"8FC2000C";
        ram_buffer(20287) := X"00000000";
        ram_buffer(20288) := X"0040F809";
        ram_buffer(20289) := X"00000000";
        ram_buffer(20290) := X"14400009";
        ram_buffer(20291) := X"24050016";
        ram_buffer(20292) := X"8E040020";
        ram_buffer(20293) := X"00000000";
        ram_buffer(20294) := X"8C820000";
        ram_buffer(20295) := X"00000000";
        ram_buffer(20296) := X"8C430000";
        ram_buffer(20297) := X"00000000";
        ram_buffer(20298) := X"0060F809";
        ram_buffer(20299) := X"AC450014";
        ram_buffer(20300) := X"8FC30000";
        ram_buffer(20301) := X"8FC20004";
        ram_buffer(20302) := X"AE030010";
        ram_buffer(20303) := X"1675FFBA";
        ram_buffer(20304) := X"AE020014";
        ram_buffer(20305) := X"8E020010";
        ram_buffer(20306) := X"00000000";
        ram_buffer(20307) := X"24430001";
        ram_buffer(20308) := X"AE030010";
        ram_buffer(20309) := X"A0400000";
        ram_buffer(20310) := X"8E020014";
        ram_buffer(20311) := X"00000000";
        ram_buffer(20312) := X"2442FFFF";
        ram_buffer(20313) := X"1440FFB0";
        ram_buffer(20314) := X"AE020014";
        ram_buffer(20315) := X"8E040020";
        ram_buffer(20316) := X"00000000";
        ram_buffer(20317) := X"8C930014";
        ram_buffer(20318) := X"00000000";
        ram_buffer(20319) := X"8E62000C";
        ram_buffer(20320) := X"00000000";
        ram_buffer(20321) := X"0040F809";
        ram_buffer(20322) := X"00000000";
        ram_buffer(20323) := X"14400009";
        ram_buffer(20324) := X"24050016";
        ram_buffer(20325) := X"8E040020";
        ram_buffer(20326) := X"00000000";
        ram_buffer(20327) := X"8C820000";
        ram_buffer(20328) := X"00000000";
        ram_buffer(20329) := X"8C430000";
        ram_buffer(20330) := X"00000000";
        ram_buffer(20331) := X"0060F809";
        ram_buffer(20332) := X"AC450014";
        ram_buffer(20333) := X"8E630000";
        ram_buffer(20334) := X"8E620004";
        ram_buffer(20335) := X"AE030010";
        ram_buffer(20336) := X"1000FF99";
        ram_buffer(20337) := X"AE020014";
        ram_buffer(20338) := X"00139880";
        ram_buffer(20339) := X"02539821";
        ram_buffer(20340) := X"8E650000";
        ram_buffer(20341) := X"00000000";
        ram_buffer(20342) := X"14A0FF5D";
        ram_buffer(20343) := X"26310016";
        ram_buffer(20344) := X"2631FFEA";
        ram_buffer(20345) := X"0C0264A0";
        ram_buffer(20346) := X"02402021";
        ram_buffer(20347) := X"00402821";
        ram_buffer(20348) := X"1000FF56";
        ram_buffer(20349) := X"AE620000";
        ram_buffer(20350) := X"8E040020";
        ram_buffer(20351) := X"00000000";
        ram_buffer(20352) := X"8C950014";
        ram_buffer(20353) := X"00000000";
        ram_buffer(20354) := X"8EA2000C";
        ram_buffer(20355) := X"00000000";
        ram_buffer(20356) := X"0040F809";
        ram_buffer(20357) := X"00000000";
        ram_buffer(20358) := X"14400009";
        ram_buffer(20359) := X"00000000";
        ram_buffer(20360) := X"8E040020";
        ram_buffer(20361) := X"00000000";
        ram_buffer(20362) := X"8C820000";
        ram_buffer(20363) := X"00000000";
        ram_buffer(20364) := X"8C430000";
        ram_buffer(20365) := X"00000000";
        ram_buffer(20366) := X"0060F809";
        ram_buffer(20367) := X"AC540014";
        ram_buffer(20368) := X"8EA30000";
        ram_buffer(20369) := X"8EA20004";
        ram_buffer(20370) := X"AE030010";
        ram_buffer(20371) := X"167EFF9B";
        ram_buffer(20372) := X"AE020014";
        ram_buffer(20373) := X"8E020010";
        ram_buffer(20374) := X"00000000";
        ram_buffer(20375) := X"24430001";
        ram_buffer(20376) := X"AE030010";
        ram_buffer(20377) := X"A0400000";
        ram_buffer(20378) := X"8E020014";
        ram_buffer(20379) := X"00000000";
        ram_buffer(20380) := X"2442FFFF";
        ram_buffer(20381) := X"1440FF91";
        ram_buffer(20382) := X"AE020014";
        ram_buffer(20383) := X"8E040020";
        ram_buffer(20384) := X"00000000";
        ram_buffer(20385) := X"8C930014";
        ram_buffer(20386) := X"00000000";
        ram_buffer(20387) := X"8E62000C";
        ram_buffer(20388) := X"00000000";
        ram_buffer(20389) := X"0040F809";
        ram_buffer(20390) := X"00000000";
        ram_buffer(20391) := X"14400009";
        ram_buffer(20392) := X"00000000";
        ram_buffer(20393) := X"8E040020";
        ram_buffer(20394) := X"00000000";
        ram_buffer(20395) := X"8C820000";
        ram_buffer(20396) := X"00000000";
        ram_buffer(20397) := X"8C430000";
        ram_buffer(20398) := X"00000000";
        ram_buffer(20399) := X"0060F809";
        ram_buffer(20400) := X"AC540014";
        ram_buffer(20401) := X"8E630000";
        ram_buffer(20402) := X"8E620004";
        ram_buffer(20403) := X"AE030010";
        ram_buffer(20404) := X"1000FF7A";
        ram_buffer(20405) := X"AE020014";
        ram_buffer(20406) := X"8E040020";
        ram_buffer(20407) := X"24050027";
        ram_buffer(20408) := X"8C820000";
        ram_buffer(20409) := X"00000000";
        ram_buffer(20410) := X"8C430000";
        ram_buffer(20411) := X"00000000";
        ram_buffer(20412) := X"0060F809";
        ram_buffer(20413) := X"AC450014";
        ram_buffer(20414) := X"8E02000C";
        ram_buffer(20415) := X"00000000";
        ram_buffer(20416) := X"1440FE60";
        ram_buffer(20417) := X"24020001";
        ram_buffer(20418) := X"1000FF2E";
        ram_buffer(20419) := X"02621004";
        ram_buffer(20420) := X"26350018";
        ram_buffer(20421) := X"0015A880";
        ram_buffer(20422) := X"0255A821";
        ram_buffer(20423) := X"8EA50000";
        ram_buffer(20424) := X"00000000";
        ram_buffer(20425) := X"10A00060";
        ram_buffer(20426) := X"00000000";
        ram_buffer(20427) := X"26230016";
        ram_buffer(20428) := X"00031880";
        ram_buffer(20429) := X"02031821";
        ram_buffer(20430) := X"8C660004";
        ram_buffer(20431) := X"0C024888";
        ram_buffer(20432) := X"02402021";
        ram_buffer(20433) := X"0274A021";
        ram_buffer(20434) := X"24020001";
        ram_buffer(20435) := X"AE820000";
        ram_buffer(20436) := X"8E4200EC";
        ram_buffer(20437) := X"1000FE60";
        ram_buffer(20438) := X"28430002";
        ram_buffer(20439) := X"26350018";
        ram_buffer(20440) := X"0015A880";
        ram_buffer(20441) := X"0255A821";
        ram_buffer(20442) := X"8EA50000";
        ram_buffer(20443) := X"00000000";
        ram_buffer(20444) := X"10A00048";
        ram_buffer(20445) := X"00000000";
        ram_buffer(20446) := X"26230016";
        ram_buffer(20447) := X"00031880";
        ram_buffer(20448) := X"02031821";
        ram_buffer(20449) := X"8C660004";
        ram_buffer(20450) := X"0C024888";
        ram_buffer(20451) := X"02402021";
        ram_buffer(20452) := X"0274A021";
        ram_buffer(20453) := X"24020001";
        ram_buffer(20454) := X"AE820000";
        ram_buffer(20455) := X"8E4200EC";
        ram_buffer(20456) := X"1000FE65";
        ram_buffer(20457) := X"28420004";
        ram_buffer(20458) := X"26350018";
        ram_buffer(20459) := X"0015A880";
        ram_buffer(20460) := X"0255A821";
        ram_buffer(20461) := X"8EA50000";
        ram_buffer(20462) := X"00000000";
        ram_buffer(20463) := X"10A00021";
        ram_buffer(20464) := X"00000000";
        ram_buffer(20465) := X"26230016";
        ram_buffer(20466) := X"00031880";
        ram_buffer(20467) := X"02031821";
        ram_buffer(20468) := X"8C660004";
        ram_buffer(20469) := X"0C024888";
        ram_buffer(20470) := X"02402021";
        ram_buffer(20471) := X"0274A021";
        ram_buffer(20472) := X"24020001";
        ram_buffer(20473) := X"AE820000";
        ram_buffer(20474) := X"8E4200EC";
        ram_buffer(20475) := X"1000FE46";
        ram_buffer(20476) := X"28430003";
        ram_buffer(20477) := X"1000FE15";
        ram_buffer(20478) := X"00008821";
        ram_buffer(20479) := X"24030001";
        ram_buffer(20480) := X"1043FE59";
        ram_buffer(20481) := X"00000000";
        ram_buffer(20482) := X"8E4400F4";
        ram_buffer(20483) := X"1000FE84";
        ram_buffer(20484) := X"00000000";
        ram_buffer(20485) := X"24030003";
        ram_buffer(20486) := X"1043FE53";
        ram_buffer(20487) := X"00000000";
        ram_buffer(20488) := X"8E4300FC";
        ram_buffer(20489) := X"1000FEBB";
        ram_buffer(20490) := X"00000000";
        ram_buffer(20491) := X"24030002";
        ram_buffer(20492) := X"1043FE4D";
        ram_buffer(20493) := X"00000000";
        ram_buffer(20494) := X"8E4400F8";
        ram_buffer(20495) := X"1000FE97";
        ram_buffer(20496) := X"00000000";
        ram_buffer(20497) := X"0C0264A0";
        ram_buffer(20498) := X"02402021";
        ram_buffer(20499) := X"00402821";
        ram_buffer(20500) := X"1000FFDC";
        ram_buffer(20501) := X"AEA20000";
        ram_buffer(20502) := X"0C0264A0";
        ram_buffer(20503) := X"02402021";
        ram_buffer(20504) := X"00402821";
        ram_buffer(20505) := X"1000FE5E";
        ram_buffer(20506) := X"AE820000";
        ram_buffer(20507) := X"0C0264A0";
        ram_buffer(20508) := X"02402021";
        ram_buffer(20509) := X"00402821";
        ram_buffer(20510) := X"1000FE96";
        ram_buffer(20511) := X"AE820000";
        ram_buffer(20512) := X"0C0264A0";
        ram_buffer(20513) := X"02402021";
        ram_buffer(20514) := X"00402821";
        ram_buffer(20515) := X"1000FE72";
        ram_buffer(20516) := X"AE820000";
        ram_buffer(20517) := X"0C0264A0";
        ram_buffer(20518) := X"02402021";
        ram_buffer(20519) := X"00402821";
        ram_buffer(20520) := X"1000FFB5";
        ram_buffer(20521) := X"AEA20000";
        ram_buffer(20522) := X"0C0264A0";
        ram_buffer(20523) := X"02402021";
        ram_buffer(20524) := X"00402821";
        ram_buffer(20525) := X"1000FF9D";
        ram_buffer(20526) := X"AEA20000";
        ram_buffer(20527) := X"8C820038";
        ram_buffer(20528) := X"27BDFFC8";
        ram_buffer(20529) := X"AFB20018";
        ram_buffer(20530) := X"AFB00010";
        ram_buffer(20531) := X"AFBF0034";
        ram_buffer(20532) := X"AFBE0030";
        ram_buffer(20533) := X"AFB7002C";
        ram_buffer(20534) := X"AFB60028";
        ram_buffer(20535) := X"AFB50024";
        ram_buffer(20536) := X"AFB40020";
        ram_buffer(20537) := X"AFB3001C";
        ram_buffer(20538) := X"AFB10014";
        ram_buffer(20539) := X"00808021";
        ram_buffer(20540) := X"10400019";
        ram_buffer(20541) := X"00A09021";
        ram_buffer(20542) := X"00021043";
        ram_buffer(20543) := X"104001A9";
        ram_buffer(20544) := X"00001821";
        ram_buffer(20545) := X"00008821";
        ram_buffer(20546) := X"00021043";
        ram_buffer(20547) := X"1440FFFE";
        ram_buffer(20548) := X"26310001";
        ram_buffer(20549) := X"00111900";
        ram_buffer(20550) := X"8E04000C";
        ram_buffer(20551) := X"8E020034";
        ram_buffer(20552) := X"10800037";
        ram_buffer(20553) := X"00032080";
        ram_buffer(20554) := X"24420016";
        ram_buffer(20555) := X"00021080";
        ram_buffer(20556) := X"02021021";
        ram_buffer(20557) := X"8C420004";
        ram_buffer(20558) := X"00031880";
        ram_buffer(20559) := X"00431821";
        ram_buffer(20560) := X"8C620000";
        ram_buffer(20561) := X"00000000";
        ram_buffer(20562) := X"24420001";
        ram_buffer(20563) := X"AC620000";
        ram_buffer(20564) := X"0C024B01";
        ram_buffer(20565) := X"02002021";
        ram_buffer(20566) := X"8E02000C";
        ram_buffer(20567) := X"00000000";
        ram_buffer(20568) := X"104000F7";
        ram_buffer(20569) := X"24140018";
        ram_buffer(20570) := X"8E020020";
        ram_buffer(20571) := X"00000000";
        ram_buffer(20572) := X"8C430134";
        ram_buffer(20573) := X"00000000";
        ram_buffer(20574) := X"14600013";
        ram_buffer(20575) := X"00000000";
        ram_buffer(20576) := X"8C4600EC";
        ram_buffer(20577) := X"00000000";
        ram_buffer(20578) := X"18C00011";
        ram_buffer(20579) := X"26040024";
        ram_buffer(20580) := X"8FBF0034";
        ram_buffer(20581) := X"8FBE0030";
        ram_buffer(20582) := X"8FB7002C";
        ram_buffer(20583) := X"8FB60028";
        ram_buffer(20584) := X"8FB50024";
        ram_buffer(20585) := X"8FB40020";
        ram_buffer(20586) := X"8FB3001C";
        ram_buffer(20587) := X"8FB20018";
        ram_buffer(20588) := X"8FB10014";
        ram_buffer(20589) := X"8FB00010";
        ram_buffer(20590) := X"00063080";
        ram_buffer(20591) := X"00002821";
        ram_buffer(20592) := X"0802801D";
        ram_buffer(20593) := X"27BD0038";
        ram_buffer(20594) := X"AE000038";
        ram_buffer(20595) := X"AE00003C";
        ram_buffer(20596) := X"8FBF0034";
        ram_buffer(20597) := X"8FBE0030";
        ram_buffer(20598) := X"8FB7002C";
        ram_buffer(20599) := X"8FB60028";
        ram_buffer(20600) := X"8FB50024";
        ram_buffer(20601) := X"8FB40020";
        ram_buffer(20602) := X"8FB3001C";
        ram_buffer(20603) := X"8FB20018";
        ram_buffer(20604) := X"8FB10014";
        ram_buffer(20605) := X"8FB00010";
        ram_buffer(20606) := X"03E00008";
        ram_buffer(20607) := X"27BD0038";
        ram_buffer(20608) := X"24420012";
        ram_buffer(20609) := X"00021080";
        ram_buffer(20610) := X"02021021";
        ram_buffer(20611) := X"8C420004";
        ram_buffer(20612) := X"00000000";
        ram_buffer(20613) := X"00431821";
        ram_buffer(20614) := X"80730400";
        ram_buffer(20615) := X"00441021";
        ram_buffer(20616) := X"8C560000";
        ram_buffer(20617) := X"8E14001C";
        ram_buffer(20618) := X"126000B7";
        ram_buffer(20619) := X"24020001";
        ram_buffer(20620) := X"02621004";
        ram_buffer(20621) := X"2442FFFF";
        ram_buffer(20622) := X"00561824";
        ram_buffer(20623) := X"0274A021";
        ram_buffer(20624) := X"24020018";
        ram_buffer(20625) := X"00541023";
        ram_buffer(20626) := X"8E160018";
        ram_buffer(20627) := X"00431004";
        ram_buffer(20628) := X"2A830008";
        ram_buffer(20629) := X"0056B025";
        ram_buffer(20630) := X"0280B821";
        ram_buffer(20631) := X"14600012";
        ram_buffer(20632) := X"241500FF";
        ram_buffer(20633) := X"8E030010";
        ram_buffer(20634) := X"00161403";
        ram_buffer(20635) := X"24640001";
        ram_buffer(20636) := X"AE040010";
        ram_buffer(20637) := X"A0620000";
        ram_buffer(20638) := X"8E030014";
        ram_buffer(20639) := X"26F7FFF8";
        ram_buffer(20640) := X"2463FFFF";
        ram_buffer(20641) := X"AE030014";
        ram_buffer(20642) := X"1060002F";
        ram_buffer(20643) := X"305300FF";
        ram_buffer(20644) := X"12750044";
        ram_buffer(20645) := X"00000000";
        ram_buffer(20646) := X"2AE20008";
        ram_buffer(20647) := X"1040FFF1";
        ram_buffer(20648) := X"0016B200";
        ram_buffer(20649) := X"32940007";
        ram_buffer(20650) := X"AE160018";
        ram_buffer(20651) := X"1220FFA8";
        ram_buffer(20652) := X"AE14001C";
        ram_buffer(20653) := X"8E03000C";
        ram_buffer(20654) := X"8E040038";
        ram_buffer(20655) := X"1460FFA4";
        ram_buffer(20656) := X"24020001";
        ram_buffer(20657) := X"02221004";
        ram_buffer(20658) := X"2442FFFF";
        ram_buffer(20659) := X"02348821";
        ram_buffer(20660) := X"24030018";
        ram_buffer(20661) := X"00711823";
        ram_buffer(20662) := X"00441024";
        ram_buffer(20663) := X"00621004";
        ram_buffer(20664) := X"2A230008";
        ram_buffer(20665) := X"14600015";
        ram_buffer(20666) := X"0056B025";
        ram_buffer(20667) := X"0220B821";
        ram_buffer(20668) := X"24140016";
        ram_buffer(20669) := X"241E00FF";
        ram_buffer(20670) := X"8E030010";
        ram_buffer(20671) := X"00161403";
        ram_buffer(20672) := X"24640001";
        ram_buffer(20673) := X"AE040010";
        ram_buffer(20674) := X"A0620000";
        ram_buffer(20675) := X"8E030014";
        ram_buffer(20676) := X"26F7FFF8";
        ram_buffer(20677) := X"2463FFFF";
        ram_buffer(20678) := X"AE030014";
        ram_buffer(20679) := X"10600042";
        ram_buffer(20680) := X"305300FF";
        ram_buffer(20681) := X"127E0057";
        ram_buffer(20682) := X"00000000";
        ram_buffer(20683) := X"2AE20008";
        ram_buffer(20684) := X"1040FFF1";
        ram_buffer(20685) := X"0016B200";
        ram_buffer(20686) := X"32310007";
        ram_buffer(20687) := X"AE160018";
        ram_buffer(20688) := X"1000FF83";
        ram_buffer(20689) := X"AE11001C";
        ram_buffer(20690) := X"8E040020";
        ram_buffer(20691) := X"00000000";
        ram_buffer(20692) := X"8C9E0014";
        ram_buffer(20693) := X"00000000";
        ram_buffer(20694) := X"8FC2000C";
        ram_buffer(20695) := X"00000000";
        ram_buffer(20696) := X"0040F809";
        ram_buffer(20697) := X"00000000";
        ram_buffer(20698) := X"14400009";
        ram_buffer(20699) := X"24050016";
        ram_buffer(20700) := X"8E040020";
        ram_buffer(20701) := X"00000000";
        ram_buffer(20702) := X"8C820000";
        ram_buffer(20703) := X"00000000";
        ram_buffer(20704) := X"8C430000";
        ram_buffer(20705) := X"00000000";
        ram_buffer(20706) := X"0060F809";
        ram_buffer(20707) := X"AC450014";
        ram_buffer(20708) := X"8FC30000";
        ram_buffer(20709) := X"8FC20004";
        ram_buffer(20710) := X"AE030010";
        ram_buffer(20711) := X"1675FFBE";
        ram_buffer(20712) := X"AE020014";
        ram_buffer(20713) := X"8E020010";
        ram_buffer(20714) := X"00000000";
        ram_buffer(20715) := X"24430001";
        ram_buffer(20716) := X"AE030010";
        ram_buffer(20717) := X"A0400000";
        ram_buffer(20718) := X"8E020014";
        ram_buffer(20719) := X"00000000";
        ram_buffer(20720) := X"2442FFFF";
        ram_buffer(20721) := X"1440FFB4";
        ram_buffer(20722) := X"AE020014";
        ram_buffer(20723) := X"8E040020";
        ram_buffer(20724) := X"00000000";
        ram_buffer(20725) := X"8C930014";
        ram_buffer(20726) := X"00000000";
        ram_buffer(20727) := X"8E62000C";
        ram_buffer(20728) := X"00000000";
        ram_buffer(20729) := X"0040F809";
        ram_buffer(20730) := X"00000000";
        ram_buffer(20731) := X"14400009";
        ram_buffer(20732) := X"24050016";
        ram_buffer(20733) := X"8E040020";
        ram_buffer(20734) := X"00000000";
        ram_buffer(20735) := X"8C820000";
        ram_buffer(20736) := X"00000000";
        ram_buffer(20737) := X"8C430000";
        ram_buffer(20738) := X"00000000";
        ram_buffer(20739) := X"0060F809";
        ram_buffer(20740) := X"AC450014";
        ram_buffer(20741) := X"8E630000";
        ram_buffer(20742) := X"8E620004";
        ram_buffer(20743) := X"AE030010";
        ram_buffer(20744) := X"1000FF9D";
        ram_buffer(20745) := X"AE020014";
        ram_buffer(20746) := X"8E040020";
        ram_buffer(20747) := X"00000000";
        ram_buffer(20748) := X"8C950014";
        ram_buffer(20749) := X"00000000";
        ram_buffer(20750) := X"8EA2000C";
        ram_buffer(20751) := X"00000000";
        ram_buffer(20752) := X"0040F809";
        ram_buffer(20753) := X"00000000";
        ram_buffer(20754) := X"14400009";
        ram_buffer(20755) := X"00000000";
        ram_buffer(20756) := X"8E040020";
        ram_buffer(20757) := X"00000000";
        ram_buffer(20758) := X"8C820000";
        ram_buffer(20759) := X"00000000";
        ram_buffer(20760) := X"8C430000";
        ram_buffer(20761) := X"00000000";
        ram_buffer(20762) := X"0060F809";
        ram_buffer(20763) := X"AC540014";
        ram_buffer(20764) := X"8EA30000";
        ram_buffer(20765) := X"8EA20004";
        ram_buffer(20766) := X"AE030010";
        ram_buffer(20767) := X"167EFFAB";
        ram_buffer(20768) := X"AE020014";
        ram_buffer(20769) := X"8E020010";
        ram_buffer(20770) := X"00000000";
        ram_buffer(20771) := X"24430001";
        ram_buffer(20772) := X"AE030010";
        ram_buffer(20773) := X"A0400000";
        ram_buffer(20774) := X"8E020014";
        ram_buffer(20775) := X"00000000";
        ram_buffer(20776) := X"2442FFFF";
        ram_buffer(20777) := X"1440FFA1";
        ram_buffer(20778) := X"AE020014";
        ram_buffer(20779) := X"8E040020";
        ram_buffer(20780) := X"00000000";
        ram_buffer(20781) := X"8C930014";
        ram_buffer(20782) := X"00000000";
        ram_buffer(20783) := X"8E62000C";
        ram_buffer(20784) := X"00000000";
        ram_buffer(20785) := X"0040F809";
        ram_buffer(20786) := X"00000000";
        ram_buffer(20787) := X"14400009";
        ram_buffer(20788) := X"00000000";
        ram_buffer(20789) := X"8E040020";
        ram_buffer(20790) := X"00000000";
        ram_buffer(20791) := X"8C820000";
        ram_buffer(20792) := X"00000000";
        ram_buffer(20793) := X"8C430000";
        ram_buffer(20794) := X"00000000";
        ram_buffer(20795) := X"0060F809";
        ram_buffer(20796) := X"AC540014";
        ram_buffer(20797) := X"8E630000";
        ram_buffer(20798) := X"8E620004";
        ram_buffer(20799) := X"AE030010";
        ram_buffer(20800) := X"1000FF8A";
        ram_buffer(20801) := X"AE020014";
        ram_buffer(20802) := X"8E040020";
        ram_buffer(20803) := X"24050027";
        ram_buffer(20804) := X"8C820000";
        ram_buffer(20805) := X"00000000";
        ram_buffer(20806) := X"8C430000";
        ram_buffer(20807) := X"00000000";
        ram_buffer(20808) := X"0060F809";
        ram_buffer(20809) := X"AC450014";
        ram_buffer(20810) := X"8E02000C";
        ram_buffer(20811) := X"00000000";
        ram_buffer(20812) := X"1440FF07";
        ram_buffer(20813) := X"24020001";
        ram_buffer(20814) := X"1000FF3E";
        ram_buffer(20815) := X"02621004";
        ram_buffer(20816) := X"8E17001C";
        ram_buffer(20817) := X"00000000";
        ram_buffer(20818) := X"26F70007";
        ram_buffer(20819) := X"0297A023";
        ram_buffer(20820) := X"8E040018";
        ram_buffer(20821) := X"2402007F";
        ram_buffer(20822) := X"02821004";
        ram_buffer(20823) := X"2AE30008";
        ram_buffer(20824) := X"14600092";
        ram_buffer(20825) := X"0044A025";
        ram_buffer(20826) := X"8E030010";
        ram_buffer(20827) := X"24130016";
        ram_buffer(20828) := X"241600FF";
        ram_buffer(20829) := X"00141403";
        ram_buffer(20830) := X"24640001";
        ram_buffer(20831) := X"AE040010";
        ram_buffer(20832) := X"A0620000";
        ram_buffer(20833) := X"8E030014";
        ram_buffer(20834) := X"305100FF";
        ram_buffer(20835) := X"2462FFFF";
        ram_buffer(20836) := X"10400035";
        ram_buffer(20837) := X"AE020014";
        ram_buffer(20838) := X"8E030010";
        ram_buffer(20839) := X"1236004A";
        ram_buffer(20840) := X"24620001";
        ram_buffer(20841) := X"26F7FFF8";
        ram_buffer(20842) := X"2AE20008";
        ram_buffer(20843) := X"1040FFF1";
        ram_buffer(20844) := X"0014A200";
        ram_buffer(20845) := X"24620001";
        ram_buffer(20846) := X"AE020010";
        ram_buffer(20847) := X"2402FFFF";
        ram_buffer(20848) := X"AE000018";
        ram_buffer(20849) := X"AE00001C";
        ram_buffer(20850) := X"A0620000";
        ram_buffer(20851) := X"8E020014";
        ram_buffer(20852) := X"00000000";
        ram_buffer(20853) := X"2442FFFF";
        ram_buffer(20854) := X"1040005C";
        ram_buffer(20855) := X"AE020014";
        ram_buffer(20856) := X"8E020010";
        ram_buffer(20857) := X"00000000";
        ram_buffer(20858) := X"24430001";
        ram_buffer(20859) := X"2652FFD0";
        ram_buffer(20860) := X"AE030010";
        ram_buffer(20861) := X"A0520000";
        ram_buffer(20862) := X"8E020014";
        ram_buffer(20863) := X"00000000";
        ram_buffer(20864) := X"2442FFFF";
        ram_buffer(20865) := X"1440FED8";
        ram_buffer(20866) := X"AE020014";
        ram_buffer(20867) := X"8E040020";
        ram_buffer(20868) := X"00000000";
        ram_buffer(20869) := X"8C910014";
        ram_buffer(20870) := X"00000000";
        ram_buffer(20871) := X"8E22000C";
        ram_buffer(20872) := X"00000000";
        ram_buffer(20873) := X"0040F809";
        ram_buffer(20874) := X"00000000";
        ram_buffer(20875) := X"14400009";
        ram_buffer(20876) := X"24050016";
        ram_buffer(20877) := X"8E040020";
        ram_buffer(20878) := X"00000000";
        ram_buffer(20879) := X"8C820000";
        ram_buffer(20880) := X"00000000";
        ram_buffer(20881) := X"8C430000";
        ram_buffer(20882) := X"00000000";
        ram_buffer(20883) := X"0060F809";
        ram_buffer(20884) := X"AC450014";
        ram_buffer(20885) := X"8E230000";
        ram_buffer(20886) := X"8E220004";
        ram_buffer(20887) := X"AE030010";
        ram_buffer(20888) := X"1000FEC1";
        ram_buffer(20889) := X"AE020014";
        ram_buffer(20890) := X"8E040020";
        ram_buffer(20891) := X"00000000";
        ram_buffer(20892) := X"8C950014";
        ram_buffer(20893) := X"00000000";
        ram_buffer(20894) := X"8EA2000C";
        ram_buffer(20895) := X"00000000";
        ram_buffer(20896) := X"0040F809";
        ram_buffer(20897) := X"00000000";
        ram_buffer(20898) := X"14400009";
        ram_buffer(20899) := X"00000000";
        ram_buffer(20900) := X"8E040020";
        ram_buffer(20901) := X"00000000";
        ram_buffer(20902) := X"8C820000";
        ram_buffer(20903) := X"00000000";
        ram_buffer(20904) := X"8C430000";
        ram_buffer(20905) := X"00000000";
        ram_buffer(20906) := X"0060F809";
        ram_buffer(20907) := X"AC530014";
        ram_buffer(20908) := X"8EA30000";
        ram_buffer(20909) := X"8EA20004";
        ram_buffer(20910) := X"AE030010";
        ram_buffer(20911) := X"1636FFB9";
        ram_buffer(20912) := X"AE020014";
        ram_buffer(20913) := X"24620001";
        ram_buffer(20914) := X"AE020010";
        ram_buffer(20915) := X"A0600000";
        ram_buffer(20916) := X"8E020014";
        ram_buffer(20917) := X"00000000";
        ram_buffer(20918) := X"2442FFFF";
        ram_buffer(20919) := X"10400004";
        ram_buffer(20920) := X"AE020014";
        ram_buffer(20921) := X"8E030010";
        ram_buffer(20922) := X"1000FFAF";
        ram_buffer(20923) := X"26F7FFF8";
        ram_buffer(20924) := X"8E040020";
        ram_buffer(20925) := X"00000000";
        ram_buffer(20926) := X"8C910014";
        ram_buffer(20927) := X"00000000";
        ram_buffer(20928) := X"8E22000C";
        ram_buffer(20929) := X"00000000";
        ram_buffer(20930) := X"0040F809";
        ram_buffer(20931) := X"00000000";
        ram_buffer(20932) := X"14400009";
        ram_buffer(20933) := X"00000000";
        ram_buffer(20934) := X"8E040020";
        ram_buffer(20935) := X"00000000";
        ram_buffer(20936) := X"8C820000";
        ram_buffer(20937) := X"00000000";
        ram_buffer(20938) := X"8C430000";
        ram_buffer(20939) := X"00000000";
        ram_buffer(20940) := X"0060F809";
        ram_buffer(20941) := X"AC530014";
        ram_buffer(20942) := X"8E230000";
        ram_buffer(20943) := X"8E220004";
        ram_buffer(20944) := X"AE030010";
        ram_buffer(20945) := X"1000FF97";
        ram_buffer(20946) := X"AE020014";
        ram_buffer(20947) := X"8E040020";
        ram_buffer(20948) := X"00000000";
        ram_buffer(20949) := X"8C910014";
        ram_buffer(20950) := X"00000000";
        ram_buffer(20951) := X"8E22000C";
        ram_buffer(20952) := X"00000000";
        ram_buffer(20953) := X"0040F809";
        ram_buffer(20954) := X"00000000";
        ram_buffer(20955) := X"14400009";
        ram_buffer(20956) := X"24050016";
        ram_buffer(20957) := X"8E040020";
        ram_buffer(20958) := X"00000000";
        ram_buffer(20959) := X"8C820000";
        ram_buffer(20960) := X"00000000";
        ram_buffer(20961) := X"8C430000";
        ram_buffer(20962) := X"00000000";
        ram_buffer(20963) := X"0060F809";
        ram_buffer(20964) := X"AC450014";
        ram_buffer(20965) := X"8E230004";
        ram_buffer(20966) := X"8E220000";
        ram_buffer(20967) := X"1000FF92";
        ram_buffer(20968) := X"AE030014";
        ram_buffer(20969) := X"1000FE5C";
        ram_buffer(20970) := X"00008821";
        ram_buffer(20971) := X"8E030010";
        ram_buffer(20972) := X"1000FF81";
        ram_buffer(20973) := X"24620001";
        ram_buffer(20974) := X"27BDFFB0";
        ram_buffer(20975) := X"8C820014";
        ram_buffer(20976) := X"AFB5003C";
        ram_buffer(20977) := X"0080A821";
        ram_buffer(20978) := X"AFBE0048";
        ram_buffer(20979) := X"8C460000";
        ram_buffer(20980) := X"8C9E0164";
        ram_buffer(20981) := X"8EA30140";
        ram_buffer(20982) := X"8C440004";
        ram_buffer(20983) := X"8EA200C0";
        ram_buffer(20984) := X"AFB20030";
        ram_buffer(20985) := X"AFBF004C";
        ram_buffer(20986) := X"AFB70044";
        ram_buffer(20987) := X"AFB60040";
        ram_buffer(20988) := X"AFB40038";
        ram_buffer(20989) := X"AFB30034";
        ram_buffer(20990) := X"AFB1002C";
        ram_buffer(20991) := X"AFB00028";
        ram_buffer(20992) := X"AFA30020";
        ram_buffer(20993) := X"00A09021";
        ram_buffer(20994) := X"AFC60010";
        ram_buffer(20995) := X"10400005";
        ram_buffer(20996) := X"AFC40014";
        ram_buffer(20997) := X"8FC20044";
        ram_buffer(20998) := X"00000000";
        ram_buffer(20999) := X"1040013F";
        ram_buffer(21000) := X"00000000";
        ram_buffer(21001) := X"8EA20108";
        ram_buffer(21002) := X"00000000";
        ram_buffer(21003) := X"1840002E";
        ram_buffer(21004) := X"00000000";
        ram_buffer(21005) := X"26B4010C";
        ram_buffer(21006) := X"00009821";
        ram_buffer(21007) := X"241100FF";
        ram_buffer(21008) := X"8E840000";
        ram_buffer(21009) := X"8E420000";
        ram_buffer(21010) := X"00042880";
        ram_buffer(21011) := X"84460000";
        ram_buffer(21012) := X"03C52821";
        ram_buffer(21013) := X"8FA30020";
        ram_buffer(21014) := X"8CA20024";
        ram_buffer(21015) := X"2484003C";
        ram_buffer(21016) := X"00663007";
        ram_buffer(21017) := X"00042080";
        ram_buffer(21018) := X"02A42021";
        ram_buffer(21019) := X"00C21023";
        ram_buffer(21020) := X"8C870000";
        ram_buffer(21021) := X"0440010E";
        ram_buffer(21022) := X"ACA60024";
        ram_buffer(21023) := X"1040011E";
        ram_buffer(21024) := X"00000000";
        ram_buffer(21025) := X"AFA20018";
        ram_buffer(21026) := X"0000B821";
        ram_buffer(21027) := X"00021043";
        ram_buffer(21028) := X"1440FFFE";
        ram_buffer(21029) := X"26F70001";
        ram_buffer(21030) := X"8FC4000C";
        ram_buffer(21031) := X"8CE20014";
        ram_buffer(21032) := X"1080002B";
        ram_buffer(21033) := X"00172880";
        ram_buffer(21034) := X"24420016";
        ram_buffer(21035) := X"00021080";
        ram_buffer(21036) := X"03C21021";
        ram_buffer(21037) := X"8C420004";
        ram_buffer(21038) := X"00000000";
        ram_buffer(21039) := X"00452821";
        ram_buffer(21040) := X"8CA20000";
        ram_buffer(21041) := X"00000000";
        ram_buffer(21042) := X"24420001";
        ram_buffer(21043) := X"ACA20000";
        ram_buffer(21044) := X"8EA20108";
        ram_buffer(21045) := X"26730001";
        ram_buffer(21046) := X"0262102A";
        ram_buffer(21047) := X"26520004";
        ram_buffer(21048) := X"1440FFD7";
        ram_buffer(21049) := X"26940004";
        ram_buffer(21050) := X"8EA20014";
        ram_buffer(21051) := X"8FC60010";
        ram_buffer(21052) := X"8FC50014";
        ram_buffer(21053) := X"8EA400C0";
        ram_buffer(21054) := X"AC460000";
        ram_buffer(21055) := X"10800007";
        ram_buffer(21056) := X"AC450004";
        ram_buffer(21057) := X"8FC20044";
        ram_buffer(21058) := X"00000000";
        ram_buffer(21059) := X"104000FD";
        ram_buffer(21060) := X"00000000";
        ram_buffer(21061) := X"2442FFFF";
        ram_buffer(21062) := X"AFC20044";
        ram_buffer(21063) := X"8FBF004C";
        ram_buffer(21064) := X"8FBE0048";
        ram_buffer(21065) := X"8FB70044";
        ram_buffer(21066) := X"8FB60040";
        ram_buffer(21067) := X"8FB5003C";
        ram_buffer(21068) := X"8FB40038";
        ram_buffer(21069) := X"8FB30034";
        ram_buffer(21070) := X"8FB20030";
        ram_buffer(21071) := X"8FB1002C";
        ram_buffer(21072) := X"8FB00028";
        ram_buffer(21073) := X"24020001";
        ram_buffer(21074) := X"03E00008";
        ram_buffer(21075) := X"27BD0050";
        ram_buffer(21076) := X"24420012";
        ram_buffer(21077) := X"00021080";
        ram_buffer(21078) := X"03C21021";
        ram_buffer(21079) := X"8C420004";
        ram_buffer(21080) := X"00172080";
        ram_buffer(21081) := X"00573021";
        ram_buffer(21082) := X"80D00400";
        ram_buffer(21083) := X"00441021";
        ram_buffer(21084) := X"8C560000";
        ram_buffer(21085) := X"8FC6001C";
        ram_buffer(21086) := X"120000D1";
        ram_buffer(21087) := X"24020001";
        ram_buffer(21088) := X"02021004";
        ram_buffer(21089) := X"02061821";
        ram_buffer(21090) := X"24040018";
        ram_buffer(21091) := X"2442FFFF";
        ram_buffer(21092) := X"00561024";
        ram_buffer(21093) := X"00833823";
        ram_buffer(21094) := X"8FC60018";
        ram_buffer(21095) := X"00E21004";
        ram_buffer(21096) := X"28640008";
        ram_buffer(21097) := X"0046B025";
        ram_buffer(21098) := X"AFA3001C";
        ram_buffer(21099) := X"00608021";
        ram_buffer(21100) := X"14800015";
        ram_buffer(21101) := X"00601021";
        ram_buffer(21102) := X"8FC40010";
        ram_buffer(21103) := X"00161403";
        ram_buffer(21104) := X"24860001";
        ram_buffer(21105) := X"AFC60010";
        ram_buffer(21106) := X"A0820000";
        ram_buffer(21107) := X"8FC40014";
        ram_buffer(21108) := X"2610FFF8";
        ram_buffer(21109) := X"2484FFFF";
        ram_buffer(21110) := X"AFC40014";
        ram_buffer(21111) := X"1080003A";
        ram_buffer(21112) := X"304600FF";
        ram_buffer(21113) := X"10D10053";
        ram_buffer(21114) := X"00000000";
        ram_buffer(21115) := X"2A020008";
        ram_buffer(21116) := X"1040FFF1";
        ram_buffer(21117) := X"0016B200";
        ram_buffer(21118) := X"8FA2001C";
        ram_buffer(21119) := X"00000000";
        ram_buffer(21120) := X"30420007";
        ram_buffer(21121) := X"AFA2001C";
        ram_buffer(21122) := X"AFD60018";
        ram_buffer(21123) := X"12E0FFB0";
        ram_buffer(21124) := X"AFC2001C";
        ram_buffer(21125) := X"8FC2000C";
        ram_buffer(21126) := X"00000000";
        ram_buffer(21127) := X"1440FFAC";
        ram_buffer(21128) := X"24020001";
        ram_buffer(21129) := X"8FA3001C";
        ram_buffer(21130) := X"00000000";
        ram_buffer(21131) := X"02E31821";
        ram_buffer(21132) := X"00602021";
        ram_buffer(21133) := X"02E21004";
        ram_buffer(21134) := X"AFA30014";
        ram_buffer(21135) := X"8FA30018";
        ram_buffer(21136) := X"2442FFFF";
        ram_buffer(21137) := X"24050018";
        ram_buffer(21138) := X"00431824";
        ram_buffer(21139) := X"00A41023";
        ram_buffer(21140) := X"00431004";
        ram_buffer(21141) := X"00801821";
        ram_buffer(21142) := X"28840008";
        ram_buffer(21143) := X"14800016";
        ram_buffer(21144) := X"0056B825";
        ram_buffer(21145) := X"00608021";
        ram_buffer(21146) := X"8FC40010";
        ram_buffer(21147) := X"00171403";
        ram_buffer(21148) := X"24860001";
        ram_buffer(21149) := X"AFC60010";
        ram_buffer(21150) := X"A0820000";
        ram_buffer(21151) := X"8FC40014";
        ram_buffer(21152) := X"2610FFF8";
        ram_buffer(21153) := X"2484FFFF";
        ram_buffer(21154) := X"AFC40014";
        ram_buffer(21155) := X"1080004D";
        ram_buffer(21156) := X"305600FF";
        ram_buffer(21157) := X"12D10065";
        ram_buffer(21158) := X"00000000";
        ram_buffer(21159) := X"2A020008";
        ram_buffer(21160) := X"1040FFF1";
        ram_buffer(21161) := X"0017BA00";
        ram_buffer(21162) := X"8FA20014";
        ram_buffer(21163) := X"00000000";
        ram_buffer(21164) := X"30420007";
        ram_buffer(21165) := X"AFA20014";
        ram_buffer(21166) := X"8FA20014";
        ram_buffer(21167) := X"AFD70018";
        ram_buffer(21168) := X"1000FF83";
        ram_buffer(21169) := X"AFC2001C";
        ram_buffer(21170) := X"8FC40020";
        ram_buffer(21171) := X"AFA60014";
        ram_buffer(21172) := X"8C890014";
        ram_buffer(21173) := X"00000000";
        ram_buffer(21174) := X"8D22000C";
        ram_buffer(21175) := X"00000000";
        ram_buffer(21176) := X"0040F809";
        ram_buffer(21177) := X"AFA90010";
        ram_buffer(21178) := X"8FA90010";
        ram_buffer(21179) := X"8FA60014";
        ram_buffer(21180) := X"1440000B";
        ram_buffer(21181) := X"24030016";
        ram_buffer(21182) := X"8FC40020";
        ram_buffer(21183) := X"00000000";
        ram_buffer(21184) := X"8C820000";
        ram_buffer(21185) := X"AFA90014";
        ram_buffer(21186) := X"8C4A0000";
        ram_buffer(21187) := X"AC430014";
        ram_buffer(21188) := X"0140F809";
        ram_buffer(21189) := X"AFA60010";
        ram_buffer(21190) := X"8FA90014";
        ram_buffer(21191) := X"8FA60010";
        ram_buffer(21192) := X"8D240000";
        ram_buffer(21193) := X"8D220004";
        ram_buffer(21194) := X"AFC40010";
        ram_buffer(21195) := X"14D1FFAF";
        ram_buffer(21196) := X"AFC20014";
        ram_buffer(21197) := X"8FC20010";
        ram_buffer(21198) := X"00000000";
        ram_buffer(21199) := X"24440001";
        ram_buffer(21200) := X"AFC40010";
        ram_buffer(21201) := X"A0400000";
        ram_buffer(21202) := X"8FC20014";
        ram_buffer(21203) := X"00000000";
        ram_buffer(21204) := X"2442FFFF";
        ram_buffer(21205) := X"1440FFA5";
        ram_buffer(21206) := X"AFC20014";
        ram_buffer(21207) := X"8FC40020";
        ram_buffer(21208) := X"00000000";
        ram_buffer(21209) := X"8C860014";
        ram_buffer(21210) := X"00000000";
        ram_buffer(21211) := X"8CC2000C";
        ram_buffer(21212) := X"00000000";
        ram_buffer(21213) := X"0040F809";
        ram_buffer(21214) := X"AFA60010";
        ram_buffer(21215) := X"8FA60010";
        ram_buffer(21216) := X"1440000B";
        ram_buffer(21217) := X"00000000";
        ram_buffer(21218) := X"8FC40020";
        ram_buffer(21219) := X"24030016";
        ram_buffer(21220) := X"8C820000";
        ram_buffer(21221) := X"00000000";
        ram_buffer(21222) := X"8C490000";
        ram_buffer(21223) := X"00000000";
        ram_buffer(21224) := X"0120F809";
        ram_buffer(21225) := X"AC430014";
        ram_buffer(21226) := X"8FA60010";
        ram_buffer(21227) := X"00000000";
        ram_buffer(21228) := X"8CC40000";
        ram_buffer(21229) := X"8CC20004";
        ram_buffer(21230) := X"AFC40010";
        ram_buffer(21231) := X"1000FF8B";
        ram_buffer(21232) := X"AFC20014";
        ram_buffer(21233) := X"8FC40020";
        ram_buffer(21234) := X"00000000";
        ram_buffer(21235) := X"8C860014";
        ram_buffer(21236) := X"00000000";
        ram_buffer(21237) := X"8CC2000C";
        ram_buffer(21238) := X"00000000";
        ram_buffer(21239) := X"0040F809";
        ram_buffer(21240) := X"AFA60010";
        ram_buffer(21241) := X"8FA60010";
        ram_buffer(21242) := X"1440000B";
        ram_buffer(21243) := X"24030016";
        ram_buffer(21244) := X"8FC40020";
        ram_buffer(21245) := X"00000000";
        ram_buffer(21246) := X"8C820000";
        ram_buffer(21247) := X"00000000";
        ram_buffer(21248) := X"8C480000";
        ram_buffer(21249) := X"00000000";
        ram_buffer(21250) := X"0100F809";
        ram_buffer(21251) := X"AC430014";
        ram_buffer(21252) := X"8FA60010";
        ram_buffer(21253) := X"00000000";
        ram_buffer(21254) := X"8CC40000";
        ram_buffer(21255) := X"8CC20004";
        ram_buffer(21256) := X"AFC40010";
        ram_buffer(21257) := X"16D1FF9D";
        ram_buffer(21258) := X"AFC20014";
        ram_buffer(21259) := X"8FC20010";
        ram_buffer(21260) := X"00000000";
        ram_buffer(21261) := X"24440001";
        ram_buffer(21262) := X"AFC40010";
        ram_buffer(21263) := X"A0400000";
        ram_buffer(21264) := X"8FC20014";
        ram_buffer(21265) := X"00000000";
        ram_buffer(21266) := X"2442FFFF";
        ram_buffer(21267) := X"1440FF93";
        ram_buffer(21268) := X"AFC20014";
        ram_buffer(21269) := X"8FC40020";
        ram_buffer(21270) := X"00000000";
        ram_buffer(21271) := X"8C960014";
        ram_buffer(21272) := X"00000000";
        ram_buffer(21273) := X"8EC2000C";
        ram_buffer(21274) := X"00000000";
        ram_buffer(21275) := X"0040F809";
        ram_buffer(21276) := X"00000000";
        ram_buffer(21277) := X"14400009";
        ram_buffer(21278) := X"24030016";
        ram_buffer(21279) := X"8FC40020";
        ram_buffer(21280) := X"00000000";
        ram_buffer(21281) := X"8C820000";
        ram_buffer(21282) := X"00000000";
        ram_buffer(21283) := X"8C460000";
        ram_buffer(21284) := X"00000000";
        ram_buffer(21285) := X"00C0F809";
        ram_buffer(21286) := X"AC430014";
        ram_buffer(21287) := X"8EC40000";
        ram_buffer(21288) := X"8EC20004";
        ram_buffer(21289) := X"AFC40010";
        ram_buffer(21290) := X"1000FF7C";
        ram_buffer(21291) := X"AFC20014";
        ram_buffer(21292) := X"2443FFFF";
        ram_buffer(21293) := X"AFA30018";
        ram_buffer(21294) := X"1000FEF3";
        ram_buffer(21295) := X"00021023";
        ram_buffer(21296) := X"8FC40020";
        ram_buffer(21297) := X"24030027";
        ram_buffer(21298) := X"8C820000";
        ram_buffer(21299) := X"AFA60010";
        ram_buffer(21300) := X"8C480000";
        ram_buffer(21301) := X"00000000";
        ram_buffer(21302) := X"0100F809";
        ram_buffer(21303) := X"AC430014";
        ram_buffer(21304) := X"8FC2000C";
        ram_buffer(21305) := X"8FA60010";
        ram_buffer(21306) := X"1440FEF9";
        ram_buffer(21307) := X"24020001";
        ram_buffer(21308) := X"1000FF24";
        ram_buffer(21309) := X"02021004";
        ram_buffer(21310) := X"AFA00018";
        ram_buffer(21311) := X"1000FEE6";
        ram_buffer(21312) := X"0000B821";
        ram_buffer(21313) := X"8FC50048";
        ram_buffer(21314) := X"00801021";
        ram_buffer(21315) := X"24A40001";
        ram_buffer(21316) := X"30840007";
        ram_buffer(21317) := X"1000FEFF";
        ram_buffer(21318) := X"AFC40048";
        ram_buffer(21319) := X"8FC50048";
        ram_buffer(21320) := X"0C02502F";
        ram_buffer(21321) := X"03C02021";
        ram_buffer(21322) := X"1000FEBE";
        ram_buffer(21323) := X"00000000";
        ram_buffer(21324) := X"8C820014";
        ram_buffer(21325) := X"27BDFFC0";
        ram_buffer(21326) := X"00801821";
        ram_buffer(21327) := X"8C460004";
        ram_buffer(21328) := X"AFB70034";
        ram_buffer(21329) := X"AFA40040";
        ram_buffer(21330) := X"8C970164";
        ram_buffer(21331) := X"8C440000";
        ram_buffer(21332) := X"8C6200C0";
        ram_buffer(21333) := X"8C630140";
        ram_buffer(21334) := X"AFB20020";
        ram_buffer(21335) := X"AFBF003C";
        ram_buffer(21336) := X"AFBE0038";
        ram_buffer(21337) := X"AFB60030";
        ram_buffer(21338) := X"AFB5002C";
        ram_buffer(21339) := X"AFB40028";
        ram_buffer(21340) := X"AFB30024";
        ram_buffer(21341) := X"AFB1001C";
        ram_buffer(21342) := X"AFB00018";
        ram_buffer(21343) := X"AFA30010";
        ram_buffer(21344) := X"00A09021";
        ram_buffer(21345) := X"AEE40010";
        ram_buffer(21346) := X"10400005";
        ram_buffer(21347) := X"AEE60014";
        ram_buffer(21348) := X"8EE20044";
        ram_buffer(21349) := X"00000000";
        ram_buffer(21350) := X"1040008F";
        ram_buffer(21351) := X"00000000";
        ram_buffer(21352) := X"8FA20040";
        ram_buffer(21353) := X"00000000";
        ram_buffer(21354) := X"8C470108";
        ram_buffer(21355) := X"00000000";
        ram_buffer(21356) := X"18E00030";
        ram_buffer(21357) := X"00000000";
        ram_buffer(21358) := X"8EF3001C";
        ram_buffer(21359) := X"00008821";
        ram_buffer(21360) := X"241000FF";
        ram_buffer(21361) := X"8EE2000C";
        ram_buffer(21362) := X"00000000";
        ram_buffer(21363) := X"14400024";
        ram_buffer(21364) := X"26760001";
        ram_buffer(21365) := X"8E420000";
        ram_buffer(21366) := X"24030018";
        ram_buffer(21367) := X"00762823";
        ram_buffer(21368) := X"84420000";
        ram_buffer(21369) := X"8FA30010";
        ram_buffer(21370) := X"8EE90018";
        ram_buffer(21371) := X"00621007";
        ram_buffer(21372) := X"30420001";
        ram_buffer(21373) := X"00A21004";
        ram_buffer(21374) := X"2AC80008";
        ram_buffer(21375) := X"15000015";
        ram_buffer(21376) := X"0049A825";
        ram_buffer(21377) := X"00151403";
        ram_buffer(21378) := X"24870001";
        ram_buffer(21379) := X"AEE70010";
        ram_buffer(21380) := X"A0820000";
        ram_buffer(21381) := X"8EE40014";
        ram_buffer(21382) := X"305E00FF";
        ram_buffer(21383) := X"2482FFFF";
        ram_buffer(21384) := X"1040002E";
        ram_buffer(21385) := X"AEE20014";
        ram_buffer(21386) := X"8EE40010";
        ram_buffer(21387) := X"13D00043";
        ram_buffer(21388) := X"24820001";
        ram_buffer(21389) := X"26D6FFF8";
        ram_buffer(21390) := X"2AC20008";
        ram_buffer(21391) := X"1040FFF1";
        ram_buffer(21392) := X"0015AA00";
        ram_buffer(21393) := X"8FA20040";
        ram_buffer(21394) := X"2673FFF9";
        ram_buffer(21395) := X"8C470108";
        ram_buffer(21396) := X"32760007";
        ram_buffer(21397) := X"AEF50018";
        ram_buffer(21398) := X"AEF6001C";
        ram_buffer(21399) := X"02C09821";
        ram_buffer(21400) := X"26310001";
        ram_buffer(21401) := X"0227102A";
        ram_buffer(21402) := X"1440FFD6";
        ram_buffer(21403) := X"26520004";
        ram_buffer(21404) := X"8FA20040";
        ram_buffer(21405) := X"8FA30040";
        ram_buffer(21406) := X"8C420014";
        ram_buffer(21407) := X"8EE60014";
        ram_buffer(21408) := X"8C6500C0";
        ram_buffer(21409) := X"AC440000";
        ram_buffer(21410) := X"10A00007";
        ram_buffer(21411) := X"AC460004";
        ram_buffer(21412) := X"8EE20044";
        ram_buffer(21413) := X"00000000";
        ram_buffer(21414) := X"10400049";
        ram_buffer(21415) := X"00000000";
        ram_buffer(21416) := X"2442FFFF";
        ram_buffer(21417) := X"AEE20044";
        ram_buffer(21418) := X"8FBF003C";
        ram_buffer(21419) := X"8FBE0038";
        ram_buffer(21420) := X"8FB70034";
        ram_buffer(21421) := X"8FB60030";
        ram_buffer(21422) := X"8FB5002C";
        ram_buffer(21423) := X"8FB40028";
        ram_buffer(21424) := X"8FB30024";
        ram_buffer(21425) := X"8FB20020";
        ram_buffer(21426) := X"8FB1001C";
        ram_buffer(21427) := X"8FB00018";
        ram_buffer(21428) := X"24020001";
        ram_buffer(21429) := X"03E00008";
        ram_buffer(21430) := X"27BD0040";
        ram_buffer(21431) := X"8EE40020";
        ram_buffer(21432) := X"00000000";
        ram_buffer(21433) := X"8C940014";
        ram_buffer(21434) := X"00000000";
        ram_buffer(21435) := X"8E82000C";
        ram_buffer(21436) := X"00000000";
        ram_buffer(21437) := X"0040F809";
        ram_buffer(21438) := X"00000000";
        ram_buffer(21439) := X"14400009";
        ram_buffer(21440) := X"24030016";
        ram_buffer(21441) := X"8EE40020";
        ram_buffer(21442) := X"00000000";
        ram_buffer(21443) := X"8C820000";
        ram_buffer(21444) := X"00000000";
        ram_buffer(21445) := X"8C480000";
        ram_buffer(21446) := X"00000000";
        ram_buffer(21447) := X"0100F809";
        ram_buffer(21448) := X"AC430014";
        ram_buffer(21449) := X"8E840000";
        ram_buffer(21450) := X"8E820004";
        ram_buffer(21451) := X"AEE40010";
        ram_buffer(21452) := X"17D0FFC0";
        ram_buffer(21453) := X"AEE20014";
        ram_buffer(21454) := X"24820001";
        ram_buffer(21455) := X"AEE20010";
        ram_buffer(21456) := X"A0800000";
        ram_buffer(21457) := X"8EE20014";
        ram_buffer(21458) := X"00000000";
        ram_buffer(21459) := X"2442FFFF";
        ram_buffer(21460) := X"10400004";
        ram_buffer(21461) := X"AEE20014";
        ram_buffer(21462) := X"8EE40010";
        ram_buffer(21463) := X"1000FFB6";
        ram_buffer(21464) := X"26D6FFF8";
        ram_buffer(21465) := X"8EE40020";
        ram_buffer(21466) := X"00000000";
        ram_buffer(21467) := X"8C9E0014";
        ram_buffer(21468) := X"00000000";
        ram_buffer(21469) := X"8FC2000C";
        ram_buffer(21470) := X"00000000";
        ram_buffer(21471) := X"0040F809";
        ram_buffer(21472) := X"00000000";
        ram_buffer(21473) := X"14400009";
        ram_buffer(21474) := X"24030016";
        ram_buffer(21475) := X"8EE40020";
        ram_buffer(21476) := X"00000000";
        ram_buffer(21477) := X"8C820000";
        ram_buffer(21478) := X"00000000";
        ram_buffer(21479) := X"8C470000";
        ram_buffer(21480) := X"00000000";
        ram_buffer(21481) := X"00E0F809";
        ram_buffer(21482) := X"AC430014";
        ram_buffer(21483) := X"8FC40000";
        ram_buffer(21484) := X"8FC20004";
        ram_buffer(21485) := X"AEE40010";
        ram_buffer(21486) := X"1000FF9E";
        ram_buffer(21487) := X"AEE20014";
        ram_buffer(21488) := X"8EE40048";
        ram_buffer(21489) := X"00A01021";
        ram_buffer(21490) := X"24840001";
        ram_buffer(21491) := X"30840007";
        ram_buffer(21492) := X"1000FFB3";
        ram_buffer(21493) := X"AEE40048";
        ram_buffer(21494) := X"8EE50048";
        ram_buffer(21495) := X"0C02502F";
        ram_buffer(21496) := X"02E02021";
        ram_buffer(21497) := X"8EE40010";
        ram_buffer(21498) := X"1000FF6D";
        ram_buffer(21499) := X"00000000";
        ram_buffer(21500) := X"8C820014";
        ram_buffer(21501) := X"27BDFEA0";
        ram_buffer(21502) := X"00801821";
        ram_buffer(21503) := X"8C460000";
        ram_buffer(21504) := X"AFB70154";
        ram_buffer(21505) := X"AFA40160";
        ram_buffer(21506) := X"8C970164";
        ram_buffer(21507) := X"8C440004";
        ram_buffer(21508) := X"8C6200C0";
        ram_buffer(21509) := X"8C630138";
        ram_buffer(21510) := X"AFB1013C";
        ram_buffer(21511) := X"AFA30134";
        ram_buffer(21512) := X"8FA30160";
        ram_buffer(21513) := X"AFB00138";
        ram_buffer(21514) := X"AFBF015C";
        ram_buffer(21515) := X"AFBE0158";
        ram_buffer(21516) := X"AFB60150";
        ram_buffer(21517) := X"AFB5014C";
        ram_buffer(21518) := X"AFB40148";
        ram_buffer(21519) := X"AFB30144";
        ram_buffer(21520) := X"AFB20140";
        ram_buffer(21521) := X"8C700140";
        ram_buffer(21522) := X"00A08821";
        ram_buffer(21523) := X"AEE60010";
        ram_buffer(21524) := X"10400005";
        ram_buffer(21525) := X"AEE40014";
        ram_buffer(21526) := X"8EE20044";
        ram_buffer(21527) := X"00000000";
        ram_buffer(21528) := X"104004C3";
        ram_buffer(21529) := X"00000000";
        ram_buffer(21530) := X"8FA20160";
        ram_buffer(21531) := X"8E230000";
        ram_buffer(21532) := X"8C420134";
        ram_buffer(21533) := X"8FA70134";
        ram_buffer(21534) := X"AFA20124";
        ram_buffer(21535) := X"AFA30130";
        ram_buffer(21536) := X"00401821";
        ram_buffer(21537) := X"00E2102A";
        ram_buffer(21538) := X"14400099";
        ram_buffer(21539) := X"3C04100D";
        ram_buffer(21540) := X"00031080";
        ram_buffer(21541) := X"24848968";
        ram_buffer(21542) := X"00822021";
        ram_buffer(21543) := X"00802821";
        ram_buffer(21544) := X"AFA40128";
        ram_buffer(21545) := X"27A40010";
        ram_buffer(21546) := X"00821021";
        ram_buffer(21547) := X"24E90001";
        ram_buffer(21548) := X"AFA2011C";
        ram_buffer(21549) := X"00403021";
        ram_buffer(21550) := X"00602021";
        ram_buffer(21551) := X"00003821";
        ram_buffer(21552) := X"10000006";
        ram_buffer(21553) := X"24080001";
        ram_buffer(21554) := X"24840001";
        ram_buffer(21555) := X"8FA70120";
        ram_buffer(21556) := X"24A50004";
        ram_buffer(21557) := X"10890012";
        ram_buffer(21558) := X"24C60004";
        ram_buffer(21559) := X"8CA20000";
        ram_buffer(21560) := X"8FA30130";
        ram_buffer(21561) := X"00021040";
        ram_buffer(21562) := X"00621021";
        ram_buffer(21563) := X"84420000";
        ram_buffer(21564) := X"00000000";
        ram_buffer(21565) := X"04400052";
        ram_buffer(21566) := X"AFA70120";
        ram_buffer(21567) := X"02021007";
        ram_buffer(21568) := X"1448FFF1";
        ram_buffer(21569) := X"ACC20000";
        ram_buffer(21570) := X"AFA40120";
        ram_buffer(21571) := X"24840001";
        ram_buffer(21572) := X"8FA70120";
        ram_buffer(21573) := X"24A50004";
        ram_buffer(21574) := X"1489FFF0";
        ram_buffer(21575) := X"24C60004";
        ram_buffer(21576) := X"8EF30040";
        ram_buffer(21577) := X"8EE2003C";
        ram_buffer(21578) := X"AFA00110";
        ram_buffer(21579) := X"02629821";
        ram_buffer(21580) := X"AFA00114";
        ram_buffer(21581) := X"241000FF";
        ram_buffer(21582) := X"8FA2011C";
        ram_buffer(21583) := X"00000000";
        ram_buffer(21584) := X"8C420000";
        ram_buffer(21585) := X"00000000";
        ram_buffer(21586) := X"10400223";
        ram_buffer(21587) := X"AFA2012C";
        ram_buffer(21588) := X"8FA20114";
        ram_buffer(21589) := X"00000000";
        ram_buffer(21590) := X"28420010";
        ram_buffer(21591) := X"14400275";
        ram_buffer(21592) := X"00000000";
        ram_buffer(21593) := X"8FA20120";
        ram_buffer(21594) := X"8FA30124";
        ram_buffer(21595) := X"00000000";
        ram_buffer(21596) := X"0043102A";
        ram_buffer(21597) := X"1440026F";
        ram_buffer(21598) := X"00000000";
        ram_buffer(21599) := X"8FA20114";
        ram_buffer(21600) := X"8EFE000C";
        ram_buffer(21601) := X"2454FFF0";
        ram_buffer(21602) := X"8EE20038";
        ram_buffer(21603) := X"00000000";
        ram_buffer(21604) := X"10400018";
        ram_buffer(21605) := X"00021043";
        ram_buffer(21606) := X"10400230";
        ram_buffer(21607) := X"00000000";
        ram_buffer(21608) := X"00009021";
        ram_buffer(21609) := X"00021043";
        ram_buffer(21610) := X"1440FFFE";
        ram_buffer(21611) := X"26520001";
        ram_buffer(21612) := X"00122100";
        ram_buffer(21613) := X"8EE20034";
        ram_buffer(21614) := X"13C00142";
        ram_buffer(21615) := X"00042880";
        ram_buffer(21616) := X"24420016";
        ram_buffer(21617) := X"00021080";
        ram_buffer(21618) := X"02E21021";
        ram_buffer(21619) := X"8C420004";
        ram_buffer(21620) := X"00042080";
        ram_buffer(21621) := X"00442021";
        ram_buffer(21622) := X"8C820000";
        ram_buffer(21623) := X"00000000";
        ram_buffer(21624) := X"24420001";
        ram_buffer(21625) := X"AC820000";
        ram_buffer(21626) := X"0C024B01";
        ram_buffer(21627) := X"02E02021";
        ram_buffer(21628) := X"8EFE000C";
        ram_buffer(21629) := X"8EE20034";
        ram_buffer(21630) := X"13C0005E";
        ram_buffer(21631) := X"00000000";
        ram_buffer(21632) := X"24420016";
        ram_buffer(21633) := X"00021080";
        ram_buffer(21634) := X"02E21021";
        ram_buffer(21635) := X"8C440004";
        ram_buffer(21636) := X"00000000";
        ram_buffer(21637) := X"8C8203C0";
        ram_buffer(21638) := X"00000000";
        ram_buffer(21639) := X"24420001";
        ram_buffer(21640) := X"AC8203C0";
        ram_buffer(21641) := X"2A820010";
        ram_buffer(21642) := X"AFB40114";
        ram_buffer(21643) := X"8EF30040";
        ram_buffer(21644) := X"14400005";
        ram_buffer(21645) := X"2694FFF0";
        ram_buffer(21646) := X"1000FFD3";
        ram_buffer(21647) := X"AFA00110";
        ram_buffer(21648) := X"1000FFAE";
        ram_buffer(21649) := X"00021023";
        ram_buffer(21650) := X"0000F021";
        ram_buffer(21651) := X"8FA3012C";
        ram_buffer(21652) := X"00000000";
        ram_buffer(21653) := X"28620002";
        ram_buffer(21654) := X"14400207";
        ram_buffer(21655) := X"30640001";
        ram_buffer(21656) := X"027E1021";
        ram_buffer(21657) := X"27C30001";
        ram_buffer(21658) := X"AFA30110";
        ram_buffer(21659) := X"A0440000";
        ram_buffer(21660) := X"8FA20124";
        ram_buffer(21661) := X"8FA30134";
        ram_buffer(21662) := X"24420001";
        ram_buffer(21663) := X"AFA20124";
        ram_buffer(21664) := X"0062102A";
        ram_buffer(21665) := X"8FA3011C";
        ram_buffer(21666) := X"00000000";
        ram_buffer(21667) := X"24630004";
        ram_buffer(21668) := X"AFA3011C";
        ram_buffer(21669) := X"8FA30128";
        ram_buffer(21670) := X"00000000";
        ram_buffer(21671) := X"24630004";
        ram_buffer(21672) := X"1040FFA5";
        ram_buffer(21673) := X"AFA30128";
        ram_buffer(21674) := X"8FA20114";
        ram_buffer(21675) := X"00000000";
        ram_buffer(21676) := X"10400457";
        ram_buffer(21677) := X"00000000";
        ram_buffer(21678) := X"8EE2003C";
        ram_buffer(21679) := X"8EE40038";
        ram_buffer(21680) := X"8FA30110";
        ram_buffer(21681) := X"24840001";
        ram_buffer(21682) := X"0062F021";
        ram_buffer(21683) := X"24027FFF";
        ram_buffer(21684) := X"AEE40038";
        ram_buffer(21685) := X"10820004";
        ram_buffer(21686) := X"AEFE003C";
        ram_buffer(21687) := X"2FDE03AA";
        ram_buffer(21688) := X"17C00003";
        ram_buffer(21689) := X"00000000";
        ram_buffer(21690) := X"0C024CF4";
        ram_buffer(21691) := X"02E02021";
        ram_buffer(21692) := X"8FA20160";
        ram_buffer(21693) := X"8FA30160";
        ram_buffer(21694) := X"8C420014";
        ram_buffer(21695) := X"8EE60010";
        ram_buffer(21696) := X"8EE40014";
        ram_buffer(21697) := X"8C6500C0";
        ram_buffer(21698) := X"AC460000";
        ram_buffer(21699) := X"10A0000C";
        ram_buffer(21700) := X"AC440004";
        ram_buffer(21701) := X"8EE20044";
        ram_buffer(21702) := X"00000000";
        ram_buffer(21703) := X"14400007";
        ram_buffer(21704) := X"2442FFFF";
        ram_buffer(21705) := X"8EE40048";
        ram_buffer(21706) := X"00A01021";
        ram_buffer(21707) := X"24840001";
        ram_buffer(21708) := X"30840007";
        ram_buffer(21709) := X"AEE40048";
        ram_buffer(21710) := X"2442FFFF";
        ram_buffer(21711) := X"AEE20044";
        ram_buffer(21712) := X"8FBF015C";
        ram_buffer(21713) := X"8FBE0158";
        ram_buffer(21714) := X"8FB70154";
        ram_buffer(21715) := X"8FB60150";
        ram_buffer(21716) := X"8FB5014C";
        ram_buffer(21717) := X"8FB40148";
        ram_buffer(21718) := X"8FB30144";
        ram_buffer(21719) := X"8FB20140";
        ram_buffer(21720) := X"8FB1013C";
        ram_buffer(21721) := X"8FB00138";
        ram_buffer(21722) := X"24020001";
        ram_buffer(21723) := X"03E00008";
        ram_buffer(21724) := X"27BD0160";
        ram_buffer(21725) := X"24420012";
        ram_buffer(21726) := X"00021080";
        ram_buffer(21727) := X"02E21021";
        ram_buffer(21728) := X"8C420004";
        ram_buffer(21729) := X"8EF2001C";
        ram_buffer(21730) := X"805104F0";
        ram_buffer(21731) := X"8C5603C0";
        ram_buffer(21732) := X"12200196";
        ram_buffer(21733) := X"24030027";
        ram_buffer(21734) := X"24020001";
        ram_buffer(21735) := X"02221004";
        ram_buffer(21736) := X"02321821";
        ram_buffer(21737) := X"24040018";
        ram_buffer(21738) := X"2442FFFF";
        ram_buffer(21739) := X"00561024";
        ram_buffer(21740) := X"8EE60018";
        ram_buffer(21741) := X"0083B023";
        ram_buffer(21742) := X"02C21004";
        ram_buffer(21743) := X"28640008";
        ram_buffer(21744) := X"AFA30118";
        ram_buffer(21745) := X"148001A8";
        ram_buffer(21746) := X"0046B025";
        ram_buffer(21747) := X"00609021";
        ram_buffer(21748) := X"8EE40010";
        ram_buffer(21749) := X"00161403";
        ram_buffer(21750) := X"24870001";
        ram_buffer(21751) := X"AEE70010";
        ram_buffer(21752) := X"A0820000";
        ram_buffer(21753) := X"8EE40014";
        ram_buffer(21754) := X"2652FFF8";
        ram_buffer(21755) := X"2484FFFF";
        ram_buffer(21756) := X"AEE40014";
        ram_buffer(21757) := X"1080003C";
        ram_buffer(21758) := X"305100FF";
        ram_buffer(21759) := X"12300051";
        ram_buffer(21760) := X"00000000";
        ram_buffer(21761) := X"2A420008";
        ram_buffer(21762) := X"1040FFF1";
        ram_buffer(21763) := X"0016B200";
        ram_buffer(21764) := X"8FA30118";
        ram_buffer(21765) := X"8EE2000C";
        ram_buffer(21766) := X"30630007";
        ram_buffer(21767) := X"AFA30118";
        ram_buffer(21768) := X"AEF60018";
        ram_buffer(21769) := X"AEE3001C";
        ram_buffer(21770) := X"1440009F";
        ram_buffer(21771) := X"AFB40114";
        ram_buffer(21772) := X"8FA20110";
        ram_buffer(21773) := X"00000000";
        ram_buffer(21774) := X"1040009B";
        ram_buffer(21775) := X"02621021";
        ram_buffer(21776) := X"8FB20118";
        ram_buffer(21777) := X"26710001";
        ram_buffer(21778) := X"AFA20110";
        ram_buffer(21779) := X"17C0001F";
        ram_buffer(21780) := X"26560001";
        ram_buffer(21781) := X"9222FFFF";
        ram_buffer(21782) := X"24030018";
        ram_buffer(21783) := X"30420001";
        ram_buffer(21784) := X"00762823";
        ram_buffer(21785) := X"8EE70018";
        ram_buffer(21786) := X"00A21004";
        ram_buffer(21787) := X"2AC40008";
        ram_buffer(21788) := X"14800013";
        ram_buffer(21789) := X"00479825";
        ram_buffer(21790) := X"8EE40010";
        ram_buffer(21791) := X"00131403";
        ram_buffer(21792) := X"24870001";
        ram_buffer(21793) := X"AEE70010";
        ram_buffer(21794) := X"A0820000";
        ram_buffer(21795) := X"8EE40014";
        ram_buffer(21796) := X"26D6FFF8";
        ram_buffer(21797) := X"2484FFFF";
        ram_buffer(21798) := X"AEE40014";
        ram_buffer(21799) := X"1080004A";
        ram_buffer(21800) := X"305E00FF";
        ram_buffer(21801) := X"13D0005F";
        ram_buffer(21802) := X"00000000";
        ram_buffer(21803) := X"2AC20008";
        ram_buffer(21804) := X"1040FFF1";
        ram_buffer(21805) := X"00139A00";
        ram_buffer(21806) := X"2652FFF9";
        ram_buffer(21807) := X"32560007";
        ram_buffer(21808) := X"AEF30018";
        ram_buffer(21809) := X"AEF6001C";
        ram_buffer(21810) := X"02C09021";
        ram_buffer(21811) := X"8FA20110";
        ram_buffer(21812) := X"00000000";
        ram_buffer(21813) := X"10510074";
        ram_buffer(21814) := X"26310001";
        ram_buffer(21815) := X"8EFE000C";
        ram_buffer(21816) := X"1000FFDA";
        ram_buffer(21817) := X"00000000";
        ram_buffer(21818) := X"8EE40020";
        ram_buffer(21819) := X"00000000";
        ram_buffer(21820) := X"8C950014";
        ram_buffer(21821) := X"00000000";
        ram_buffer(21822) := X"8EA2000C";
        ram_buffer(21823) := X"00000000";
        ram_buffer(21824) := X"0040F809";
        ram_buffer(21825) := X"00000000";
        ram_buffer(21826) := X"14400009";
        ram_buffer(21827) := X"24030016";
        ram_buffer(21828) := X"8EE40020";
        ram_buffer(21829) := X"00000000";
        ram_buffer(21830) := X"8C820000";
        ram_buffer(21831) := X"00000000";
        ram_buffer(21832) := X"8C480000";
        ram_buffer(21833) := X"00000000";
        ram_buffer(21834) := X"0100F809";
        ram_buffer(21835) := X"AC430014";
        ram_buffer(21836) := X"8EA40000";
        ram_buffer(21837) := X"8EA20004";
        ram_buffer(21838) := X"AEE40010";
        ram_buffer(21839) := X"1630FFB1";
        ram_buffer(21840) := X"AEE20014";
        ram_buffer(21841) := X"8EE20010";
        ram_buffer(21842) := X"00000000";
        ram_buffer(21843) := X"24440001";
        ram_buffer(21844) := X"AEE40010";
        ram_buffer(21845) := X"A0400000";
        ram_buffer(21846) := X"8EE20014";
        ram_buffer(21847) := X"00000000";
        ram_buffer(21848) := X"2442FFFF";
        ram_buffer(21849) := X"1440FFA7";
        ram_buffer(21850) := X"AEE20014";
        ram_buffer(21851) := X"8EE40020";
        ram_buffer(21852) := X"00000000";
        ram_buffer(21853) := X"8C910014";
        ram_buffer(21854) := X"00000000";
        ram_buffer(21855) := X"8E22000C";
        ram_buffer(21856) := X"00000000";
        ram_buffer(21857) := X"0040F809";
        ram_buffer(21858) := X"00000000";
        ram_buffer(21859) := X"14400009";
        ram_buffer(21860) := X"24030016";
        ram_buffer(21861) := X"8EE40020";
        ram_buffer(21862) := X"00000000";
        ram_buffer(21863) := X"8C820000";
        ram_buffer(21864) := X"00000000";
        ram_buffer(21865) := X"8C470000";
        ram_buffer(21866) := X"00000000";
        ram_buffer(21867) := X"00E0F809";
        ram_buffer(21868) := X"AC430014";
        ram_buffer(21869) := X"8E240000";
        ram_buffer(21870) := X"8E220004";
        ram_buffer(21871) := X"AEE40010";
        ram_buffer(21872) := X"1000FF90";
        ram_buffer(21873) := X"AEE20014";
        ram_buffer(21874) := X"8EE40020";
        ram_buffer(21875) := X"00000000";
        ram_buffer(21876) := X"8C950014";
        ram_buffer(21877) := X"00000000";
        ram_buffer(21878) := X"8EA2000C";
        ram_buffer(21879) := X"00000000";
        ram_buffer(21880) := X"0040F809";
        ram_buffer(21881) := X"00000000";
        ram_buffer(21882) := X"14400009";
        ram_buffer(21883) := X"24030016";
        ram_buffer(21884) := X"8EE40020";
        ram_buffer(21885) := X"00000000";
        ram_buffer(21886) := X"8C820000";
        ram_buffer(21887) := X"00000000";
        ram_buffer(21888) := X"8C480000";
        ram_buffer(21889) := X"00000000";
        ram_buffer(21890) := X"0100F809";
        ram_buffer(21891) := X"AC430014";
        ram_buffer(21892) := X"8EA40000";
        ram_buffer(21893) := X"8EA20004";
        ram_buffer(21894) := X"AEE40010";
        ram_buffer(21895) := X"17D0FFA3";
        ram_buffer(21896) := X"AEE20014";
        ram_buffer(21897) := X"8EE20010";
        ram_buffer(21898) := X"00000000";
        ram_buffer(21899) := X"24440001";
        ram_buffer(21900) := X"AEE40010";
        ram_buffer(21901) := X"A0400000";
        ram_buffer(21902) := X"8EE20014";
        ram_buffer(21903) := X"00000000";
        ram_buffer(21904) := X"2442FFFF";
        ram_buffer(21905) := X"1440FF99";
        ram_buffer(21906) := X"AEE20014";
        ram_buffer(21907) := X"8EE40020";
        ram_buffer(21908) := X"00000000";
        ram_buffer(21909) := X"8C9E0014";
        ram_buffer(21910) := X"00000000";
        ram_buffer(21911) := X"8FC2000C";
        ram_buffer(21912) := X"00000000";
        ram_buffer(21913) := X"0040F809";
        ram_buffer(21914) := X"00000000";
        ram_buffer(21915) := X"14400009";
        ram_buffer(21916) := X"24030016";
        ram_buffer(21917) := X"8EE40020";
        ram_buffer(21918) := X"00000000";
        ram_buffer(21919) := X"8C820000";
        ram_buffer(21920) := X"00000000";
        ram_buffer(21921) := X"8C470000";
        ram_buffer(21922) := X"00000000";
        ram_buffer(21923) := X"00E0F809";
        ram_buffer(21924) := X"AC430014";
        ram_buffer(21925) := X"8FC40000";
        ram_buffer(21926) := X"8FC20004";
        ram_buffer(21927) := X"AEE40010";
        ram_buffer(21928) := X"1000FF82";
        ram_buffer(21929) := X"AEE20014";
        ram_buffer(21930) := X"2A820010";
        ram_buffer(21931) := X"8EF30040";
        ram_buffer(21932) := X"1440FEE5";
        ram_buffer(21933) := X"2694FFF0";
        ram_buffer(21934) := X"8EFE000C";
        ram_buffer(21935) := X"1000FEB2";
        ram_buffer(21936) := X"AFA00110";
        ram_buffer(21937) := X"24420012";
        ram_buffer(21938) := X"00021080";
        ram_buffer(21939) := X"02E21021";
        ram_buffer(21940) := X"8C420004";
        ram_buffer(21941) := X"00000000";
        ram_buffer(21942) := X"00442021";
        ram_buffer(21943) := X"80910400";
        ram_buffer(21944) := X"00451021";
        ram_buffer(21945) := X"8C560000";
        ram_buffer(21946) := X"8EFE001C";
        ram_buffer(21947) := X"122000CD";
        ram_buffer(21948) := X"24020001";
        ram_buffer(21949) := X"02221004";
        ram_buffer(21950) := X"023E1821";
        ram_buffer(21951) := X"2442FFFF";
        ram_buffer(21952) := X"24040018";
        ram_buffer(21953) := X"00832023";
        ram_buffer(21954) := X"00561024";
        ram_buffer(21955) := X"8EE50018";
        ram_buffer(21956) := X"00821004";
        ram_buffer(21957) := X"28640008";
        ram_buffer(21958) := X"0045F025";
        ram_buffer(21959) := X"AFA30114";
        ram_buffer(21960) := X"00608821";
        ram_buffer(21961) := X"14800015";
        ram_buffer(21962) := X"00601021";
        ram_buffer(21963) := X"8EE40010";
        ram_buffer(21964) := X"001E1403";
        ram_buffer(21965) := X"24870001";
        ram_buffer(21966) := X"AEE70010";
        ram_buffer(21967) := X"A0820000";
        ram_buffer(21968) := X"8EE40014";
        ram_buffer(21969) := X"2631FFF8";
        ram_buffer(21970) := X"2484FFFF";
        ram_buffer(21971) := X"AEE40014";
        ram_buffer(21972) := X"10800031";
        ram_buffer(21973) := X"305600FF";
        ram_buffer(21974) := X"12D00046";
        ram_buffer(21975) := X"00000000";
        ram_buffer(21976) := X"2A220008";
        ram_buffer(21977) := X"1040FFF1";
        ram_buffer(21978) := X"001EF200";
        ram_buffer(21979) := X"8FA20114";
        ram_buffer(21980) := X"00000000";
        ram_buffer(21981) := X"30420007";
        ram_buffer(21982) := X"AFA20114";
        ram_buffer(21983) := X"AEFE0018";
        ram_buffer(21984) := X"1240FE99";
        ram_buffer(21985) := X"AEE2001C";
        ram_buffer(21986) := X"8EE4000C";
        ram_buffer(21987) := X"8EF60038";
        ram_buffer(21988) := X"1480FE95";
        ram_buffer(21989) := X"00401821";
        ram_buffer(21990) := X"24020001";
        ram_buffer(21991) := X"02421004";
        ram_buffer(21992) := X"00728821";
        ram_buffer(21993) := X"2442FFFF";
        ram_buffer(21994) := X"24030018";
        ram_buffer(21995) := X"00561024";
        ram_buffer(21996) := X"0071B023";
        ram_buffer(21997) := X"02C2B004";
        ram_buffer(21998) := X"2A220008";
        ram_buffer(21999) := X"14400013";
        ram_buffer(22000) := X"02DEB025";
        ram_buffer(22001) := X"0220F021";
        ram_buffer(22002) := X"8EE40010";
        ram_buffer(22003) := X"00161403";
        ram_buffer(22004) := X"24860001";
        ram_buffer(22005) := X"AEE60010";
        ram_buffer(22006) := X"A0820000";
        ram_buffer(22007) := X"8EE40014";
        ram_buffer(22008) := X"27DEFFF8";
        ram_buffer(22009) := X"2484FFFF";
        ram_buffer(22010) := X"AEE40014";
        ram_buffer(22011) := X"10800042";
        ram_buffer(22012) := X"305200FF";
        ram_buffer(22013) := X"12500057";
        ram_buffer(22014) := X"00000000";
        ram_buffer(22015) := X"2BC20008";
        ram_buffer(22016) := X"1040FFF1";
        ram_buffer(22017) := X"0016B200";
        ram_buffer(22018) := X"32310007";
        ram_buffer(22019) := X"AEF60018";
        ram_buffer(22020) := X"1000FE75";
        ram_buffer(22021) := X"AEF1001C";
        ram_buffer(22022) := X"8EE40020";
        ram_buffer(22023) := X"00000000";
        ram_buffer(22024) := X"8C950014";
        ram_buffer(22025) := X"00000000";
        ram_buffer(22026) := X"8EA2000C";
        ram_buffer(22027) := X"00000000";
        ram_buffer(22028) := X"0040F809";
        ram_buffer(22029) := X"00000000";
        ram_buffer(22030) := X"14400009";
        ram_buffer(22031) := X"24030016";
        ram_buffer(22032) := X"8EE40020";
        ram_buffer(22033) := X"00000000";
        ram_buffer(22034) := X"8C820000";
        ram_buffer(22035) := X"00000000";
        ram_buffer(22036) := X"8C480000";
        ram_buffer(22037) := X"00000000";
        ram_buffer(22038) := X"0100F809";
        ram_buffer(22039) := X"AC430014";
        ram_buffer(22040) := X"8EA40000";
        ram_buffer(22041) := X"8EA20004";
        ram_buffer(22042) := X"AEE40010";
        ram_buffer(22043) := X"16D0FFBC";
        ram_buffer(22044) := X"AEE20014";
        ram_buffer(22045) := X"8EE20010";
        ram_buffer(22046) := X"00000000";
        ram_buffer(22047) := X"24440001";
        ram_buffer(22048) := X"AEE40010";
        ram_buffer(22049) := X"A0400000";
        ram_buffer(22050) := X"8EE20014";
        ram_buffer(22051) := X"00000000";
        ram_buffer(22052) := X"2442FFFF";
        ram_buffer(22053) := X"1440FFB2";
        ram_buffer(22054) := X"AEE20014";
        ram_buffer(22055) := X"8EE40020";
        ram_buffer(22056) := X"00000000";
        ram_buffer(22057) := X"8C960014";
        ram_buffer(22058) := X"00000000";
        ram_buffer(22059) := X"8EC2000C";
        ram_buffer(22060) := X"00000000";
        ram_buffer(22061) := X"0040F809";
        ram_buffer(22062) := X"00000000";
        ram_buffer(22063) := X"14400009";
        ram_buffer(22064) := X"00000000";
        ram_buffer(22065) := X"8EE40020";
        ram_buffer(22066) := X"24030016";
        ram_buffer(22067) := X"8C820000";
        ram_buffer(22068) := X"00000000";
        ram_buffer(22069) := X"8C470000";
        ram_buffer(22070) := X"00000000";
        ram_buffer(22071) := X"00E0F809";
        ram_buffer(22072) := X"AC430014";
        ram_buffer(22073) := X"8EC40000";
        ram_buffer(22074) := X"8EC20004";
        ram_buffer(22075) := X"AEE40010";
        ram_buffer(22076) := X"1000FF9B";
        ram_buffer(22077) := X"AEE20014";
        ram_buffer(22078) := X"8EE40020";
        ram_buffer(22079) := X"00000000";
        ram_buffer(22080) := X"8C950014";
        ram_buffer(22081) := X"00000000";
        ram_buffer(22082) := X"8EA2000C";
        ram_buffer(22083) := X"00000000";
        ram_buffer(22084) := X"0040F809";
        ram_buffer(22085) := X"00000000";
        ram_buffer(22086) := X"14400009";
        ram_buffer(22087) := X"24030016";
        ram_buffer(22088) := X"8EE40020";
        ram_buffer(22089) := X"00000000";
        ram_buffer(22090) := X"8C820000";
        ram_buffer(22091) := X"00000000";
        ram_buffer(22092) := X"8C470000";
        ram_buffer(22093) := X"00000000";
        ram_buffer(22094) := X"00E0F809";
        ram_buffer(22095) := X"AC430014";
        ram_buffer(22096) := X"8EA40000";
        ram_buffer(22097) := X"8EA20004";
        ram_buffer(22098) := X"AEE40010";
        ram_buffer(22099) := X"1650FFAB";
        ram_buffer(22100) := X"AEE20014";
        ram_buffer(22101) := X"8EE20010";
        ram_buffer(22102) := X"00000000";
        ram_buffer(22103) := X"24440001";
        ram_buffer(22104) := X"AEE40010";
        ram_buffer(22105) := X"A0400000";
        ram_buffer(22106) := X"8EE20014";
        ram_buffer(22107) := X"00000000";
        ram_buffer(22108) := X"2442FFFF";
        ram_buffer(22109) := X"1440FFA1";
        ram_buffer(22110) := X"AEE20014";
        ram_buffer(22111) := X"8EE40020";
        ram_buffer(22112) := X"00000000";
        ram_buffer(22113) := X"8C920014";
        ram_buffer(22114) := X"00000000";
        ram_buffer(22115) := X"8E42000C";
        ram_buffer(22116) := X"00000000";
        ram_buffer(22117) := X"0040F809";
        ram_buffer(22118) := X"00000000";
        ram_buffer(22119) := X"14400009";
        ram_buffer(22120) := X"24030016";
        ram_buffer(22121) := X"8EE40020";
        ram_buffer(22122) := X"00000000";
        ram_buffer(22123) := X"8C820000";
        ram_buffer(22124) := X"00000000";
        ram_buffer(22125) := X"8C460000";
        ram_buffer(22126) := X"00000000";
        ram_buffer(22127) := X"00C0F809";
        ram_buffer(22128) := X"AC430014";
        ram_buffer(22129) := X"8E440000";
        ram_buffer(22130) := X"8E420004";
        ram_buffer(22131) := X"AEE40010";
        ram_buffer(22132) := X"1000FF8A";
        ram_buffer(22133) := X"AEE20014";
        ram_buffer(22134) := X"8FA20114";
        ram_buffer(22135) := X"00000000";
        ram_buffer(22136) := X"24420001";
        ram_buffer(22137) := X"1000FE22";
        ram_buffer(22138) := X"AFA20114";
        ram_buffer(22139) := X"8EE40020";
        ram_buffer(22140) := X"00000000";
        ram_buffer(22141) := X"8C820000";
        ram_buffer(22142) := X"00000000";
        ram_buffer(22143) := X"8C460000";
        ram_buffer(22144) := X"00000000";
        ram_buffer(22145) := X"00C0F809";
        ram_buffer(22146) := X"AC430014";
        ram_buffer(22147) := X"8EE2000C";
        ram_buffer(22148) := X"00000000";
        ram_buffer(22149) := X"1040FE60";
        ram_buffer(22150) := X"00000000";
        ram_buffer(22151) := X"1000FE01";
        ram_buffer(22152) := X"0040F021";
        ram_buffer(22153) := X"8EE40020";
        ram_buffer(22154) := X"24030027";
        ram_buffer(22155) := X"8C820000";
        ram_buffer(22156) := X"00000000";
        ram_buffer(22157) := X"8C460000";
        ram_buffer(22158) := X"00000000";
        ram_buffer(22159) := X"00C0F809";
        ram_buffer(22160) := X"AC430014";
        ram_buffer(22161) := X"8EE2000C";
        ram_buffer(22162) := X"00000000";
        ram_buffer(22163) := X"1440FDE6";
        ram_buffer(22164) := X"24020001";
        ram_buffer(22165) := X"1000FF28";
        ram_buffer(22166) := X"02221004";
        ram_buffer(22167) := X"00002021";
        ram_buffer(22168) := X"1000FDD4";
        ram_buffer(22169) := X"00009021";
        ram_buffer(22170) := X"AEF60018";
        ram_buffer(22171) := X"AEE3001C";
        ram_buffer(22172) := X"1000FE6F";
        ram_buffer(22173) := X"AFB40114";
        ram_buffer(22174) := X"8EE20038";
        ram_buffer(22175) := X"00000000";
        ram_buffer(22176) := X"10400018";
        ram_buffer(22177) := X"00021043";
        ram_buffer(22178) := X"1040025F";
        ram_buffer(22179) := X"00002021";
        ram_buffer(22180) := X"0000A021";
        ram_buffer(22181) := X"00021043";
        ram_buffer(22182) := X"1440FFFE";
        ram_buffer(22183) := X"26940001";
        ram_buffer(22184) := X"00142100";
        ram_buffer(22185) := X"8EE6000C";
        ram_buffer(22186) := X"8EE20034";
        ram_buffer(22187) := X"10C00024";
        ram_buffer(22188) := X"00043080";
        ram_buffer(22189) := X"24420016";
        ram_buffer(22190) := X"00021080";
        ram_buffer(22191) := X"02E21021";
        ram_buffer(22192) := X"8C420004";
        ram_buffer(22193) := X"00042080";
        ram_buffer(22194) := X"00442021";
        ram_buffer(22195) := X"8C820000";
        ram_buffer(22196) := X"00000000";
        ram_buffer(22197) := X"24420001";
        ram_buffer(22198) := X"AC820000";
        ram_buffer(22199) := X"0C024B01";
        ram_buffer(22200) := X"02E02021";
        ram_buffer(22201) := X"8FA20114";
        ram_buffer(22202) := X"8EF4000C";
        ram_buffer(22203) := X"00022100";
        ram_buffer(22204) := X"8EE20034";
        ram_buffer(22205) := X"12800095";
        ram_buffer(22206) := X"24840001";
        ram_buffer(22207) := X"24420016";
        ram_buffer(22208) := X"00021080";
        ram_buffer(22209) := X"02E21021";
        ram_buffer(22210) := X"8C420004";
        ram_buffer(22211) := X"00042080";
        ram_buffer(22212) := X"00442021";
        ram_buffer(22213) := X"8C820000";
        ram_buffer(22214) := X"00000000";
        ram_buffer(22215) := X"24420001";
        ram_buffer(22216) := X"AC820000";
        ram_buffer(22217) := X"8EF30040";
        ram_buffer(22218) := X"AFA00110";
        ram_buffer(22219) := X"1000FDD0";
        ram_buffer(22220) := X"AFA00114";
        ram_buffer(22221) := X"8FBE0110";
        ram_buffer(22222) := X"1000FDC4";
        ram_buffer(22223) := X"00000000";
        ram_buffer(22224) := X"24420012";
        ram_buffer(22225) := X"00021080";
        ram_buffer(22226) := X"02E21021";
        ram_buffer(22227) := X"8C420004";
        ram_buffer(22228) := X"00000000";
        ram_buffer(22229) := X"00442021";
        ram_buffer(22230) := X"80910400";
        ram_buffer(22231) := X"00461021";
        ram_buffer(22232) := X"8C520000";
        ram_buffer(22233) := X"8EF5001C";
        ram_buffer(22234) := X"122001BF";
        ram_buffer(22235) := X"24020001";
        ram_buffer(22236) := X"02221004";
        ram_buffer(22237) := X"02353021";
        ram_buffer(22238) := X"2442FFFF";
        ram_buffer(22239) := X"24030018";
        ram_buffer(22240) := X"00521024";
        ram_buffer(22241) := X"8EE70018";
        ram_buffer(22242) := X"00669023";
        ram_buffer(22243) := X"02421004";
        ram_buffer(22244) := X"28C40008";
        ram_buffer(22245) := X"00479025";
        ram_buffer(22246) := X"14800012";
        ram_buffer(22247) := X"00C0B021";
        ram_buffer(22248) := X"8EE20010";
        ram_buffer(22249) := X"00128C03";
        ram_buffer(22250) := X"24440001";
        ram_buffer(22251) := X"AEE40010";
        ram_buffer(22252) := X"A0510000";
        ram_buffer(22253) := X"8EE20014";
        ram_buffer(22254) := X"26D6FFF8";
        ram_buffer(22255) := X"2442FFFF";
        ram_buffer(22256) := X"AEE20014";
        ram_buffer(22257) := X"1040002E";
        ram_buffer(22258) := X"323500FF";
        ram_buffer(22259) := X"12B00045";
        ram_buffer(22260) := X"00000000";
        ram_buffer(22261) := X"2AC20008";
        ram_buffer(22262) := X"1040FFF1";
        ram_buffer(22263) := X"00129200";
        ram_buffer(22264) := X"30C60007";
        ram_buffer(22265) := X"AEF20018";
        ram_buffer(22266) := X"1280FFBC";
        ram_buffer(22267) := X"AEE6001C";
        ram_buffer(22268) := X"8EE4000C";
        ram_buffer(22269) := X"8EE70038";
        ram_buffer(22270) := X"1480FFB8";
        ram_buffer(22271) := X"24020001";
        ram_buffer(22272) := X"02821004";
        ram_buffer(22273) := X"00D48821";
        ram_buffer(22274) := X"2442FFFF";
        ram_buffer(22275) := X"24030018";
        ram_buffer(22276) := X"00712023";
        ram_buffer(22277) := X"00471024";
        ram_buffer(22278) := X"00821004";
        ram_buffer(22279) := X"2A240008";
        ram_buffer(22280) := X"14800014";
        ram_buffer(22281) := X"00529025";
        ram_buffer(22282) := X"0220A021";
        ram_buffer(22283) := X"8EE20010";
        ram_buffer(22284) := X"00122403";
        ram_buffer(22285) := X"24450001";
        ram_buffer(22286) := X"AEE50010";
        ram_buffer(22287) := X"A0440000";
        ram_buffer(22288) := X"8EE20014";
        ram_buffer(22289) := X"308300FF";
        ram_buffer(22290) := X"2442FFFF";
        ram_buffer(22291) := X"2694FFF8";
        ram_buffer(22292) := X"AEE20014";
        ram_buffer(22293) := X"10400192";
        ram_buffer(22294) := X"0060A821";
        ram_buffer(22295) := X"12B001AA";
        ram_buffer(22296) := X"00000000";
        ram_buffer(22297) := X"2A820008";
        ram_buffer(22298) := X"1040FFF0";
        ram_buffer(22299) := X"00129200";
        ram_buffer(22300) := X"32310007";
        ram_buffer(22301) := X"AEF20018";
        ram_buffer(22302) := X"1000FF98";
        ram_buffer(22303) := X"AEF1001C";
        ram_buffer(22304) := X"8EE40020";
        ram_buffer(22305) := X"AFA60110";
        ram_buffer(22306) := X"8C910014";
        ram_buffer(22307) := X"00000000";
        ram_buffer(22308) := X"8E22000C";
        ram_buffer(22309) := X"00000000";
        ram_buffer(22310) := X"0040F809";
        ram_buffer(22311) := X"00000000";
        ram_buffer(22312) := X"8FA60110";
        ram_buffer(22313) := X"1440000A";
        ram_buffer(22314) := X"24030016";
        ram_buffer(22315) := X"8EE40020";
        ram_buffer(22316) := X"00000000";
        ram_buffer(22317) := X"8C820000";
        ram_buffer(22318) := X"00000000";
        ram_buffer(22319) := X"8C480000";
        ram_buffer(22320) := X"00000000";
        ram_buffer(22321) := X"0100F809";
        ram_buffer(22322) := X"AC430014";
        ram_buffer(22323) := X"8FA60110";
        ram_buffer(22324) := X"8E240000";
        ram_buffer(22325) := X"8E220004";
        ram_buffer(22326) := X"AEE40010";
        ram_buffer(22327) := X"16B0FFBD";
        ram_buffer(22328) := X"AEE20014";
        ram_buffer(22329) := X"8EE20010";
        ram_buffer(22330) := X"00000000";
        ram_buffer(22331) := X"24440001";
        ram_buffer(22332) := X"AEE40010";
        ram_buffer(22333) := X"A0400000";
        ram_buffer(22334) := X"8EE20014";
        ram_buffer(22335) := X"00000000";
        ram_buffer(22336) := X"2442FFFF";
        ram_buffer(22337) := X"1440FFB3";
        ram_buffer(22338) := X"AEE20014";
        ram_buffer(22339) := X"8EE40020";
        ram_buffer(22340) := X"AFA60110";
        ram_buffer(22341) := X"8C910014";
        ram_buffer(22342) := X"00000000";
        ram_buffer(22343) := X"8E22000C";
        ram_buffer(22344) := X"00000000";
        ram_buffer(22345) := X"0040F809";
        ram_buffer(22346) := X"00000000";
        ram_buffer(22347) := X"8FA60110";
        ram_buffer(22348) := X"104001AA";
        ram_buffer(22349) := X"24030016";
        ram_buffer(22350) := X"8E240000";
        ram_buffer(22351) := X"8E220004";
        ram_buffer(22352) := X"AEE40010";
        ram_buffer(22353) := X"1000FFA3";
        ram_buffer(22354) := X"AEE20014";
        ram_buffer(22355) := X"24420012";
        ram_buffer(22356) := X"00021080";
        ram_buffer(22357) := X"02E21021";
        ram_buffer(22358) := X"8C420004";
        ram_buffer(22359) := X"00042880";
        ram_buffer(22360) := X"00442021";
        ram_buffer(22361) := X"80910400";
        ram_buffer(22362) := X"00451021";
        ram_buffer(22363) := X"8C520000";
        ram_buffer(22364) := X"8EF6001C";
        ram_buffer(22365) := X"12200119";
        ram_buffer(22366) := X"24020001";
        ram_buffer(22367) := X"02221004";
        ram_buffer(22368) := X"2442FFFF";
        ram_buffer(22369) := X"02368821";
        ram_buffer(22370) := X"24030018";
        ram_buffer(22371) := X"00521024";
        ram_buffer(22372) := X"8EE50018";
        ram_buffer(22373) := X"00719023";
        ram_buffer(22374) := X"02421004";
        ram_buffer(22375) := X"2A240008";
        ram_buffer(22376) := X"14800125";
        ram_buffer(22377) := X"00459025";
        ram_buffer(22378) := X"0220B021";
        ram_buffer(22379) := X"8EE20010";
        ram_buffer(22380) := X"00122403";
        ram_buffer(22381) := X"24450001";
        ram_buffer(22382) := X"AEE50010";
        ram_buffer(22383) := X"A0440000";
        ram_buffer(22384) := X"8EE20014";
        ram_buffer(22385) := X"308300FF";
        ram_buffer(22386) := X"2442FFFF";
        ram_buffer(22387) := X"26D6FFF8";
        ram_buffer(22388) := X"AEE20014";
        ram_buffer(22389) := X"1040005A";
        ram_buffer(22390) := X"0060A821";
        ram_buffer(22391) := X"12B00072";
        ram_buffer(22392) := X"00000000";
        ram_buffer(22393) := X"2AC20008";
        ram_buffer(22394) := X"1040FFF0";
        ram_buffer(22395) := X"00129200";
        ram_buffer(22396) := X"32310007";
        ram_buffer(22397) := X"8FA20128";
        ram_buffer(22398) := X"AEF1001C";
        ram_buffer(22399) := X"8C420000";
        ram_buffer(22400) := X"8FA30130";
        ram_buffer(22401) := X"00021040";
        ram_buffer(22402) := X"00621021";
        ram_buffer(22403) := X"94420000";
        ram_buffer(22404) := X"8EE4000C";
        ram_buffer(22405) := X"00021027";
        ram_buffer(22406) := X"3042FFFF";
        ram_buffer(22407) := X"AEF20018";
        ram_buffer(22408) := X"1480FF40";
        ram_buffer(22409) := X"000213C2";
        ram_buffer(22410) := X"26360001";
        ram_buffer(22411) := X"24030018";
        ram_buffer(22412) := X"00762023";
        ram_buffer(22413) := X"00821004";
        ram_buffer(22414) := X"2AC40008";
        ram_buffer(22415) := X"14800014";
        ram_buffer(22416) := X"02429025";
        ram_buffer(22417) := X"8EE40010";
        ram_buffer(22418) := X"00121403";
        ram_buffer(22419) := X"24850001";
        ram_buffer(22420) := X"AEE50010";
        ram_buffer(22421) := X"A0820000";
        ram_buffer(22422) := X"8EE40014";
        ram_buffer(22423) := X"26D6FFF8";
        ram_buffer(22424) := X"2484FFFF";
        ram_buffer(22425) := X"AEE40014";
        ram_buffer(22426) := X"10800069";
        ram_buffer(22427) := X"305400FF";
        ram_buffer(22428) := X"12900081";
        ram_buffer(22429) := X"00000000";
        ram_buffer(22430) := X"2AC20008";
        ram_buffer(22431) := X"1040FFF1";
        ram_buffer(22432) := X"00129200";
        ram_buffer(22433) := X"2631FFF9";
        ram_buffer(22434) := X"8EF4000C";
        ram_buffer(22435) := X"32360007";
        ram_buffer(22436) := X"AEF20018";
        ram_buffer(22437) := X"1680FF23";
        ram_buffer(22438) := X"AEF6001C";
        ram_buffer(22439) := X"13C0FF21";
        ram_buffer(22440) := X"02C09021";
        ram_buffer(22441) := X"26710001";
        ram_buffer(22442) := X"027EA821";
        ram_buffer(22443) := X"1680001F";
        ram_buffer(22444) := X"26540001";
        ram_buffer(22445) := X"9222FFFF";
        ram_buffer(22446) := X"24030018";
        ram_buffer(22447) := X"0074B023";
        ram_buffer(22448) := X"30420001";
        ram_buffer(22449) := X"8EE50018";
        ram_buffer(22450) := X"02C21004";
        ram_buffer(22451) := X"2A840008";
        ram_buffer(22452) := X"14800013";
        ram_buffer(22453) := X"0045B025";
        ram_buffer(22454) := X"8EE40010";
        ram_buffer(22455) := X"00161403";
        ram_buffer(22456) := X"24850001";
        ram_buffer(22457) := X"AEE50010";
        ram_buffer(22458) := X"A0820000";
        ram_buffer(22459) := X"8EE40014";
        ram_buffer(22460) := X"2694FFF8";
        ram_buffer(22461) := X"2484FFFF";
        ram_buffer(22462) := X"AEE40014";
        ram_buffer(22463) := X"1080007F";
        ram_buffer(22464) := X"305300FF";
        ram_buffer(22465) := X"12700094";
        ram_buffer(22466) := X"00000000";
        ram_buffer(22467) := X"2A820008";
        ram_buffer(22468) := X"1040FFF1";
        ram_buffer(22469) := X"0016B200";
        ram_buffer(22470) := X"2652FFF9";
        ram_buffer(22471) := X"32540007";
        ram_buffer(22472) := X"AEF60018";
        ram_buffer(22473) := X"AEF4001C";
        ram_buffer(22474) := X"02809021";
        ram_buffer(22475) := X"1235FEFD";
        ram_buffer(22476) := X"26310001";
        ram_buffer(22477) := X"8EF4000C";
        ram_buffer(22478) := X"1000FFDC";
        ram_buffer(22479) := X"00000000";
        ram_buffer(22480) := X"8EE40020";
        ram_buffer(22481) := X"00000000";
        ram_buffer(22482) := X"8C850014";
        ram_buffer(22483) := X"00000000";
        ram_buffer(22484) := X"8CA2000C";
        ram_buffer(22485) := X"00000000";
        ram_buffer(22486) := X"0040F809";
        ram_buffer(22487) := X"AFA50110";
        ram_buffer(22488) := X"8FA50110";
        ram_buffer(22489) := X"1440000B";
        ram_buffer(22490) := X"24030016";
        ram_buffer(22491) := X"8EE40020";
        ram_buffer(22492) := X"00000000";
        ram_buffer(22493) := X"8C820000";
        ram_buffer(22494) := X"00000000";
        ram_buffer(22495) := X"8C460000";
        ram_buffer(22496) := X"00000000";
        ram_buffer(22497) := X"00C0F809";
        ram_buffer(22498) := X"AC430014";
        ram_buffer(22499) := X"8FA50110";
        ram_buffer(22500) := X"00000000";
        ram_buffer(22501) := X"8CA40000";
        ram_buffer(22502) := X"8CA20004";
        ram_buffer(22503) := X"AEE40010";
        ram_buffer(22504) := X"16B0FF90";
        ram_buffer(22505) := X"AEE20014";
        ram_buffer(22506) := X"8EE20010";
        ram_buffer(22507) := X"00000000";
        ram_buffer(22508) := X"24440001";
        ram_buffer(22509) := X"AEE40010";
        ram_buffer(22510) := X"A0400000";
        ram_buffer(22511) := X"8EE20014";
        ram_buffer(22512) := X"00000000";
        ram_buffer(22513) := X"2442FFFF";
        ram_buffer(22514) := X"1440FF86";
        ram_buffer(22515) := X"AEE20014";
        ram_buffer(22516) := X"8EE40020";
        ram_buffer(22517) := X"00000000";
        ram_buffer(22518) := X"8C850014";
        ram_buffer(22519) := X"00000000";
        ram_buffer(22520) := X"8CA2000C";
        ram_buffer(22521) := X"00000000";
        ram_buffer(22522) := X"0040F809";
        ram_buffer(22523) := X"AFA50110";
        ram_buffer(22524) := X"8FA50110";
        ram_buffer(22525) := X"104000EE";
        ram_buffer(22526) := X"24030016";
        ram_buffer(22527) := X"8CA40000";
        ram_buffer(22528) := X"8CA20004";
        ram_buffer(22529) := X"AEE40010";
        ram_buffer(22530) := X"1000FF76";
        ram_buffer(22531) := X"AEE20014";
        ram_buffer(22532) := X"8EE40020";
        ram_buffer(22533) := X"00000000";
        ram_buffer(22534) := X"8C850014";
        ram_buffer(22535) := X"00000000";
        ram_buffer(22536) := X"8CA2000C";
        ram_buffer(22537) := X"00000000";
        ram_buffer(22538) := X"0040F809";
        ram_buffer(22539) := X"AFA50110";
        ram_buffer(22540) := X"8FA50110";
        ram_buffer(22541) := X"1440000B";
        ram_buffer(22542) := X"24030016";
        ram_buffer(22543) := X"8EE40020";
        ram_buffer(22544) := X"00000000";
        ram_buffer(22545) := X"8C820000";
        ram_buffer(22546) := X"00000000";
        ram_buffer(22547) := X"8C460000";
        ram_buffer(22548) := X"00000000";
        ram_buffer(22549) := X"00C0F809";
        ram_buffer(22550) := X"AC430014";
        ram_buffer(22551) := X"8FA50110";
        ram_buffer(22552) := X"00000000";
        ram_buffer(22553) := X"8CA40000";
        ram_buffer(22554) := X"8CA20004";
        ram_buffer(22555) := X"AEE40010";
        ram_buffer(22556) := X"1690FF81";
        ram_buffer(22557) := X"AEE20014";
        ram_buffer(22558) := X"8EE20010";
        ram_buffer(22559) := X"00000000";
        ram_buffer(22560) := X"24440001";
        ram_buffer(22561) := X"AEE40010";
        ram_buffer(22562) := X"A0400000";
        ram_buffer(22563) := X"8EE20014";
        ram_buffer(22564) := X"00000000";
        ram_buffer(22565) := X"2442FFFF";
        ram_buffer(22566) := X"1440FF77";
        ram_buffer(22567) := X"AEE20014";
        ram_buffer(22568) := X"8EE40020";
        ram_buffer(22569) := X"00000000";
        ram_buffer(22570) := X"8C940014";
        ram_buffer(22571) := X"00000000";
        ram_buffer(22572) := X"8E82000C";
        ram_buffer(22573) := X"00000000";
        ram_buffer(22574) := X"0040F809";
        ram_buffer(22575) := X"00000000";
        ram_buffer(22576) := X"14400009";
        ram_buffer(22577) := X"24030016";
        ram_buffer(22578) := X"8EE40020";
        ram_buffer(22579) := X"00000000";
        ram_buffer(22580) := X"8C820000";
        ram_buffer(22581) := X"00000000";
        ram_buffer(22582) := X"8C450000";
        ram_buffer(22583) := X"00000000";
        ram_buffer(22584) := X"00A0F809";
        ram_buffer(22585) := X"AC430014";
        ram_buffer(22586) := X"8E840000";
        ram_buffer(22587) := X"8E820004";
        ram_buffer(22588) := X"AEE40010";
        ram_buffer(22589) := X"1000FF60";
        ram_buffer(22590) := X"AEE20014";
        ram_buffer(22591) := X"8EE40020";
        ram_buffer(22592) := X"00000000";
        ram_buffer(22593) := X"8C9E0014";
        ram_buffer(22594) := X"00000000";
        ram_buffer(22595) := X"8FC2000C";
        ram_buffer(22596) := X"00000000";
        ram_buffer(22597) := X"0040F809";
        ram_buffer(22598) := X"00000000";
        ram_buffer(22599) := X"14400009";
        ram_buffer(22600) := X"24030016";
        ram_buffer(22601) := X"8EE40020";
        ram_buffer(22602) := X"00000000";
        ram_buffer(22603) := X"8C820000";
        ram_buffer(22604) := X"00000000";
        ram_buffer(22605) := X"8C460000";
        ram_buffer(22606) := X"00000000";
        ram_buffer(22607) := X"00C0F809";
        ram_buffer(22608) := X"AC430014";
        ram_buffer(22609) := X"8FC40000";
        ram_buffer(22610) := X"8FC20004";
        ram_buffer(22611) := X"AEE40010";
        ram_buffer(22612) := X"1670FF6E";
        ram_buffer(22613) := X"AEE20014";
        ram_buffer(22614) := X"8EE20010";
        ram_buffer(22615) := X"00000000";
        ram_buffer(22616) := X"24440001";
        ram_buffer(22617) := X"AEE40010";
        ram_buffer(22618) := X"A0400000";
        ram_buffer(22619) := X"8EE20014";
        ram_buffer(22620) := X"00000000";
        ram_buffer(22621) := X"2442FFFF";
        ram_buffer(22622) := X"1440FF64";
        ram_buffer(22623) := X"AEE20014";
        ram_buffer(22624) := X"8EE40020";
        ram_buffer(22625) := X"00000000";
        ram_buffer(22626) := X"8C930014";
        ram_buffer(22627) := X"00000000";
        ram_buffer(22628) := X"8E62000C";
        ram_buffer(22629) := X"00000000";
        ram_buffer(22630) := X"0040F809";
        ram_buffer(22631) := X"00000000";
        ram_buffer(22632) := X"14400009";
        ram_buffer(22633) := X"24030016";
        ram_buffer(22634) := X"8EE40020";
        ram_buffer(22635) := X"00000000";
        ram_buffer(22636) := X"8C820000";
        ram_buffer(22637) := X"00000000";
        ram_buffer(22638) := X"8C450000";
        ram_buffer(22639) := X"00000000";
        ram_buffer(22640) := X"00A0F809";
        ram_buffer(22641) := X"AC430014";
        ram_buffer(22642) := X"8E640000";
        ram_buffer(22643) := X"8E620004";
        ram_buffer(22644) := X"AEE40010";
        ram_buffer(22645) := X"1000FF4D";
        ram_buffer(22646) := X"AEE20014";
        ram_buffer(22647) := X"8EE40020";
        ram_buffer(22648) := X"24030027";
        ram_buffer(22649) := X"8C850000";
        ram_buffer(22650) := X"00000000";
        ram_buffer(22651) := X"8CA20000";
        ram_buffer(22652) := X"00000000";
        ram_buffer(22653) := X"0040F809";
        ram_buffer(22654) := X"ACA30014";
        ram_buffer(22655) := X"8EE2000C";
        ram_buffer(22656) := X"00000000";
        ram_buffer(22657) := X"1440FE47";
        ram_buffer(22658) := X"24020001";
        ram_buffer(22659) := X"02221004";
        ram_buffer(22660) := X"2442FFFF";
        ram_buffer(22661) := X"02368821";
        ram_buffer(22662) := X"24030018";
        ram_buffer(22663) := X"00521024";
        ram_buffer(22664) := X"8EE50018";
        ram_buffer(22665) := X"00719023";
        ram_buffer(22666) := X"02421004";
        ram_buffer(22667) := X"2A240008";
        ram_buffer(22668) := X"1080FEDD";
        ram_buffer(22669) := X"00459025";
        ram_buffer(22670) := X"8FA20128";
        ram_buffer(22671) := X"AEF1001C";
        ram_buffer(22672) := X"8C420000";
        ram_buffer(22673) := X"8FA30130";
        ram_buffer(22674) := X"00021040";
        ram_buffer(22675) := X"00621021";
        ram_buffer(22676) := X"94420000";
        ram_buffer(22677) := X"AEF20018";
        ram_buffer(22678) := X"00021027";
        ram_buffer(22679) := X"3042FFFF";
        ram_buffer(22680) := X"1000FEF1";
        ram_buffer(22681) := X"000213C2";
        ram_buffer(22682) := X"8EE40020";
        ram_buffer(22683) := X"24030027";
        ram_buffer(22684) := X"8C870000";
        ram_buffer(22685) := X"00000000";
        ram_buffer(22686) := X"8CE20000";
        ram_buffer(22687) := X"00000000";
        ram_buffer(22688) := X"0040F809";
        ram_buffer(22689) := X"ACE30014";
        ram_buffer(22690) := X"8EE2000C";
        ram_buffer(22691) := X"00000000";
        ram_buffer(22692) := X"1440FE12";
        ram_buffer(22693) := X"24020001";
        ram_buffer(22694) := X"1000FE36";
        ram_buffer(22695) := X"02221004";
        ram_buffer(22696) := X"8EE40020";
        ram_buffer(22697) := X"00000000";
        ram_buffer(22698) := X"8C850014";
        ram_buffer(22699) := X"00000000";
        ram_buffer(22700) := X"8CA2000C";
        ram_buffer(22701) := X"00000000";
        ram_buffer(22702) := X"0040F809";
        ram_buffer(22703) := X"AFA50110";
        ram_buffer(22704) := X"8FA50110";
        ram_buffer(22705) := X"1440000B";
        ram_buffer(22706) := X"24030016";
        ram_buffer(22707) := X"8EE40020";
        ram_buffer(22708) := X"00000000";
        ram_buffer(22709) := X"8C820000";
        ram_buffer(22710) := X"00000000";
        ram_buffer(22711) := X"8C460000";
        ram_buffer(22712) := X"00000000";
        ram_buffer(22713) := X"00C0F809";
        ram_buffer(22714) := X"AC430014";
        ram_buffer(22715) := X"8FA50110";
        ram_buffer(22716) := X"00000000";
        ram_buffer(22717) := X"8CA40000";
        ram_buffer(22718) := X"8CA20004";
        ram_buffer(22719) := X"AEE40010";
        ram_buffer(22720) := X"16B0FE58";
        ram_buffer(22721) := X"AEE20014";
        ram_buffer(22722) := X"8EE20010";
        ram_buffer(22723) := X"00000000";
        ram_buffer(22724) := X"24440001";
        ram_buffer(22725) := X"AEE40010";
        ram_buffer(22726) := X"A0400000";
        ram_buffer(22727) := X"8EE20014";
        ram_buffer(22728) := X"00000000";
        ram_buffer(22729) := X"2442FFFF";
        ram_buffer(22730) := X"1440FE4E";
        ram_buffer(22731) := X"AEE20014";
        ram_buffer(22732) := X"8EE40020";
        ram_buffer(22733) := X"00000000";
        ram_buffer(22734) := X"8C850014";
        ram_buffer(22735) := X"00000000";
        ram_buffer(22736) := X"8CA2000C";
        ram_buffer(22737) := X"00000000";
        ram_buffer(22738) := X"0040F809";
        ram_buffer(22739) := X"AFA50110";
        ram_buffer(22740) := X"8FA50110";
        ram_buffer(22741) := X"1040000B";
        ram_buffer(22742) := X"24030016";
        ram_buffer(22743) := X"8CA40000";
        ram_buffer(22744) := X"8CA20004";
        ram_buffer(22745) := X"AEE40010";
        ram_buffer(22746) := X"1000FE3E";
        ram_buffer(22747) := X"AEE20014";
        ram_buffer(22748) := X"8EE50048";
        ram_buffer(22749) := X"0C02502F";
        ram_buffer(22750) := X"02E02021";
        ram_buffer(22751) := X"1000FB3A";
        ram_buffer(22752) := X"00000000";
        ram_buffer(22753) := X"8EE40020";
        ram_buffer(22754) := X"00000000";
        ram_buffer(22755) := X"8C820000";
        ram_buffer(22756) := X"00000000";
        ram_buffer(22757) := X"8C460000";
        ram_buffer(22758) := X"00000000";
        ram_buffer(22759) := X"00C0F809";
        ram_buffer(22760) := X"AC430014";
        ram_buffer(22761) := X"8FA50110";
        ram_buffer(22762) := X"1000FFEC";
        ram_buffer(22763) := X"00000000";
        ram_buffer(22764) := X"8EE40020";
        ram_buffer(22765) := X"00000000";
        ram_buffer(22766) := X"8C820000";
        ram_buffer(22767) := X"00000000";
        ram_buffer(22768) := X"8C460000";
        ram_buffer(22769) := X"00000000";
        ram_buffer(22770) := X"00C0F809";
        ram_buffer(22771) := X"AC430014";
        ram_buffer(22772) := X"8FA50110";
        ram_buffer(22773) := X"1000FF09";
        ram_buffer(22774) := X"00000000";
        ram_buffer(22775) := X"8EE40020";
        ram_buffer(22776) := X"00000000";
        ram_buffer(22777) := X"8C820000";
        ram_buffer(22778) := X"00000000";
        ram_buffer(22779) := X"8C470000";
        ram_buffer(22780) := X"00000000";
        ram_buffer(22781) := X"00E0F809";
        ram_buffer(22782) := X"AC430014";
        ram_buffer(22783) := X"8FA60110";
        ram_buffer(22784) := X"1000FE4D";
        ram_buffer(22785) := X"00000000";
        ram_buffer(22786) := X"1000FDA6";
        ram_buffer(22787) := X"0000A021";
        ram_buffer(22788) := X"8FA20110";
        ram_buffer(22789) := X"00000000";
        ram_buffer(22790) := X"1040FBB5";
        ram_buffer(22791) := X"00000000";
        ram_buffer(22792) := X"1000FBA5";
        ram_buffer(22793) := X"00000000";
        ram_buffer(22794) := X"8C820014";
        ram_buffer(22795) := X"27BDFFA0";
        ram_buffer(22796) := X"00801821";
        ram_buffer(22797) := X"8C460000";
        ram_buffer(22798) := X"AFBE0058";
        ram_buffer(22799) := X"AFA40060";
        ram_buffer(22800) := X"8C9E0164";
        ram_buffer(22801) := X"8C440004";
        ram_buffer(22802) := X"8C6200C0";
        ram_buffer(22803) := X"8C630138";
        ram_buffer(22804) := X"AFB00038";
        ram_buffer(22805) := X"AFA3001C";
        ram_buffer(22806) := X"8FA30060";
        ram_buffer(22807) := X"AFBF005C";
        ram_buffer(22808) := X"8C630140";
        ram_buffer(22809) := X"AFB70054";
        ram_buffer(22810) := X"AFB60050";
        ram_buffer(22811) := X"AFB5004C";
        ram_buffer(22812) := X"AFB40048";
        ram_buffer(22813) := X"AFB30044";
        ram_buffer(22814) := X"AFB20040";
        ram_buffer(22815) := X"AFB1003C";
        ram_buffer(22816) := X"AFA3002C";
        ram_buffer(22817) := X"00A08021";
        ram_buffer(22818) := X"AFC60010";
        ram_buffer(22819) := X"10400005";
        ram_buffer(22820) := X"AFC40014";
        ram_buffer(22821) := X"8FC20044";
        ram_buffer(22822) := X"00000000";
        ram_buffer(22823) := X"104001F7";
        ram_buffer(22824) := X"00000000";
        ram_buffer(22825) := X"8FA20060";
        ram_buffer(22826) := X"8E030000";
        ram_buffer(22827) := X"8C420134";
        ram_buffer(22828) := X"8FA4001C";
        ram_buffer(22829) := X"AFA20014";
        ram_buffer(22830) := X"AFA30020";
        ram_buffer(22831) := X"00401821";
        ram_buffer(22832) := X"0082102A";
        ram_buffer(22833) := X"1440005D";
        ram_buffer(22834) := X"3C02100D";
        ram_buffer(22835) := X"0003A080";
        ram_buffer(22836) := X"24428968";
        ram_buffer(22837) := X"0054A021";
        ram_buffer(22838) := X"AFA00010";
        ram_buffer(22839) := X"241100FF";
        ram_buffer(22840) := X"8E820000";
        ram_buffer(22841) := X"8FA30020";
        ram_buffer(22842) := X"00021040";
        ram_buffer(22843) := X"00621021";
        ram_buffer(22844) := X"84500000";
        ram_buffer(22845) := X"00000000";
        ram_buffer(22846) := X"1200006C";
        ram_buffer(22847) := X"00000000";
        ram_buffer(22848) := X"060000E6";
        ram_buffer(22849) := X"00000000";
        ram_buffer(22850) := X"8FA2002C";
        ram_buffer(22851) := X"00000000";
        ram_buffer(22852) := X"00501007";
        ram_buffer(22853) := X"AFA20018";
        ram_buffer(22854) := X"AFA20028";
        ram_buffer(22855) := X"10400063";
        ram_buffer(22856) := X"00000000";
        ram_buffer(22857) := X"8FC20038";
        ram_buffer(22858) := X"00000000";
        ram_buffer(22859) := X"144001AB";
        ram_buffer(22860) := X"00021043";
        ram_buffer(22861) := X"8FA20010";
        ram_buffer(22862) := X"8FC40034";
        ram_buffer(22863) := X"28420010";
        ram_buffer(22864) := X"8FC7000C";
        ram_buffer(22865) := X"8FD2001C";
        ram_buffer(22866) := X"14400014";
        ram_buffer(22867) := X"00000000";
        ram_buffer(22868) := X"8FB70010";
        ram_buffer(22869) := X"10E0005A";
        ram_buffer(22870) := X"24820016";
        ram_buffer(22871) := X"00021080";
        ram_buffer(22872) := X"03C21021";
        ram_buffer(22873) := X"8C450004";
        ram_buffer(22874) := X"00000000";
        ram_buffer(22875) := X"8CA203C0";
        ram_buffer(22876) := X"00000000";
        ram_buffer(22877) := X"24420001";
        ram_buffer(22878) := X"ACA203C0";
        ram_buffer(22879) := X"26F7FFF0";
        ram_buffer(22880) := X"2AE20010";
        ram_buffer(22881) := X"1040FFF3";
        ram_buffer(22882) := X"00000000";
        ram_buffer(22883) := X"8FA20010";
        ram_buffer(22884) := X"00000000";
        ram_buffer(22885) := X"3042000F";
        ram_buffer(22886) := X"AFA20010";
        ram_buffer(22887) := X"8FA20018";
        ram_buffer(22888) := X"00000000";
        ram_buffer(22889) := X"00028043";
        ram_buffer(22890) := X"12000004";
        ram_buffer(22891) := X"24050001";
        ram_buffer(22892) := X"00108043";
        ram_buffer(22893) := X"1600FFFE";
        ram_buffer(22894) := X"24A50001";
        ram_buffer(22895) := X"8FA20010";
        ram_buffer(22896) := X"00000000";
        ram_buffer(22897) := X"00029900";
        ram_buffer(22898) := X"10E000BD";
        ram_buffer(22899) := X"02659821";
        ram_buffer(22900) := X"24820016";
        ram_buffer(22901) := X"00021080";
        ram_buffer(22902) := X"03C21021";
        ram_buffer(22903) := X"8C420004";
        ram_buffer(22904) := X"00139880";
        ram_buffer(22905) := X"00539821";
        ram_buffer(22906) := X"8E620000";
        ram_buffer(22907) := X"00000000";
        ram_buffer(22908) := X"24420001";
        ram_buffer(22909) := X"AE620000";
        ram_buffer(22910) := X"AFA00010";
        ram_buffer(22911) := X"8FA20014";
        ram_buffer(22912) := X"8FA3001C";
        ram_buffer(22913) := X"24420001";
        ram_buffer(22914) := X"AFA20014";
        ram_buffer(22915) := X"0062102A";
        ram_buffer(22916) := X"1040FFB3";
        ram_buffer(22917) := X"26940004";
        ram_buffer(22918) := X"8FA20010";
        ram_buffer(22919) := X"00000000";
        ram_buffer(22920) := X"10400006";
        ram_buffer(22921) := X"24047FFF";
        ram_buffer(22922) := X"8FC20038";
        ram_buffer(22923) := X"00000000";
        ram_buffer(22924) := X"24420001";
        ram_buffer(22925) := X"10440255";
        ram_buffer(22926) := X"AFC20038";
        ram_buffer(22927) := X"8FA20060";
        ram_buffer(22928) := X"8FA30060";
        ram_buffer(22929) := X"8C420014";
        ram_buffer(22930) := X"8FC60010";
        ram_buffer(22931) := X"8FC50014";
        ram_buffer(22932) := X"8C6400C0";
        ram_buffer(22933) := X"AC460000";
        ram_buffer(22934) := X"10800007";
        ram_buffer(22935) := X"AC450004";
        ram_buffer(22936) := X"8FC20044";
        ram_buffer(22937) := X"00000000";
        ram_buffer(22938) := X"10400156";
        ram_buffer(22939) := X"00000000";
        ram_buffer(22940) := X"2442FFFF";
        ram_buffer(22941) := X"AFC20044";
        ram_buffer(22942) := X"8FBF005C";
        ram_buffer(22943) := X"8FBE0058";
        ram_buffer(22944) := X"8FB70054";
        ram_buffer(22945) := X"8FB60050";
        ram_buffer(22946) := X"8FB5004C";
        ram_buffer(22947) := X"8FB40048";
        ram_buffer(22948) := X"8FB30044";
        ram_buffer(22949) := X"8FB20040";
        ram_buffer(22950) := X"8FB1003C";
        ram_buffer(22951) := X"8FB00038";
        ram_buffer(22952) := X"24020001";
        ram_buffer(22953) := X"03E00008";
        ram_buffer(22954) := X"27BD0060";
        ram_buffer(22955) := X"8FA20010";
        ram_buffer(22956) := X"00000000";
        ram_buffer(22957) := X"24420001";
        ram_buffer(22958) := X"1000FFD0";
        ram_buffer(22959) := X"AFA20010";
        ram_buffer(22960) := X"24840012";
        ram_buffer(22961) := X"00042080";
        ram_buffer(22962) := X"03C42021";
        ram_buffer(22963) := X"8C820004";
        ram_buffer(22964) := X"00000000";
        ram_buffer(22965) := X"805604F0";
        ram_buffer(22966) := X"8C5003C0";
        ram_buffer(22967) := X"12C0005F";
        ram_buffer(22968) := X"24030027";
        ram_buffer(22969) := X"24020001";
        ram_buffer(22970) := X"02C21004";
        ram_buffer(22971) := X"02D29021";
        ram_buffer(22972) := X"2442FFFF";
        ram_buffer(22973) := X"24030018";
        ram_buffer(22974) := X"00501024";
        ram_buffer(22975) := X"00723023";
        ram_buffer(22976) := X"8FC50018";
        ram_buffer(22977) := X"00C21004";
        ram_buffer(22978) := X"2A440008";
        ram_buffer(22979) := X"14800014";
        ram_buffer(22980) := X"0045B025";
        ram_buffer(22981) := X"02408021";
        ram_buffer(22982) := X"8FC40010";
        ram_buffer(22983) := X"00161403";
        ram_buffer(22984) := X"24850001";
        ram_buffer(22985) := X"AFC50010";
        ram_buffer(22986) := X"A0820000";
        ram_buffer(22987) := X"8FC40014";
        ram_buffer(22988) := X"2610FFF8";
        ram_buffer(22989) := X"2484FFFF";
        ram_buffer(22990) := X"AFC40014";
        ram_buffer(22991) := X"1080000C";
        ram_buffer(22992) := X"305300FF";
        ram_buffer(22993) := X"12710021";
        ram_buffer(22994) := X"00000000";
        ram_buffer(22995) := X"2A020008";
        ram_buffer(22996) := X"1040FFF1";
        ram_buffer(22997) := X"0016B200";
        ram_buffer(22998) := X"8FC7000C";
        ram_buffer(22999) := X"32520007";
        ram_buffer(23000) := X"8FC40034";
        ram_buffer(23001) := X"AFD60018";
        ram_buffer(23002) := X"1000FF84";
        ram_buffer(23003) := X"AFD2001C";
        ram_buffer(23004) := X"8FC40020";
        ram_buffer(23005) := X"00000000";
        ram_buffer(23006) := X"8C950014";
        ram_buffer(23007) := X"00000000";
        ram_buffer(23008) := X"8EA2000C";
        ram_buffer(23009) := X"00000000";
        ram_buffer(23010) := X"0040F809";
        ram_buffer(23011) := X"00000000";
        ram_buffer(23012) := X"14400009";
        ram_buffer(23013) := X"24030016";
        ram_buffer(23014) := X"8FC40020";
        ram_buffer(23015) := X"00000000";
        ram_buffer(23016) := X"8C820000";
        ram_buffer(23017) := X"00000000";
        ram_buffer(23018) := X"8C4A0000";
        ram_buffer(23019) := X"00000000";
        ram_buffer(23020) := X"0140F809";
        ram_buffer(23021) := X"AC430014";
        ram_buffer(23022) := X"8EA40000";
        ram_buffer(23023) := X"8EA20004";
        ram_buffer(23024) := X"AFC40010";
        ram_buffer(23025) := X"1671FFE1";
        ram_buffer(23026) := X"AFC20014";
        ram_buffer(23027) := X"8FC20010";
        ram_buffer(23028) := X"00000000";
        ram_buffer(23029) := X"24440001";
        ram_buffer(23030) := X"AFC40010";
        ram_buffer(23031) := X"A0400000";
        ram_buffer(23032) := X"8FC20014";
        ram_buffer(23033) := X"00000000";
        ram_buffer(23034) := X"2442FFFF";
        ram_buffer(23035) := X"1440FFD7";
        ram_buffer(23036) := X"AFC20014";
        ram_buffer(23037) := X"8FC40020";
        ram_buffer(23038) := X"00000000";
        ram_buffer(23039) := X"8C850014";
        ram_buffer(23040) := X"00000000";
        ram_buffer(23041) := X"8CA2000C";
        ram_buffer(23042) := X"00000000";
        ram_buffer(23043) := X"0040F809";
        ram_buffer(23044) := X"AFA50024";
        ram_buffer(23045) := X"8FA50024";
        ram_buffer(23046) := X"1440000B";
        ram_buffer(23047) := X"24030016";
        ram_buffer(23048) := X"8FC40020";
        ram_buffer(23049) := X"00000000";
        ram_buffer(23050) := X"8C820000";
        ram_buffer(23051) := X"00000000";
        ram_buffer(23052) := X"8C490000";
        ram_buffer(23053) := X"00000000";
        ram_buffer(23054) := X"0120F809";
        ram_buffer(23055) := X"AC430014";
        ram_buffer(23056) := X"8FA50024";
        ram_buffer(23057) := X"00000000";
        ram_buffer(23058) := X"8CA40000";
        ram_buffer(23059) := X"8CA20004";
        ram_buffer(23060) := X"AFC40010";
        ram_buffer(23061) := X"1000FFBD";
        ram_buffer(23062) := X"AFC20014";
        ram_buffer(23063) := X"8FC40020";
        ram_buffer(23064) := X"00000000";
        ram_buffer(23065) := X"8C820000";
        ram_buffer(23066) := X"AFA70024";
        ram_buffer(23067) := X"8C490000";
        ram_buffer(23068) := X"00000000";
        ram_buffer(23069) := X"0120F809";
        ram_buffer(23070) := X"AC430014";
        ram_buffer(23071) := X"8FC2000C";
        ram_buffer(23072) := X"8FA70024";
        ram_buffer(23073) := X"1040FF97";
        ram_buffer(23074) := X"00000000";
        ram_buffer(23075) := X"8FC40034";
        ram_buffer(23076) := X"8FD2001C";
        ram_buffer(23077) := X"1000FF39";
        ram_buffer(23078) := X"00403821";
        ram_buffer(23079) := X"8FA2002C";
        ram_buffer(23080) := X"00108023";
        ram_buffer(23081) := X"00501007";
        ram_buffer(23082) := X"AFA20018";
        ram_buffer(23083) := X"00021027";
        ram_buffer(23084) := X"AFA20028";
        ram_buffer(23085) := X"8FA20018";
        ram_buffer(23086) := X"1000FF18";
        ram_buffer(23087) := X"00000000";
        ram_buffer(23088) := X"24820012";
        ram_buffer(23089) := X"00021080";
        ram_buffer(23090) := X"03C21021";
        ram_buffer(23091) := X"8C420004";
        ram_buffer(23092) := X"00132080";
        ram_buffer(23093) := X"00539821";
        ram_buffer(23094) := X"82700400";
        ram_buffer(23095) := X"00441021";
        ram_buffer(23096) := X"8C530000";
        ram_buffer(23097) := X"120000D6";
        ram_buffer(23098) := X"24020001";
        ram_buffer(23099) := X"02021004";
        ram_buffer(23100) := X"0212A821";
        ram_buffer(23101) := X"2442FFFF";
        ram_buffer(23102) := X"24030018";
        ram_buffer(23103) := X"00531024";
        ram_buffer(23104) := X"00752023";
        ram_buffer(23105) := X"8FD30018";
        ram_buffer(23106) := X"00821004";
        ram_buffer(23107) := X"2AA40008";
        ram_buffer(23108) := X"14800014";
        ram_buffer(23109) := X"00539825";
        ram_buffer(23110) := X"02A08021";
        ram_buffer(23111) := X"8FC40010";
        ram_buffer(23112) := X"00131403";
        ram_buffer(23113) := X"24870001";
        ram_buffer(23114) := X"AFC70010";
        ram_buffer(23115) := X"A0820000";
        ram_buffer(23116) := X"8FC40014";
        ram_buffer(23117) := X"2610FFF8";
        ram_buffer(23118) := X"2484FFFF";
        ram_buffer(23119) := X"AFC40014";
        ram_buffer(23120) := X"1080002C";
        ram_buffer(23121) := X"305200FF";
        ram_buffer(23122) := X"12510043";
        ram_buffer(23123) := X"00000000";
        ram_buffer(23124) := X"2A020008";
        ram_buffer(23125) := X"1040FFF1";
        ram_buffer(23126) := X"00139A00";
        ram_buffer(23127) := X"8FC7000C";
        ram_buffer(23128) := X"32B50007";
        ram_buffer(23129) := X"AFD30018";
        ram_buffer(23130) := X"14E0FF23";
        ram_buffer(23131) := X"AFD5001C";
        ram_buffer(23132) := X"24020001";
        ram_buffer(23133) := X"8FA30028";
        ram_buffer(23134) := X"00A21004";
        ram_buffer(23135) := X"2442FFFF";
        ram_buffer(23136) := X"00B5A821";
        ram_buffer(23137) := X"00431024";
        ram_buffer(23138) := X"24030018";
        ram_buffer(23139) := X"00752023";
        ram_buffer(23140) := X"00821004";
        ram_buffer(23141) := X"2AA40008";
        ram_buffer(23142) := X"14800013";
        ram_buffer(23143) := X"00539825";
        ram_buffer(23144) := X"02A08021";
        ram_buffer(23145) := X"8FC40010";
        ram_buffer(23146) := X"00131403";
        ram_buffer(23147) := X"24860001";
        ram_buffer(23148) := X"AFC60010";
        ram_buffer(23149) := X"A0820000";
        ram_buffer(23150) := X"8FC40014";
        ram_buffer(23151) := X"2610FFF8";
        ram_buffer(23152) := X"2484FFFF";
        ram_buffer(23153) := X"AFC40014";
        ram_buffer(23154) := X"10800046";
        ram_buffer(23155) := X"305200FF";
        ram_buffer(23156) := X"1251005B";
        ram_buffer(23157) := X"00000000";
        ram_buffer(23158) := X"2A020008";
        ram_buffer(23159) := X"1040FFF1";
        ram_buffer(23160) := X"00139A00";
        ram_buffer(23161) := X"32B50007";
        ram_buffer(23162) := X"AFD30018";
        ram_buffer(23163) := X"1000FF02";
        ram_buffer(23164) := X"AFD5001C";
        ram_buffer(23165) := X"8FC40020";
        ram_buffer(23166) := X"AFA50010";
        ram_buffer(23167) := X"8C970014";
        ram_buffer(23168) := X"00000000";
        ram_buffer(23169) := X"8EE2000C";
        ram_buffer(23170) := X"00000000";
        ram_buffer(23171) := X"0040F809";
        ram_buffer(23172) := X"00000000";
        ram_buffer(23173) := X"8FA50010";
        ram_buffer(23174) := X"1440000A";
        ram_buffer(23175) := X"24030016";
        ram_buffer(23176) := X"8FC40020";
        ram_buffer(23177) := X"00000000";
        ram_buffer(23178) := X"8C820000";
        ram_buffer(23179) := X"00000000";
        ram_buffer(23180) := X"8C480000";
        ram_buffer(23181) := X"00000000";
        ram_buffer(23182) := X"0100F809";
        ram_buffer(23183) := X"AC430014";
        ram_buffer(23184) := X"8FA50010";
        ram_buffer(23185) := X"8EE40000";
        ram_buffer(23186) := X"8EE20004";
        ram_buffer(23187) := X"AFC40010";
        ram_buffer(23188) := X"1651FFBF";
        ram_buffer(23189) := X"AFC20014";
        ram_buffer(23190) := X"8FC20010";
        ram_buffer(23191) := X"00000000";
        ram_buffer(23192) := X"24440001";
        ram_buffer(23193) := X"AFC40010";
        ram_buffer(23194) := X"A0400000";
        ram_buffer(23195) := X"8FC20014";
        ram_buffer(23196) := X"00000000";
        ram_buffer(23197) := X"2442FFFF";
        ram_buffer(23198) := X"1440FFB5";
        ram_buffer(23199) := X"AFC20014";
        ram_buffer(23200) := X"8FC40020";
        ram_buffer(23201) := X"AFA50010";
        ram_buffer(23202) := X"8C920014";
        ram_buffer(23203) := X"00000000";
        ram_buffer(23204) := X"8E42000C";
        ram_buffer(23205) := X"00000000";
        ram_buffer(23206) := X"0040F809";
        ram_buffer(23207) := X"00000000";
        ram_buffer(23208) := X"8FA50010";
        ram_buffer(23209) := X"1440000A";
        ram_buffer(23210) := X"24030016";
        ram_buffer(23211) := X"8FC40020";
        ram_buffer(23212) := X"00000000";
        ram_buffer(23213) := X"8C820000";
        ram_buffer(23214) := X"00000000";
        ram_buffer(23215) := X"8C470000";
        ram_buffer(23216) := X"00000000";
        ram_buffer(23217) := X"00E0F809";
        ram_buffer(23218) := X"AC430014";
        ram_buffer(23219) := X"8FA50010";
        ram_buffer(23220) := X"8E440000";
        ram_buffer(23221) := X"8E420004";
        ram_buffer(23222) := X"AFC40010";
        ram_buffer(23223) := X"1000FF9C";
        ram_buffer(23224) := X"AFC20014";
        ram_buffer(23225) := X"8FC40020";
        ram_buffer(23226) := X"00000000";
        ram_buffer(23227) := X"8C970014";
        ram_buffer(23228) := X"00000000";
        ram_buffer(23229) := X"8EE2000C";
        ram_buffer(23230) := X"00000000";
        ram_buffer(23231) := X"0040F809";
        ram_buffer(23232) := X"00000000";
        ram_buffer(23233) := X"14400009";
        ram_buffer(23234) := X"24030016";
        ram_buffer(23235) := X"8FC40020";
        ram_buffer(23236) := X"00000000";
        ram_buffer(23237) := X"8C820000";
        ram_buffer(23238) := X"00000000";
        ram_buffer(23239) := X"8C470000";
        ram_buffer(23240) := X"00000000";
        ram_buffer(23241) := X"00E0F809";
        ram_buffer(23242) := X"AC430014";
        ram_buffer(23243) := X"8EE40000";
        ram_buffer(23244) := X"8EE20004";
        ram_buffer(23245) := X"AFC40010";
        ram_buffer(23246) := X"1651FFA7";
        ram_buffer(23247) := X"AFC20014";
        ram_buffer(23248) := X"8FC20010";
        ram_buffer(23249) := X"00000000";
        ram_buffer(23250) := X"24440001";
        ram_buffer(23251) := X"AFC40010";
        ram_buffer(23252) := X"A0400000";
        ram_buffer(23253) := X"8FC20014";
        ram_buffer(23254) := X"00000000";
        ram_buffer(23255) := X"2442FFFF";
        ram_buffer(23256) := X"1440FF9D";
        ram_buffer(23257) := X"AFC20014";
        ram_buffer(23258) := X"8FC40020";
        ram_buffer(23259) := X"00000000";
        ram_buffer(23260) := X"8C920014";
        ram_buffer(23261) := X"00000000";
        ram_buffer(23262) := X"8E42000C";
        ram_buffer(23263) := X"00000000";
        ram_buffer(23264) := X"0040F809";
        ram_buffer(23265) := X"00000000";
        ram_buffer(23266) := X"14400009";
        ram_buffer(23267) := X"24030016";
        ram_buffer(23268) := X"8FC40020";
        ram_buffer(23269) := X"00000000";
        ram_buffer(23270) := X"8C820000";
        ram_buffer(23271) := X"00000000";
        ram_buffer(23272) := X"8C460000";
        ram_buffer(23273) := X"00000000";
        ram_buffer(23274) := X"00C0F809";
        ram_buffer(23275) := X"AC430014";
        ram_buffer(23276) := X"8E440000";
        ram_buffer(23277) := X"8E420004";
        ram_buffer(23278) := X"AFC40010";
        ram_buffer(23279) := X"1000FF86";
        ram_buffer(23280) := X"AFC20014";
        ram_buffer(23281) := X"8FC50048";
        ram_buffer(23282) := X"00801021";
        ram_buffer(23283) := X"24A40001";
        ram_buffer(23284) := X"30840007";
        ram_buffer(23285) := X"1000FEA6";
        ram_buffer(23286) := X"AFC40048";
        ram_buffer(23287) := X"10400108";
        ram_buffer(23288) := X"00002021";
        ram_buffer(23289) := X"00002821";
        ram_buffer(23290) := X"00021043";
        ram_buffer(23291) := X"1440FFFE";
        ram_buffer(23292) := X"24A50001";
        ram_buffer(23293) := X"00052100";
        ram_buffer(23294) := X"8FC6000C";
        ram_buffer(23295) := X"8FC20034";
        ram_buffer(23296) := X"10C00023";
        ram_buffer(23297) := X"00043080";
        ram_buffer(23298) := X"24420016";
        ram_buffer(23299) := X"00021080";
        ram_buffer(23300) := X"03C21021";
        ram_buffer(23301) := X"8C420004";
        ram_buffer(23302) := X"00042080";
        ram_buffer(23303) := X"00442021";
        ram_buffer(23304) := X"8C820000";
        ram_buffer(23305) := X"00000000";
        ram_buffer(23306) := X"24420001";
        ram_buffer(23307) := X"AC820000";
        ram_buffer(23308) := X"0C024B01";
        ram_buffer(23309) := X"03C02021";
        ram_buffer(23310) := X"1000FE3E";
        ram_buffer(23311) := X"00000000";
        ram_buffer(23312) := X"8FC40020";
        ram_buffer(23313) := X"24030027";
        ram_buffer(23314) := X"8C820000";
        ram_buffer(23315) := X"AFA70018";
        ram_buffer(23316) := X"8C460000";
        ram_buffer(23317) := X"AC430014";
        ram_buffer(23318) := X"00C0F809";
        ram_buffer(23319) := X"AFA50010";
        ram_buffer(23320) := X"8FC2000C";
        ram_buffer(23321) := X"8FA50010";
        ram_buffer(23322) := X"8FA70018";
        ram_buffer(23323) := X"1440FE62";
        ram_buffer(23324) := X"24020001";
        ram_buffer(23325) := X"1000FF1E";
        ram_buffer(23326) := X"02021004";
        ram_buffer(23327) := X"8FC50048";
        ram_buffer(23328) := X"0C02502F";
        ram_buffer(23329) := X"03C02021";
        ram_buffer(23330) := X"1000FE06";
        ram_buffer(23331) := X"00000000";
        ram_buffer(23332) := X"24420012";
        ram_buffer(23333) := X"00021080";
        ram_buffer(23334) := X"03C21021";
        ram_buffer(23335) := X"8C420004";
        ram_buffer(23336) := X"00000000";
        ram_buffer(23337) := X"00442021";
        ram_buffer(23338) := X"80920400";
        ram_buffer(23339) := X"00461021";
        ram_buffer(23340) := X"8C570000";
        ram_buffer(23341) := X"8FC7001C";
        ram_buffer(23342) := X"124000B8";
        ram_buffer(23343) := X"24020001";
        ram_buffer(23344) := X"02421004";
        ram_buffer(23345) := X"2442FFFF";
        ram_buffer(23346) := X"02479021";
        ram_buffer(23347) := X"24030018";
        ram_buffer(23348) := X"00571024";
        ram_buffer(23349) := X"00723823";
        ram_buffer(23350) := X"8FC60018";
        ram_buffer(23351) := X"00E21004";
        ram_buffer(23352) := X"2A440008";
        ram_buffer(23353) := X"00463825";
        ram_buffer(23354) := X"14800012";
        ram_buffer(23355) := X"0240B821";
        ram_buffer(23356) := X"8FC40010";
        ram_buffer(23357) := X"00071403";
        ram_buffer(23358) := X"24860001";
        ram_buffer(23359) := X"AFC60010";
        ram_buffer(23360) := X"A0820000";
        ram_buffer(23361) := X"8FC40014";
        ram_buffer(23362) := X"26F7FFF8";
        ram_buffer(23363) := X"2484FFFF";
        ram_buffer(23364) := X"AFC40014";
        ram_buffer(23365) := X"1080002D";
        ram_buffer(23366) := X"305000FF";
        ram_buffer(23367) := X"12110046";
        ram_buffer(23368) := X"00000000";
        ram_buffer(23369) := X"2AE20008";
        ram_buffer(23370) := X"1040FFF1";
        ram_buffer(23371) := X"00073A00";
        ram_buffer(23372) := X"32520007";
        ram_buffer(23373) := X"AFC70018";
        ram_buffer(23374) := X"10A0FFBD";
        ram_buffer(23375) := X"AFD2001C";
        ram_buffer(23376) := X"8FC4000C";
        ram_buffer(23377) := X"8FC60038";
        ram_buffer(23378) := X"1480FFB9";
        ram_buffer(23379) := X"24020001";
        ram_buffer(23380) := X"00A21004";
        ram_buffer(23381) := X"00B2A821";
        ram_buffer(23382) := X"2442FFFF";
        ram_buffer(23383) := X"24030018";
        ram_buffer(23384) := X"00752023";
        ram_buffer(23385) := X"00461024";
        ram_buffer(23386) := X"00821004";
        ram_buffer(23387) := X"2AA40008";
        ram_buffer(23388) := X"14800013";
        ram_buffer(23389) := X"0047B825";
        ram_buffer(23390) := X"02A09021";
        ram_buffer(23391) := X"8FC40010";
        ram_buffer(23392) := X"00171403";
        ram_buffer(23393) := X"24850001";
        ram_buffer(23394) := X"AFC50010";
        ram_buffer(23395) := X"A0820000";
        ram_buffer(23396) := X"8FC40014";
        ram_buffer(23397) := X"2652FFF8";
        ram_buffer(23398) := X"2484FFFF";
        ram_buffer(23399) := X"AFC40014";
        ram_buffer(23400) := X"1080004A";
        ram_buffer(23401) := X"305000FF";
        ram_buffer(23402) := X"1211005F";
        ram_buffer(23403) := X"00000000";
        ram_buffer(23404) := X"2A420008";
        ram_buffer(23405) := X"1040FFF1";
        ram_buffer(23406) := X"0017BA00";
        ram_buffer(23407) := X"32B50007";
        ram_buffer(23408) := X"AFD70018";
        ram_buffer(23409) := X"1000FF9A";
        ram_buffer(23410) := X"AFD5001C";
        ram_buffer(23411) := X"8FC40020";
        ram_buffer(23412) := X"AFA70030";
        ram_buffer(23413) := X"8C930014";
        ram_buffer(23414) := X"AFA50024";
        ram_buffer(23415) := X"8E62000C";
        ram_buffer(23416) := X"00000000";
        ram_buffer(23417) := X"0040F809";
        ram_buffer(23418) := X"00000000";
        ram_buffer(23419) := X"8FA50024";
        ram_buffer(23420) := X"8FA70030";
        ram_buffer(23421) := X"1440000B";
        ram_buffer(23422) := X"24030016";
        ram_buffer(23423) := X"8FC40020";
        ram_buffer(23424) := X"00000000";
        ram_buffer(23425) := X"8C820000";
        ram_buffer(23426) := X"00000000";
        ram_buffer(23427) := X"8C4A0000";
        ram_buffer(23428) := X"00000000";
        ram_buffer(23429) := X"0140F809";
        ram_buffer(23430) := X"AC430014";
        ram_buffer(23431) := X"8FA70030";
        ram_buffer(23432) := X"8FA50024";
        ram_buffer(23433) := X"8E640000";
        ram_buffer(23434) := X"8E620004";
        ram_buffer(23435) := X"AFC40010";
        ram_buffer(23436) := X"1611FFBC";
        ram_buffer(23437) := X"AFC20014";
        ram_buffer(23438) := X"8FC20010";
        ram_buffer(23439) := X"00000000";
        ram_buffer(23440) := X"24440001";
        ram_buffer(23441) := X"AFC40010";
        ram_buffer(23442) := X"A0400000";
        ram_buffer(23443) := X"8FC20014";
        ram_buffer(23444) := X"00000000";
        ram_buffer(23445) := X"2442FFFF";
        ram_buffer(23446) := X"1440FFB2";
        ram_buffer(23447) := X"AFC20014";
        ram_buffer(23448) := X"8FC40020";
        ram_buffer(23449) := X"AFA70030";
        ram_buffer(23450) := X"8C900014";
        ram_buffer(23451) := X"AFA50024";
        ram_buffer(23452) := X"8E02000C";
        ram_buffer(23453) := X"00000000";
        ram_buffer(23454) := X"0040F809";
        ram_buffer(23455) := X"00000000";
        ram_buffer(23456) := X"8FA50024";
        ram_buffer(23457) := X"8FA70030";
        ram_buffer(23458) := X"1440000B";
        ram_buffer(23459) := X"24030016";
        ram_buffer(23460) := X"8FC40020";
        ram_buffer(23461) := X"00000000";
        ram_buffer(23462) := X"8C820000";
        ram_buffer(23463) := X"00000000";
        ram_buffer(23464) := X"8C490000";
        ram_buffer(23465) := X"00000000";
        ram_buffer(23466) := X"0120F809";
        ram_buffer(23467) := X"AC430014";
        ram_buffer(23468) := X"8FA70030";
        ram_buffer(23469) := X"8FA50024";
        ram_buffer(23470) := X"8E040000";
        ram_buffer(23471) := X"8E020004";
        ram_buffer(23472) := X"AFC40010";
        ram_buffer(23473) := X"1000FF97";
        ram_buffer(23474) := X"AFC20014";
        ram_buffer(23475) := X"8FC40020";
        ram_buffer(23476) := X"00000000";
        ram_buffer(23477) := X"8C930014";
        ram_buffer(23478) := X"00000000";
        ram_buffer(23479) := X"8E62000C";
        ram_buffer(23480) := X"00000000";
        ram_buffer(23481) := X"0040F809";
        ram_buffer(23482) := X"00000000";
        ram_buffer(23483) := X"14400009";
        ram_buffer(23484) := X"24030016";
        ram_buffer(23485) := X"8FC40020";
        ram_buffer(23486) := X"00000000";
        ram_buffer(23487) := X"8C820000";
        ram_buffer(23488) := X"00000000";
        ram_buffer(23489) := X"8C490000";
        ram_buffer(23490) := X"00000000";
        ram_buffer(23491) := X"0120F809";
        ram_buffer(23492) := X"AC430014";
        ram_buffer(23493) := X"8E640000";
        ram_buffer(23494) := X"8E620004";
        ram_buffer(23495) := X"AFC40010";
        ram_buffer(23496) := X"1611FFA3";
        ram_buffer(23497) := X"AFC20014";
        ram_buffer(23498) := X"8FC20010";
        ram_buffer(23499) := X"00000000";
        ram_buffer(23500) := X"24440001";
        ram_buffer(23501) := X"AFC40010";
        ram_buffer(23502) := X"A0400000";
        ram_buffer(23503) := X"8FC20014";
        ram_buffer(23504) := X"00000000";
        ram_buffer(23505) := X"2442FFFF";
        ram_buffer(23506) := X"1440FF99";
        ram_buffer(23507) := X"AFC20014";
        ram_buffer(23508) := X"8FC40020";
        ram_buffer(23509) := X"00000000";
        ram_buffer(23510) := X"8C900014";
        ram_buffer(23511) := X"00000000";
        ram_buffer(23512) := X"8E02000C";
        ram_buffer(23513) := X"00000000";
        ram_buffer(23514) := X"0040F809";
        ram_buffer(23515) := X"00000000";
        ram_buffer(23516) := X"10400019";
        ram_buffer(23517) := X"24030016";
        ram_buffer(23518) := X"8E040000";
        ram_buffer(23519) := X"8E020004";
        ram_buffer(23520) := X"AFC40010";
        ram_buffer(23521) := X"1000FF8A";
        ram_buffer(23522) := X"AFC20014";
        ram_buffer(23523) := X"0C024CF4";
        ram_buffer(23524) := X"03C02021";
        ram_buffer(23525) := X"1000FDA9";
        ram_buffer(23526) := X"00000000";
        ram_buffer(23527) := X"8FC40020";
        ram_buffer(23528) := X"24030027";
        ram_buffer(23529) := X"8C820000";
        ram_buffer(23530) := X"AFA70030";
        ram_buffer(23531) := X"8C480000";
        ram_buffer(23532) := X"AC430014";
        ram_buffer(23533) := X"0100F809";
        ram_buffer(23534) := X"AFA50024";
        ram_buffer(23535) := X"8FC2000C";
        ram_buffer(23536) := X"8FA50024";
        ram_buffer(23537) := X"8FA70030";
        ram_buffer(23538) := X"1440FF19";
        ram_buffer(23539) := X"24020001";
        ram_buffer(23540) := X"1000FF3C";
        ram_buffer(23541) := X"02421004";
        ram_buffer(23542) := X"8FC40020";
        ram_buffer(23543) := X"00000000";
        ram_buffer(23544) := X"8C820000";
        ram_buffer(23545) := X"00000000";
        ram_buffer(23546) := X"8C480000";
        ram_buffer(23547) := X"00000000";
        ram_buffer(23548) := X"0100F809";
        ram_buffer(23549) := X"AC430014";
        ram_buffer(23550) := X"1000FFDF";
        ram_buffer(23551) := X"00000000";
        ram_buffer(23552) := X"1000FEFD";
        ram_buffer(23553) := X"00002821";
        ram_buffer(23554) := X"8C820004";
        ram_buffer(23555) := X"27BDFFE0";
        ram_buffer(23556) := X"8C420000";
        ram_buffer(23557) := X"2406006C";
        ram_buffer(23558) := X"AFBF001C";
        ram_buffer(23559) := X"AFB10018";
        ram_buffer(23560) := X"AFB00014";
        ram_buffer(23561) := X"24050001";
        ram_buffer(23562) := X"0040F809";
        ram_buffer(23563) := X"00808821";
        ram_buffer(23564) := X"00408021";
        ram_buffer(23565) := X"AE220164";
        ram_buffer(23566) := X"3C021009";
        ram_buffer(23567) := X"24422944";
        ram_buffer(23568) := X"2604004C";
        ram_buffer(23569) := X"24060010";
        ram_buffer(23570) := X"AE020000";
        ram_buffer(23571) := X"0C02801D";
        ram_buffer(23572) := X"00002821";
        ram_buffer(23573) := X"2604005C";
        ram_buffer(23574) := X"24060010";
        ram_buffer(23575) := X"0C02801D";
        ram_buffer(23576) := X"00002821";
        ram_buffer(23577) := X"8FBF001C";
        ram_buffer(23578) := X"AE000040";
        ram_buffer(23579) := X"8FB10018";
        ram_buffer(23580) := X"8FB00014";
        ram_buffer(23581) := X"03E00008";
        ram_buffer(23582) := X"27BD0020";
        ram_buffer(23583) := X"8C830160";
        ram_buffer(23584) := X"27BDFF18";
        ram_buffer(23585) := X"8C820034";
        ram_buffer(23586) := X"AFA300B8";
        ram_buffer(23587) := X"8C83003C";
        ram_buffer(23588) := X"AFBF00E4";
        ram_buffer(23589) := X"AFBE00E0";
        ram_buffer(23590) := X"AFB700DC";
        ram_buffer(23591) := X"AFB600D8";
        ram_buffer(23592) := X"AFB500D4";
        ram_buffer(23593) := X"AFB400D0";
        ram_buffer(23594) := X"AFB300CC";
        ram_buffer(23595) := X"AFB200C8";
        ram_buffer(23596) := X"AFB100C4";
        ram_buffer(23597) := X"AFB000C0";
        ram_buffer(23598) := X"AFA30010";
        ram_buffer(23599) := X"18400140";
        ram_buffer(23600) := X"AFA000B4";
        ram_buffer(23601) := X"8F828028";
        ram_buffer(23602) := X"0080B821";
        ram_buffer(23603) := X"AFA20094";
        ram_buffer(23604) := X"00402021";
        ram_buffer(23605) := X"8F82802C";
        ram_buffer(23606) := X"8F838034";
        ram_buffer(23607) := X"00402821";
        ram_buffer(23608) := X"AFA200A8";
        ram_buffer(23609) := X"8F828030";
        ram_buffer(23610) := X"AFA3009C";
        ram_buffer(23611) := X"AFA20098";
        ram_buffer(23612) := X"8F828038";
        ram_buffer(23613) := X"8F83803C";
        ram_buffer(23614) := X"AFA200A0";
        ram_buffer(23615) := X"3C02100D";
        ram_buffer(23616) := X"3C08100D";
        ram_buffer(23617) := X"244288E8";
        ram_buffer(23618) := X"AFA300A4";
        ram_buffer(23619) := X"25168968";
        ram_buffer(23620) := X"AFA20090";
        ram_buffer(23621) := X"AFA400AC";
        ram_buffer(23622) := X"AFA500B0";
        ram_buffer(23623) := X"8FA20010";
        ram_buffer(23624) := X"00000000";
        ram_buffer(23625) := X"8C510010";
        ram_buffer(23626) := X"00000000";
        ram_buffer(23627) := X"2E220004";
        ram_buffer(23628) := X"1040012F";
        ram_buffer(23629) := X"26320010";
        ram_buffer(23630) := X"00121080";
        ram_buffer(23631) := X"02E21021";
        ram_buffer(23632) := X"8C500000";
        ram_buffer(23633) := X"00000000";
        ram_buffer(23634) := X"12000129";
        ram_buffer(23635) := X"24030001";
        ram_buffer(23636) := X"8EE200BC";
        ram_buffer(23637) := X"00000000";
        ram_buffer(23638) := X"10430135";
        ram_buffer(23639) := X"00000000";
        ram_buffer(23640) := X"10400151";
        ram_buffer(23641) := X"24030002";
        ram_buffer(23642) := X"14430147";
        ram_buffer(23643) := X"2404002F";
        ram_buffer(23644) := X"8FA200B8";
        ram_buffer(23645) := X"00118880";
        ram_buffer(23646) := X"00519021";
        ram_buffer(23647) := X"8E510020";
        ram_buffer(23648) := X"00000000";
        ram_buffer(23649) := X"12200169";
        ram_buffer(23650) := X"00000000";
        ram_buffer(23651) := X"8F828028";
        ram_buffer(23652) := X"8F838044";
        ram_buffer(23653) := X"00402021";
        ram_buffer(23654) := X"AFA20014";
        ram_buffer(23655) := X"8F82802C";
        ram_buffer(23656) := X"AFA3001C";
        ram_buffer(23657) := X"00402821";
        ram_buffer(23658) := X"AFA20040";
        ram_buffer(23659) := X"8F828040";
        ram_buffer(23660) := X"8F83804C";
        ram_buffer(23661) := X"AFA20018";
        ram_buffer(23662) := X"8F828048";
        ram_buffer(23663) := X"AFA30024";
        ram_buffer(23664) := X"AFA20020";
        ram_buffer(23665) := X"8F838054";
        ram_buffer(23666) := X"8F828050";
        ram_buffer(23667) := X"AFA3002C";
        ram_buffer(23668) := X"AFA20028";
        ram_buffer(23669) := X"8F83805C";
        ram_buffer(23670) := X"8F828058";
        ram_buffer(23671) := X"8F958030";
        ram_buffer(23672) := X"8F948034";
        ram_buffer(23673) := X"AFA30034";
        ram_buffer(23674) := X"AFA20030";
        ram_buffer(23675) := X"8F838064";
        ram_buffer(23676) := X"8F828060";
        ram_buffer(23677) := X"3C08100D";
        ram_buffer(23678) := X"251E88A8";
        ram_buffer(23679) := X"AFA3003C";
        ram_buffer(23680) := X"AFA20038";
        ram_buffer(23681) := X"AFB50044";
        ram_buffer(23682) := X"AFB40048";
        ram_buffer(23683) := X"AFA4004C";
        ram_buffer(23684) := X"AFA50050";
        ram_buffer(23685) := X"AFB50054";
        ram_buffer(23686) := X"AFB40058";
        ram_buffer(23687) := X"26100002";
        ram_buffer(23688) := X"AFA4005C";
        ram_buffer(23689) := X"AFB700BC";
        ram_buffer(23690) := X"AFA50060";
        ram_buffer(23691) := X"03C0B821";
        ram_buffer(23692) := X"AFB50064";
        ram_buffer(23693) := X"AFB40068";
        ram_buffer(23694) := X"AFA4006C";
        ram_buffer(23695) := X"AFA50070";
        ram_buffer(23696) := X"AFB50074";
        ram_buffer(23697) := X"AFB40078";
        ram_buffer(23698) := X"AFA4007C";
        ram_buffer(23699) := X"AFA50080";
        ram_buffer(23700) := X"AFB50084";
        ram_buffer(23701) := X"AFB40088";
        ram_buffer(23702) := X"AFA4008C";
        ram_buffer(23703) := X"00A0F021";
        ram_buffer(23704) := X"9604FFFE";
        ram_buffer(23705) := X"8EF30004";
        ram_buffer(23706) := X"8EF20000";
        ram_buffer(23707) := X"0C031BBD";
        ram_buffer(23708) := X"26F70008";
        ram_buffer(23709) := X"00602821";
        ram_buffer(23710) := X"02603821";
        ram_buffer(23711) := X"02403021";
        ram_buffer(23712) := X"0C03174A";
        ram_buffer(23713) := X"00402021";
        ram_buffer(23714) := X"8FA60094";
        ram_buffer(23715) := X"8FA700A8";
        ram_buffer(23716) := X"00602821";
        ram_buffer(23717) := X"0C03174A";
        ram_buffer(23718) := X"00402021";
        ram_buffer(23719) := X"8FA5009C";
        ram_buffer(23720) := X"8FA40098";
        ram_buffer(23721) := X"00603821";
        ram_buffer(23722) := X"0C03144F";
        ram_buffer(23723) := X"00403021";
        ram_buffer(23724) := X"00602821";
        ram_buffer(23725) := X"0C031C96";
        ram_buffer(23726) := X"00402021";
        ram_buffer(23727) := X"96040000";
        ram_buffer(23728) := X"0C031BBD";
        ram_buffer(23729) := X"AE220000";
        ram_buffer(23730) := X"00602821";
        ram_buffer(23731) := X"02603821";
        ram_buffer(23732) := X"02403021";
        ram_buffer(23733) := X"0C03174A";
        ram_buffer(23734) := X"00402021";
        ram_buffer(23735) := X"8FA700A4";
        ram_buffer(23736) := X"8FA600A0";
        ram_buffer(23737) := X"00602821";
        ram_buffer(23738) := X"0C03174A";
        ram_buffer(23739) := X"00402021";
        ram_buffer(23740) := X"8FA600AC";
        ram_buffer(23741) := X"8FA700B0";
        ram_buffer(23742) := X"00602821";
        ram_buffer(23743) := X"0C03174A";
        ram_buffer(23744) := X"00402021";
        ram_buffer(23745) := X"00603821";
        ram_buffer(23746) := X"00403021";
        ram_buffer(23747) := X"02A02021";
        ram_buffer(23748) := X"0C03144F";
        ram_buffer(23749) := X"02802821";
        ram_buffer(23750) := X"00602821";
        ram_buffer(23751) := X"0C031C96";
        ram_buffer(23752) := X"00402021";
        ram_buffer(23753) := X"96040002";
        ram_buffer(23754) := X"0C031BBD";
        ram_buffer(23755) := X"AE220004";
        ram_buffer(23756) := X"00602821";
        ram_buffer(23757) := X"02603821";
        ram_buffer(23758) := X"02403021";
        ram_buffer(23759) := X"0C03174A";
        ram_buffer(23760) := X"00402021";
        ram_buffer(23761) := X"8FA7001C";
        ram_buffer(23762) := X"8FA60018";
        ram_buffer(23763) := X"00602821";
        ram_buffer(23764) := X"0C03174A";
        ram_buffer(23765) := X"00402021";
        ram_buffer(23766) := X"8FA60014";
        ram_buffer(23767) := X"8FA70040";
        ram_buffer(23768) := X"00602821";
        ram_buffer(23769) := X"0C03174A";
        ram_buffer(23770) := X"00402021";
        ram_buffer(23771) := X"8FA40044";
        ram_buffer(23772) := X"8FA50048";
        ram_buffer(23773) := X"00603821";
        ram_buffer(23774) := X"0C03144F";
        ram_buffer(23775) := X"00403021";
        ram_buffer(23776) := X"00602821";
        ram_buffer(23777) := X"0C031C96";
        ram_buffer(23778) := X"00402021";
        ram_buffer(23779) := X"96040004";
        ram_buffer(23780) := X"0C031BBD";
        ram_buffer(23781) := X"AE220008";
        ram_buffer(23782) := X"00602821";
        ram_buffer(23783) := X"02603821";
        ram_buffer(23784) := X"02403021";
        ram_buffer(23785) := X"0C03174A";
        ram_buffer(23786) := X"00402021";
        ram_buffer(23787) := X"8FA70024";
        ram_buffer(23788) := X"8FA60020";
        ram_buffer(23789) := X"00602821";
        ram_buffer(23790) := X"0C03174A";
        ram_buffer(23791) := X"00402021";
        ram_buffer(23792) := X"8FA6004C";
        ram_buffer(23793) := X"8FA70050";
        ram_buffer(23794) := X"00602821";
        ram_buffer(23795) := X"0C03174A";
        ram_buffer(23796) := X"00402021";
        ram_buffer(23797) := X"8FA40054";
        ram_buffer(23798) := X"8FA50058";
        ram_buffer(23799) := X"00603821";
        ram_buffer(23800) := X"0C03144F";
        ram_buffer(23801) := X"00403021";
        ram_buffer(23802) := X"00602821";
        ram_buffer(23803) := X"0C031C96";
        ram_buffer(23804) := X"00402021";
        ram_buffer(23805) := X"96040006";
        ram_buffer(23806) := X"0C031BBD";
        ram_buffer(23807) := X"AE22000C";
        ram_buffer(23808) := X"00602821";
        ram_buffer(23809) := X"02603821";
        ram_buffer(23810) := X"02403021";
        ram_buffer(23811) := X"0C03174A";
        ram_buffer(23812) := X"00402021";
        ram_buffer(23813) := X"8FA6005C";
        ram_buffer(23814) := X"8FA70060";
        ram_buffer(23815) := X"00602821";
        ram_buffer(23816) := X"0C03174A";
        ram_buffer(23817) := X"00402021";
        ram_buffer(23818) := X"8FA40064";
        ram_buffer(23819) := X"8FA50068";
        ram_buffer(23820) := X"00603821";
        ram_buffer(23821) := X"0C03144F";
        ram_buffer(23822) := X"00403021";
        ram_buffer(23823) := X"00602821";
        ram_buffer(23824) := X"0C031C96";
        ram_buffer(23825) := X"00402021";
        ram_buffer(23826) := X"96040008";
        ram_buffer(23827) := X"0C031BBD";
        ram_buffer(23828) := X"AE220010";
        ram_buffer(23829) := X"00602821";
        ram_buffer(23830) := X"02603821";
        ram_buffer(23831) := X"02403021";
        ram_buffer(23832) := X"0C03174A";
        ram_buffer(23833) := X"00402021";
        ram_buffer(23834) := X"8FA7002C";
        ram_buffer(23835) := X"8FA60028";
        ram_buffer(23836) := X"00602821";
        ram_buffer(23837) := X"0C03174A";
        ram_buffer(23838) := X"00402021";
        ram_buffer(23839) := X"8FA6006C";
        ram_buffer(23840) := X"8FA70070";
        ram_buffer(23841) := X"00602821";
        ram_buffer(23842) := X"0C03174A";
        ram_buffer(23843) := X"00402021";
        ram_buffer(23844) := X"8FA40074";
        ram_buffer(23845) := X"8FA50078";
        ram_buffer(23846) := X"00603821";
        ram_buffer(23847) := X"0C03144F";
        ram_buffer(23848) := X"00403021";
        ram_buffer(23849) := X"00602821";
        ram_buffer(23850) := X"0C031C96";
        ram_buffer(23851) := X"00402021";
        ram_buffer(23852) := X"9604000A";
        ram_buffer(23853) := X"0C031BBD";
        ram_buffer(23854) := X"AE220014";
        ram_buffer(23855) := X"00602821";
        ram_buffer(23856) := X"02603821";
        ram_buffer(23857) := X"02403021";
        ram_buffer(23858) := X"0C03174A";
        ram_buffer(23859) := X"00402021";
        ram_buffer(23860) := X"8FA70034";
        ram_buffer(23861) := X"8FA60030";
        ram_buffer(23862) := X"00602821";
        ram_buffer(23863) := X"0C03174A";
        ram_buffer(23864) := X"00402021";
        ram_buffer(23865) := X"8FA6007C";
        ram_buffer(23866) := X"8FA70080";
        ram_buffer(23867) := X"00602821";
        ram_buffer(23868) := X"0C03174A";
        ram_buffer(23869) := X"00402021";
        ram_buffer(23870) := X"8FA40084";
        ram_buffer(23871) := X"8FA50088";
        ram_buffer(23872) := X"00603821";
        ram_buffer(23873) := X"0C03144F";
        ram_buffer(23874) := X"00403021";
        ram_buffer(23875) := X"00602821";
        ram_buffer(23876) := X"0C031C96";
        ram_buffer(23877) := X"00402021";
        ram_buffer(23878) := X"9604000C";
        ram_buffer(23879) := X"0C031BBD";
        ram_buffer(23880) := X"AE220018";
        ram_buffer(23881) := X"00602821";
        ram_buffer(23882) := X"02603821";
        ram_buffer(23883) := X"02403021";
        ram_buffer(23884) := X"0C03174A";
        ram_buffer(23885) := X"00402021";
        ram_buffer(23886) := X"8FA7003C";
        ram_buffer(23887) := X"8FA60038";
        ram_buffer(23888) := X"00602821";
        ram_buffer(23889) := X"0C03174A";
        ram_buffer(23890) := X"00402021";
        ram_buffer(23891) := X"8FA6008C";
        ram_buffer(23892) := X"03C03821";
        ram_buffer(23893) := X"00602821";
        ram_buffer(23894) := X"0C03174A";
        ram_buffer(23895) := X"00402021";
        ram_buffer(23896) := X"00603821";
        ram_buffer(23897) := X"00403021";
        ram_buffer(23898) := X"02A02021";
        ram_buffer(23899) := X"0C03144F";
        ram_buffer(23900) := X"02802821";
        ram_buffer(23901) := X"00602821";
        ram_buffer(23902) := X"0C031C96";
        ram_buffer(23903) := X"00402021";
        ram_buffer(23904) := X"AE22001C";
        ram_buffer(23905) := X"8FA20090";
        ram_buffer(23906) := X"26100010";
        ram_buffer(23907) := X"16E2FF34";
        ram_buffer(23908) := X"26310020";
        ram_buffer(23909) := X"8FB700BC";
        ram_buffer(23910) := X"8FA300B4";
        ram_buffer(23911) := X"8EE20034";
        ram_buffer(23912) := X"24630001";
        ram_buffer(23913) := X"AFA300B4";
        ram_buffer(23914) := X"0062102A";
        ram_buffer(23915) := X"8FA30010";
        ram_buffer(23916) := X"00000000";
        ram_buffer(23917) := X"24630054";
        ram_buffer(23918) := X"1440FED8";
        ram_buffer(23919) := X"AFA30010";
        ram_buffer(23920) := X"8FBF00E4";
        ram_buffer(23921) := X"8FBE00E0";
        ram_buffer(23922) := X"8FB700DC";
        ram_buffer(23923) := X"8FB600D8";
        ram_buffer(23924) := X"8FB500D4";
        ram_buffer(23925) := X"8FB400D0";
        ram_buffer(23926) := X"8FB300CC";
        ram_buffer(23927) := X"8FB200C8";
        ram_buffer(23928) := X"8FB100C4";
        ram_buffer(23929) := X"8FB000C0";
        ram_buffer(23930) := X"03E00008";
        ram_buffer(23931) := X"27BD00E8";
        ram_buffer(23932) := X"8EE20000";
        ram_buffer(23933) := X"24040033";
        ram_buffer(23934) := X"AC510018";
        ram_buffer(23935) := X"8EE30000";
        ram_buffer(23936) := X"AC440014";
        ram_buffer(23937) := X"8C620000";
        ram_buffer(23938) := X"00000000";
        ram_buffer(23939) := X"0040F809";
        ram_buffer(23940) := X"02E02021";
        ram_buffer(23941) := X"00129080";
        ram_buffer(23942) := X"8EE200BC";
        ram_buffer(23943) := X"02F29021";
        ram_buffer(23944) := X"24030001";
        ram_buffer(23945) := X"8E500000";
        ram_buffer(23946) := X"1443FECD";
        ram_buffer(23947) := X"00000000";
        ram_buffer(23948) := X"8FA200B8";
        ram_buffer(23949) := X"00118880";
        ram_buffer(23950) := X"00518821";
        ram_buffer(23951) := X"8E25000C";
        ram_buffer(23952) := X"00000000";
        ram_buffer(23953) := X"10A00028";
        ram_buffer(23954) := X"24060100";
        ram_buffer(23955) := X"3C04100D";
        ram_buffer(23956) := X"248488E8";
        ram_buffer(23957) := X"96020000";
        ram_buffer(23958) := X"84830000";
        ram_buffer(23959) := X"24A50004";
        ram_buffer(23960) := X"00430018";
        ram_buffer(23961) := X"24840002";
        ram_buffer(23962) := X"26100002";
        ram_buffer(23963) := X"00001012";
        ram_buffer(23964) := X"24420400";
        ram_buffer(23965) := X"000212C3";
        ram_buffer(23966) := X"16C4FFF6";
        ram_buffer(23967) := X"ACA2FFFC";
        ram_buffer(23968) := X"1000FFC5";
        ram_buffer(23969) := X"00000000";
        ram_buffer(23970) := X"8EE20000";
        ram_buffer(23971) := X"00000000";
        ram_buffer(23972) := X"8C430000";
        ram_buffer(23973) := X"AC440014";
        ram_buffer(23974) := X"0060F809";
        ram_buffer(23975) := X"02E02021";
        ram_buffer(23976) := X"1000FFBD";
        ram_buffer(23977) := X"00000000";
        ram_buffer(23978) := X"8FA200B8";
        ram_buffer(23979) := X"00118880";
        ram_buffer(23980) := X"00518821";
        ram_buffer(23981) := X"8E22000C";
        ram_buffer(23982) := X"00000000";
        ram_buffer(23983) := X"10400013";
        ram_buffer(23984) := X"24060100";
        ram_buffer(23985) := X"24440100";
        ram_buffer(23986) := X"96030000";
        ram_buffer(23987) := X"24420004";
        ram_buffer(23988) := X"000318C0";
        ram_buffer(23989) := X"AC43FFFC";
        ram_buffer(23990) := X"1482FFFB";
        ram_buffer(23991) := X"26100002";
        ram_buffer(23992) := X"1000FFAD";
        ram_buffer(23993) := X"00000000";
        ram_buffer(23994) := X"8EE20004";
        ram_buffer(23995) := X"24050001";
        ram_buffer(23996) := X"8C420000";
        ram_buffer(23997) := X"00000000";
        ram_buffer(23998) := X"0040F809";
        ram_buffer(23999) := X"02E02021";
        ram_buffer(24000) := X"AE22000C";
        ram_buffer(24001) := X"1000FFD1";
        ram_buffer(24002) := X"00402821";
        ram_buffer(24003) := X"8EE20004";
        ram_buffer(24004) := X"00000000";
        ram_buffer(24005) := X"8C420000";
        ram_buffer(24006) := X"24050001";
        ram_buffer(24007) := X"0040F809";
        ram_buffer(24008) := X"02E02021";
        ram_buffer(24009) := X"1000FFE7";
        ram_buffer(24010) := X"AE22000C";
        ram_buffer(24011) := X"8EE20004";
        ram_buffer(24012) := X"24060100";
        ram_buffer(24013) := X"8C420000";
        ram_buffer(24014) := X"24050001";
        ram_buffer(24015) := X"0040F809";
        ram_buffer(24016) := X"02E02021";
        ram_buffer(24017) := X"AE420020";
        ram_buffer(24018) := X"1000FE90";
        ram_buffer(24019) := X"00408821";
        ram_buffer(24020) := X"8CA20010";
        ram_buffer(24021) := X"8C830160";
        ram_buffer(24022) := X"24420002";
        ram_buffer(24023) := X"00021080";
        ram_buffer(24024) := X"00621021";
        ram_buffer(24025) := X"8C420004";
        ram_buffer(24026) := X"27BDFEB0";
        ram_buffer(24027) := X"8C630008";
        ram_buffer(24028) := X"AFA20120";
        ram_buffer(24029) := X"8FA20168";
        ram_buffer(24030) := X"AFBE0148";
        ram_buffer(24031) := X"AFB40138";
        ram_buffer(24032) := X"AFBF014C";
        ram_buffer(24033) := X"AFB70144";
        ram_buffer(24034) := X"AFB60140";
        ram_buffer(24035) := X"AFB5013C";
        ram_buffer(24036) := X"AFB30134";
        ram_buffer(24037) := X"AFB20130";
        ram_buffer(24038) := X"AFB1012C";
        ram_buffer(24039) := X"AFB00128";
        ram_buffer(24040) := X"8FB40164";
        ram_buffer(24041) := X"AFA3011C";
        ram_buffer(24042) := X"8FBE0160";
        ram_buffer(24043) := X"10400140";
        ram_buffer(24044) := X"001EF080";
        ram_buffer(24045) := X"27CC0004";
        ram_buffer(24046) := X"27CB0008";
        ram_buffer(24047) := X"27CA000C";
        ram_buffer(24048) := X"27C90010";
        ram_buffer(24049) := X"27C80014";
        ram_buffer(24050) := X"27D7001C";
        ram_buffer(24051) := X"00E0A821";
        ram_buffer(24052) := X"27C70018";
        ram_buffer(24053) := X"00CC6021";
        ram_buffer(24054) := X"00DEF021";
        ram_buffer(24055) := X"00CB5821";
        ram_buffer(24056) := X"00CA5021";
        ram_buffer(24057) := X"00C99021";
        ram_buffer(24058) := X"00C88821";
        ram_buffer(24059) := X"00C78021";
        ram_buffer(24060) := X"00D7B821";
        ram_buffer(24061) := X"0000B021";
        ram_buffer(24062) := X"27B30110";
        ram_buffer(24063) := X"8FC30000";
        ram_buffer(24064) := X"8D820000";
        ram_buffer(24065) := X"00741821";
        ram_buffer(24066) := X"90640000";
        ram_buffer(24067) := X"00541021";
        ram_buffer(24068) := X"2484FF80";
        ram_buffer(24069) := X"AFA40010";
        ram_buffer(24070) := X"90650001";
        ram_buffer(24071) := X"AFAC0118";
        ram_buffer(24072) := X"24A5FF80";
        ram_buffer(24073) := X"AFA50014";
        ram_buffer(24074) := X"90650002";
        ram_buffer(24075) := X"00000000";
        ram_buffer(24076) := X"24A5FF80";
        ram_buffer(24077) := X"AFA50018";
        ram_buffer(24078) := X"90650003";
        ram_buffer(24079) := X"00000000";
        ram_buffer(24080) := X"24A5FF80";
        ram_buffer(24081) := X"AFA5001C";
        ram_buffer(24082) := X"90650004";
        ram_buffer(24083) := X"00000000";
        ram_buffer(24084) := X"24A5FF80";
        ram_buffer(24085) := X"AFA50020";
        ram_buffer(24086) := X"90650005";
        ram_buffer(24087) := X"00000000";
        ram_buffer(24088) := X"24A5FF80";
        ram_buffer(24089) := X"AFA50024";
        ram_buffer(24090) := X"90650006";
        ram_buffer(24091) := X"00000000";
        ram_buffer(24092) := X"24A5FF80";
        ram_buffer(24093) := X"AFA50028";
        ram_buffer(24094) := X"90630007";
        ram_buffer(24095) := X"00000000";
        ram_buffer(24096) := X"2463FF80";
        ram_buffer(24097) := X"AFA3002C";
        ram_buffer(24098) := X"90430000";
        ram_buffer(24099) := X"00000000";
        ram_buffer(24100) := X"2463FF80";
        ram_buffer(24101) := X"AFA30030";
        ram_buffer(24102) := X"90430001";
        ram_buffer(24103) := X"00000000";
        ram_buffer(24104) := X"2463FF80";
        ram_buffer(24105) := X"AFA30034";
        ram_buffer(24106) := X"90430002";
        ram_buffer(24107) := X"00000000";
        ram_buffer(24108) := X"2463FF80";
        ram_buffer(24109) := X"AFA30038";
        ram_buffer(24110) := X"90430003";
        ram_buffer(24111) := X"00000000";
        ram_buffer(24112) := X"2463FF80";
        ram_buffer(24113) := X"AFA3003C";
        ram_buffer(24114) := X"90430004";
        ram_buffer(24115) := X"00000000";
        ram_buffer(24116) := X"2463FF80";
        ram_buffer(24117) := X"AFA30040";
        ram_buffer(24118) := X"90430005";
        ram_buffer(24119) := X"00000000";
        ram_buffer(24120) := X"2463FF80";
        ram_buffer(24121) := X"AFA30044";
        ram_buffer(24122) := X"90430006";
        ram_buffer(24123) := X"00000000";
        ram_buffer(24124) := X"2463FF80";
        ram_buffer(24125) := X"AFA30048";
        ram_buffer(24126) := X"90420007";
        ram_buffer(24127) := X"8D630000";
        ram_buffer(24128) := X"2442FF80";
        ram_buffer(24129) := X"AFA2004C";
        ram_buffer(24130) := X"00741821";
        ram_buffer(24131) := X"90650000";
        ram_buffer(24132) := X"8D420000";
        ram_buffer(24133) := X"24A5FF80";
        ram_buffer(24134) := X"AFA50050";
        ram_buffer(24135) := X"90650001";
        ram_buffer(24136) := X"00541021";
        ram_buffer(24137) := X"24A5FF80";
        ram_buffer(24138) := X"AFA50054";
        ram_buffer(24139) := X"90650002";
        ram_buffer(24140) := X"AFAB0114";
        ram_buffer(24141) := X"24A5FF80";
        ram_buffer(24142) := X"AFA50058";
        ram_buffer(24143) := X"90650003";
        ram_buffer(24144) := X"AFAA0110";
        ram_buffer(24145) := X"24A5FF80";
        ram_buffer(24146) := X"AFA5005C";
        ram_buffer(24147) := X"90650004";
        ram_buffer(24148) := X"00000000";
        ram_buffer(24149) := X"24A5FF80";
        ram_buffer(24150) := X"AFA50060";
        ram_buffer(24151) := X"90650005";
        ram_buffer(24152) := X"00000000";
        ram_buffer(24153) := X"24A5FF80";
        ram_buffer(24154) := X"AFA50064";
        ram_buffer(24155) := X"90650006";
        ram_buffer(24156) := X"00000000";
        ram_buffer(24157) := X"24A5FF80";
        ram_buffer(24158) := X"AFA50068";
        ram_buffer(24159) := X"90630007";
        ram_buffer(24160) := X"00000000";
        ram_buffer(24161) := X"2463FF80";
        ram_buffer(24162) := X"AFA3006C";
        ram_buffer(24163) := X"90430000";
        ram_buffer(24164) := X"00000000";
        ram_buffer(24165) := X"2463FF80";
        ram_buffer(24166) := X"AFA30070";
        ram_buffer(24167) := X"90430001";
        ram_buffer(24168) := X"00000000";
        ram_buffer(24169) := X"2463FF80";
        ram_buffer(24170) := X"AFA30074";
        ram_buffer(24171) := X"90430002";
        ram_buffer(24172) := X"00000000";
        ram_buffer(24173) := X"2463FF80";
        ram_buffer(24174) := X"AFA30078";
        ram_buffer(24175) := X"90430003";
        ram_buffer(24176) := X"00000000";
        ram_buffer(24177) := X"2463FF80";
        ram_buffer(24178) := X"AFA3007C";
        ram_buffer(24179) := X"90430004";
        ram_buffer(24180) := X"00000000";
        ram_buffer(24181) := X"2463FF80";
        ram_buffer(24182) := X"AFA30080";
        ram_buffer(24183) := X"90430005";
        ram_buffer(24184) := X"00000000";
        ram_buffer(24185) := X"2463FF80";
        ram_buffer(24186) := X"AFA30084";
        ram_buffer(24187) := X"90450006";
        ram_buffer(24188) := X"8E430000";
        ram_buffer(24189) := X"24A5FF80";
        ram_buffer(24190) := X"AFA50088";
        ram_buffer(24191) := X"90420007";
        ram_buffer(24192) := X"00741821";
        ram_buffer(24193) := X"2442FF80";
        ram_buffer(24194) := X"AFA2008C";
        ram_buffer(24195) := X"90650000";
        ram_buffer(24196) := X"8E220000";
        ram_buffer(24197) := X"24A5FF80";
        ram_buffer(24198) := X"AFA50090";
        ram_buffer(24199) := X"90650001";
        ram_buffer(24200) := X"00541021";
        ram_buffer(24201) := X"24A5FF80";
        ram_buffer(24202) := X"AFA50094";
        ram_buffer(24203) := X"90650002";
        ram_buffer(24204) := X"00000000";
        ram_buffer(24205) := X"24A5FF80";
        ram_buffer(24206) := X"AFA50098";
        ram_buffer(24207) := X"90650003";
        ram_buffer(24208) := X"00000000";
        ram_buffer(24209) := X"24A5FF80";
        ram_buffer(24210) := X"AFA5009C";
        ram_buffer(24211) := X"90650004";
        ram_buffer(24212) := X"00000000";
        ram_buffer(24213) := X"24A5FF80";
        ram_buffer(24214) := X"AFA500A0";
        ram_buffer(24215) := X"90650005";
        ram_buffer(24216) := X"00000000";
        ram_buffer(24217) := X"24A5FF80";
        ram_buffer(24218) := X"AFA500A4";
        ram_buffer(24219) := X"90650006";
        ram_buffer(24220) := X"00000000";
        ram_buffer(24221) := X"24A5FF80";
        ram_buffer(24222) := X"AFA500A8";
        ram_buffer(24223) := X"90630007";
        ram_buffer(24224) := X"00000000";
        ram_buffer(24225) := X"2463FF80";
        ram_buffer(24226) := X"AFA300AC";
        ram_buffer(24227) := X"90430000";
        ram_buffer(24228) := X"00000000";
        ram_buffer(24229) := X"2463FF80";
        ram_buffer(24230) := X"AFA300B0";
        ram_buffer(24231) := X"90430001";
        ram_buffer(24232) := X"00000000";
        ram_buffer(24233) := X"2463FF80";
        ram_buffer(24234) := X"AFA300B4";
        ram_buffer(24235) := X"90430002";
        ram_buffer(24236) := X"00000000";
        ram_buffer(24237) := X"2463FF80";
        ram_buffer(24238) := X"AFA300B8";
        ram_buffer(24239) := X"90430003";
        ram_buffer(24240) := X"00000000";
        ram_buffer(24241) := X"2463FF80";
        ram_buffer(24242) := X"AFA300BC";
        ram_buffer(24243) := X"90430004";
        ram_buffer(24244) := X"00000000";
        ram_buffer(24245) := X"2463FF80";
        ram_buffer(24246) := X"AFA300C0";
        ram_buffer(24247) := X"90450005";
        ram_buffer(24248) := X"8E030000";
        ram_buffer(24249) := X"24A5FF80";
        ram_buffer(24250) := X"AFA500C4";
        ram_buffer(24251) := X"90450006";
        ram_buffer(24252) := X"00741821";
        ram_buffer(24253) := X"24A5FF80";
        ram_buffer(24254) := X"AFA500C8";
        ram_buffer(24255) := X"90450007";
        ram_buffer(24256) := X"8EE20000";
        ram_buffer(24257) := X"24A5FF80";
        ram_buffer(24258) := X"AFA500CC";
        ram_buffer(24259) := X"90650000";
        ram_buffer(24260) := X"00541021";
        ram_buffer(24261) := X"24A5FF80";
        ram_buffer(24262) := X"AFA500D0";
        ram_buffer(24263) := X"90650001";
        ram_buffer(24264) := X"00000000";
        ram_buffer(24265) := X"24A5FF80";
        ram_buffer(24266) := X"AFA500D4";
        ram_buffer(24267) := X"90650002";
        ram_buffer(24268) := X"00000000";
        ram_buffer(24269) := X"24A5FF80";
        ram_buffer(24270) := X"AFA500D8";
        ram_buffer(24271) := X"90650003";
        ram_buffer(24272) := X"00000000";
        ram_buffer(24273) := X"24A5FF80";
        ram_buffer(24274) := X"AFA500DC";
        ram_buffer(24275) := X"90650004";
        ram_buffer(24276) := X"00000000";
        ram_buffer(24277) := X"24A5FF80";
        ram_buffer(24278) := X"AFA500E0";
        ram_buffer(24279) := X"90650005";
        ram_buffer(24280) := X"00000000";
        ram_buffer(24281) := X"24A5FF80";
        ram_buffer(24282) := X"AFA500E4";
        ram_buffer(24283) := X"90650006";
        ram_buffer(24284) := X"00000000";
        ram_buffer(24285) := X"24A5FF80";
        ram_buffer(24286) := X"AFA500E8";
        ram_buffer(24287) := X"90630007";
        ram_buffer(24288) := X"00000000";
        ram_buffer(24289) := X"2463FF80";
        ram_buffer(24290) := X"AFA300EC";
        ram_buffer(24291) := X"90430000";
        ram_buffer(24292) := X"00000000";
        ram_buffer(24293) := X"2463FF80";
        ram_buffer(24294) := X"AFA300F0";
        ram_buffer(24295) := X"90430001";
        ram_buffer(24296) := X"00000000";
        ram_buffer(24297) := X"2463FF80";
        ram_buffer(24298) := X"AFA300F4";
        ram_buffer(24299) := X"90430002";
        ram_buffer(24300) := X"00000000";
        ram_buffer(24301) := X"2463FF80";
        ram_buffer(24302) := X"AFA300F8";
        ram_buffer(24303) := X"90430003";
        ram_buffer(24304) := X"00000000";
        ram_buffer(24305) := X"2463FF80";
        ram_buffer(24306) := X"AFA300FC";
        ram_buffer(24307) := X"90430004";
        ram_buffer(24308) := X"00000000";
        ram_buffer(24309) := X"2463FF80";
        ram_buffer(24310) := X"AFA30100";
        ram_buffer(24311) := X"90430005";
        ram_buffer(24312) := X"00000000";
        ram_buffer(24313) := X"2463FF80";
        ram_buffer(24314) := X"AFA30104";
        ram_buffer(24315) := X"90430006";
        ram_buffer(24316) := X"00000000";
        ram_buffer(24317) := X"2463FF80";
        ram_buffer(24318) := X"AFA30108";
        ram_buffer(24319) := X"90420007";
        ram_buffer(24320) := X"00000000";
        ram_buffer(24321) := X"2442FF80";
        ram_buffer(24322) := X"AFA2010C";
        ram_buffer(24323) := X"8FA2011C";
        ram_buffer(24324) := X"00000000";
        ram_buffer(24325) := X"0040F809";
        ram_buffer(24326) := X"27A40010";
        ram_buffer(24327) := X"8FAD0120";
        ram_buffer(24328) := X"27A50010";
        ram_buffer(24329) := X"8FAA0110";
        ram_buffer(24330) := X"8FAB0114";
        ram_buffer(24331) := X"8FAC0118";
        ram_buffer(24332) := X"1000000C";
        ram_buffer(24333) := X"02A03021";
        ram_buffer(24334) := X"15C00002";
        ram_buffer(24335) := X"004E001A";
        ram_buffer(24336) := X"0007000D";
        ram_buffer(24337) := X"00001012";
        ram_buffer(24338) := X"00021400";
        ram_buffer(24339) := X"00021403";
        ram_buffer(24340) := X"24A50004";
        ram_buffer(24341) := X"A4C20000";
        ram_buffer(24342) := X"25AD0004";
        ram_buffer(24343) := X"1265000F";
        ram_buffer(24344) := X"24C60002";
        ram_buffer(24345) := X"8CA20000";
        ram_buffer(24346) := X"8DAE0000";
        ram_buffer(24347) := X"0440001C";
        ram_buffer(24348) := X"000E1843";
        ram_buffer(24349) := X"00621021";
        ram_buffer(24350) := X"004E182A";
        ram_buffer(24351) := X"1060FFEE";
        ram_buffer(24352) := X"00000000";
        ram_buffer(24353) := X"00001021";
        ram_buffer(24354) := X"24A50004";
        ram_buffer(24355) := X"A4C20000";
        ram_buffer(24356) := X"25AD0004";
        ram_buffer(24357) := X"1665FFF3";
        ram_buffer(24358) := X"24C60002";
        ram_buffer(24359) := X"8FA20168";
        ram_buffer(24360) := X"26D60001";
        ram_buffer(24361) := X"26940008";
        ram_buffer(24362) := X"1456FED4";
        ram_buffer(24363) := X"26B50080";
        ram_buffer(24364) := X"8FBF014C";
        ram_buffer(24365) := X"8FBE0148";
        ram_buffer(24366) := X"8FB70144";
        ram_buffer(24367) := X"8FB60140";
        ram_buffer(24368) := X"8FB5013C";
        ram_buffer(24369) := X"8FB40138";
        ram_buffer(24370) := X"8FB30134";
        ram_buffer(24371) := X"8FB20130";
        ram_buffer(24372) := X"8FB1012C";
        ram_buffer(24373) := X"8FB00128";
        ram_buffer(24374) := X"03E00008";
        ram_buffer(24375) := X"27BD0150";
        ram_buffer(24376) := X"000E2043";
        ram_buffer(24377) := X"00821823";
        ram_buffer(24378) := X"006E102A";
        ram_buffer(24379) := X"1440FFE5";
        ram_buffer(24380) := X"00000000";
        ram_buffer(24381) := X"15C00002";
        ram_buffer(24382) := X"006E001A";
        ram_buffer(24383) := X"0007000D";
        ram_buffer(24384) := X"00001012";
        ram_buffer(24385) := X"00021023";
        ram_buffer(24386) := X"00021400";
        ram_buffer(24387) := X"1000FFD0";
        ram_buffer(24388) := X"00021403";
        ram_buffer(24389) := X"8CA20010";
        ram_buffer(24390) := X"8C830160";
        ram_buffer(24391) := X"24420008";
        ram_buffer(24392) := X"00021080";
        ram_buffer(24393) := X"00621021";
        ram_buffer(24394) := X"8C420000";
        ram_buffer(24395) := X"27BDFEA0";
        ram_buffer(24396) := X"8C63001C";
        ram_buffer(24397) := X"AFA20114";
        ram_buffer(24398) := X"8FA20178";
        ram_buffer(24399) := X"AFB60150";
        ram_buffer(24400) := X"AFB30144";
        ram_buffer(24401) := X"AFBF015C";
        ram_buffer(24402) := X"AFBE0158";
        ram_buffer(24403) := X"AFB70154";
        ram_buffer(24404) := X"AFB5014C";
        ram_buffer(24405) := X"AFB40148";
        ram_buffer(24406) := X"AFB20140";
        ram_buffer(24407) := X"AFB1013C";
        ram_buffer(24408) := X"AFB00138";
        ram_buffer(24409) := X"8FB30174";
        ram_buffer(24410) := X"AFA30110";
        ram_buffer(24411) := X"8FB60170";
        ram_buffer(24412) := X"10400155";
        ram_buffer(24413) := X"0016B080";
        ram_buffer(24414) := X"00C01021";
        ram_buffer(24415) := X"00564821";
        ram_buffer(24416) := X"26DE0004";
        ram_buffer(24417) := X"26D70008";
        ram_buffer(24418) := X"26C8000C";
        ram_buffer(24419) := X"26C60010";
        ram_buffer(24420) := X"26C50014";
        ram_buffer(24421) := X"26C40018";
        ram_buffer(24422) := X"26C3001C";
        ram_buffer(24423) := X"00484021";
        ram_buffer(24424) := X"00463021";
        ram_buffer(24425) := X"00452821";
        ram_buffer(24426) := X"00442021";
        ram_buffer(24427) := X"AFA90118";
        ram_buffer(24428) := X"005EF021";
        ram_buffer(24429) := X"00574821";
        ram_buffer(24430) := X"8F908068";
        ram_buffer(24431) := X"00431021";
        ram_buffer(24432) := X"AFA9011C";
        ram_buffer(24433) := X"AFA80120";
        ram_buffer(24434) := X"AFA60124";
        ram_buffer(24435) := X"AFA50128";
        ram_buffer(24436) := X"AFA4012C";
        ram_buffer(24437) := X"AFA20130";
        ram_buffer(24438) := X"00E0A021";
        ram_buffer(24439) := X"0000A821";
        ram_buffer(24440) := X"27B10110";
        ram_buffer(24441) := X"8FA20118";
        ram_buffer(24442) := X"0280B021";
        ram_buffer(24443) := X"8C520000";
        ram_buffer(24444) := X"00000000";
        ram_buffer(24445) := X"02539021";
        ram_buffer(24446) := X"92440000";
        ram_buffer(24447) := X"0C031190";
        ram_buffer(24448) := X"2484FF80";
        ram_buffer(24449) := X"AFA20010";
        ram_buffer(24450) := X"92440001";
        ram_buffer(24451) := X"0C031190";
        ram_buffer(24452) := X"2484FF80";
        ram_buffer(24453) := X"AFA20014";
        ram_buffer(24454) := X"92440002";
        ram_buffer(24455) := X"0C031190";
        ram_buffer(24456) := X"2484FF80";
        ram_buffer(24457) := X"AFA20018";
        ram_buffer(24458) := X"92440003";
        ram_buffer(24459) := X"0C031190";
        ram_buffer(24460) := X"2484FF80";
        ram_buffer(24461) := X"AFA2001C";
        ram_buffer(24462) := X"92440004";
        ram_buffer(24463) := X"0C031190";
        ram_buffer(24464) := X"2484FF80";
        ram_buffer(24465) := X"AFA20020";
        ram_buffer(24466) := X"92440005";
        ram_buffer(24467) := X"0C031190";
        ram_buffer(24468) := X"2484FF80";
        ram_buffer(24469) := X"AFA20024";
        ram_buffer(24470) := X"92440006";
        ram_buffer(24471) := X"0C031190";
        ram_buffer(24472) := X"2484FF80";
        ram_buffer(24473) := X"AFA20028";
        ram_buffer(24474) := X"92440007";
        ram_buffer(24475) := X"0C031190";
        ram_buffer(24476) := X"2484FF80";
        ram_buffer(24477) := X"8FD20000";
        ram_buffer(24478) := X"AFA2002C";
        ram_buffer(24479) := X"02539021";
        ram_buffer(24480) := X"92440000";
        ram_buffer(24481) := X"0C031190";
        ram_buffer(24482) := X"2484FF80";
        ram_buffer(24483) := X"AFA20030";
        ram_buffer(24484) := X"92440001";
        ram_buffer(24485) := X"0C031190";
        ram_buffer(24486) := X"2484FF80";
        ram_buffer(24487) := X"AFA20034";
        ram_buffer(24488) := X"92440002";
        ram_buffer(24489) := X"0C031190";
        ram_buffer(24490) := X"2484FF80";
        ram_buffer(24491) := X"AFA20038";
        ram_buffer(24492) := X"92440003";
        ram_buffer(24493) := X"0C031190";
        ram_buffer(24494) := X"2484FF80";
        ram_buffer(24495) := X"AFA2003C";
        ram_buffer(24496) := X"92440004";
        ram_buffer(24497) := X"0C031190";
        ram_buffer(24498) := X"2484FF80";
        ram_buffer(24499) := X"AFA20040";
        ram_buffer(24500) := X"92440005";
        ram_buffer(24501) := X"0C031190";
        ram_buffer(24502) := X"2484FF80";
        ram_buffer(24503) := X"AFA20044";
        ram_buffer(24504) := X"92440006";
        ram_buffer(24505) := X"0C031190";
        ram_buffer(24506) := X"2484FF80";
        ram_buffer(24507) := X"AFA20048";
        ram_buffer(24508) := X"92440007";
        ram_buffer(24509) := X"0C031190";
        ram_buffer(24510) := X"2484FF80";
        ram_buffer(24511) := X"8FA3011C";
        ram_buffer(24512) := X"AFA2004C";
        ram_buffer(24513) := X"8C720000";
        ram_buffer(24514) := X"00000000";
        ram_buffer(24515) := X"02539021";
        ram_buffer(24516) := X"92440000";
        ram_buffer(24517) := X"0C031190";
        ram_buffer(24518) := X"2484FF80";
        ram_buffer(24519) := X"AFA20050";
        ram_buffer(24520) := X"92440001";
        ram_buffer(24521) := X"0C031190";
        ram_buffer(24522) := X"2484FF80";
        ram_buffer(24523) := X"AFA20054";
        ram_buffer(24524) := X"92440002";
        ram_buffer(24525) := X"0C031190";
        ram_buffer(24526) := X"2484FF80";
        ram_buffer(24527) := X"AFA20058";
        ram_buffer(24528) := X"92440003";
        ram_buffer(24529) := X"0C031190";
        ram_buffer(24530) := X"2484FF80";
        ram_buffer(24531) := X"AFA2005C";
        ram_buffer(24532) := X"92440004";
        ram_buffer(24533) := X"0C031190";
        ram_buffer(24534) := X"2484FF80";
        ram_buffer(24535) := X"AFA20060";
        ram_buffer(24536) := X"92440005";
        ram_buffer(24537) := X"0C031190";
        ram_buffer(24538) := X"2484FF80";
        ram_buffer(24539) := X"AFA20064";
        ram_buffer(24540) := X"92440006";
        ram_buffer(24541) := X"0C031190";
        ram_buffer(24542) := X"2484FF80";
        ram_buffer(24543) := X"AFA20068";
        ram_buffer(24544) := X"92440007";
        ram_buffer(24545) := X"0C031190";
        ram_buffer(24546) := X"2484FF80";
        ram_buffer(24547) := X"8FA30120";
        ram_buffer(24548) := X"AFA2006C";
        ram_buffer(24549) := X"8C720000";
        ram_buffer(24550) := X"00000000";
        ram_buffer(24551) := X"02539021";
        ram_buffer(24552) := X"92440000";
        ram_buffer(24553) := X"0C031190";
        ram_buffer(24554) := X"2484FF80";
        ram_buffer(24555) := X"AFA20070";
        ram_buffer(24556) := X"92440001";
        ram_buffer(24557) := X"0C031190";
        ram_buffer(24558) := X"2484FF80";
        ram_buffer(24559) := X"AFA20074";
        ram_buffer(24560) := X"92440002";
        ram_buffer(24561) := X"0C031190";
        ram_buffer(24562) := X"2484FF80";
        ram_buffer(24563) := X"AFA20078";
        ram_buffer(24564) := X"92440003";
        ram_buffer(24565) := X"0C031190";
        ram_buffer(24566) := X"2484FF80";
        ram_buffer(24567) := X"AFA2007C";
        ram_buffer(24568) := X"92440004";
        ram_buffer(24569) := X"0C031190";
        ram_buffer(24570) := X"2484FF80";
        ram_buffer(24571) := X"AFA20080";
        ram_buffer(24572) := X"92440005";
        ram_buffer(24573) := X"0C031190";
        ram_buffer(24574) := X"2484FF80";
        ram_buffer(24575) := X"AFA20084";
        ram_buffer(24576) := X"92440006";
        ram_buffer(24577) := X"0C031190";
        ram_buffer(24578) := X"2484FF80";
        ram_buffer(24579) := X"AFA20088";
        ram_buffer(24580) := X"92440007";
        ram_buffer(24581) := X"0C031190";
        ram_buffer(24582) := X"2484FF80";
        ram_buffer(24583) := X"8FA30124";
        ram_buffer(24584) := X"AFA2008C";
        ram_buffer(24585) := X"8C720000";
        ram_buffer(24586) := X"00000000";
        ram_buffer(24587) := X"02539021";
        ram_buffer(24588) := X"92440000";
        ram_buffer(24589) := X"0C031190";
        ram_buffer(24590) := X"2484FF80";
        ram_buffer(24591) := X"AFA20090";
        ram_buffer(24592) := X"92440001";
        ram_buffer(24593) := X"0C031190";
        ram_buffer(24594) := X"2484FF80";
        ram_buffer(24595) := X"AFA20094";
        ram_buffer(24596) := X"92440002";
        ram_buffer(24597) := X"0C031190";
        ram_buffer(24598) := X"2484FF80";
        ram_buffer(24599) := X"AFA20098";
        ram_buffer(24600) := X"92440003";
        ram_buffer(24601) := X"0C031190";
        ram_buffer(24602) := X"2484FF80";
        ram_buffer(24603) := X"AFA2009C";
        ram_buffer(24604) := X"92440004";
        ram_buffer(24605) := X"0C031190";
        ram_buffer(24606) := X"2484FF80";
        ram_buffer(24607) := X"AFA200A0";
        ram_buffer(24608) := X"92440005";
        ram_buffer(24609) := X"0C031190";
        ram_buffer(24610) := X"2484FF80";
        ram_buffer(24611) := X"AFA200A4";
        ram_buffer(24612) := X"92440006";
        ram_buffer(24613) := X"0C031190";
        ram_buffer(24614) := X"2484FF80";
        ram_buffer(24615) := X"AFA200A8";
        ram_buffer(24616) := X"92440007";
        ram_buffer(24617) := X"0C031190";
        ram_buffer(24618) := X"2484FF80";
        ram_buffer(24619) := X"8FA30128";
        ram_buffer(24620) := X"AFA200AC";
        ram_buffer(24621) := X"8C720000";
        ram_buffer(24622) := X"00000000";
        ram_buffer(24623) := X"02539021";
        ram_buffer(24624) := X"92440000";
        ram_buffer(24625) := X"0C031190";
        ram_buffer(24626) := X"2484FF80";
        ram_buffer(24627) := X"AFA200B0";
        ram_buffer(24628) := X"92440001";
        ram_buffer(24629) := X"0C031190";
        ram_buffer(24630) := X"2484FF80";
        ram_buffer(24631) := X"AFA200B4";
        ram_buffer(24632) := X"92440002";
        ram_buffer(24633) := X"0C031190";
        ram_buffer(24634) := X"2484FF80";
        ram_buffer(24635) := X"AFA200B8";
        ram_buffer(24636) := X"92440003";
        ram_buffer(24637) := X"0C031190";
        ram_buffer(24638) := X"2484FF80";
        ram_buffer(24639) := X"AFA200BC";
        ram_buffer(24640) := X"92440004";
        ram_buffer(24641) := X"0C031190";
        ram_buffer(24642) := X"2484FF80";
        ram_buffer(24643) := X"AFA200C0";
        ram_buffer(24644) := X"92440005";
        ram_buffer(24645) := X"0C031190";
        ram_buffer(24646) := X"2484FF80";
        ram_buffer(24647) := X"AFA200C4";
        ram_buffer(24648) := X"92440006";
        ram_buffer(24649) := X"0C031190";
        ram_buffer(24650) := X"2484FF80";
        ram_buffer(24651) := X"AFA200C8";
        ram_buffer(24652) := X"92440007";
        ram_buffer(24653) := X"0C031190";
        ram_buffer(24654) := X"2484FF80";
        ram_buffer(24655) := X"8FA3012C";
        ram_buffer(24656) := X"AFA200CC";
        ram_buffer(24657) := X"8C720000";
        ram_buffer(24658) := X"00000000";
        ram_buffer(24659) := X"02539021";
        ram_buffer(24660) := X"92440000";
        ram_buffer(24661) := X"0C031190";
        ram_buffer(24662) := X"2484FF80";
        ram_buffer(24663) := X"AFA200D0";
        ram_buffer(24664) := X"92440001";
        ram_buffer(24665) := X"0C031190";
        ram_buffer(24666) := X"2484FF80";
        ram_buffer(24667) := X"AFA200D4";
        ram_buffer(24668) := X"92440002";
        ram_buffer(24669) := X"0C031190";
        ram_buffer(24670) := X"2484FF80";
        ram_buffer(24671) := X"AFA200D8";
        ram_buffer(24672) := X"92440003";
        ram_buffer(24673) := X"0C031190";
        ram_buffer(24674) := X"2484FF80";
        ram_buffer(24675) := X"AFA200DC";
        ram_buffer(24676) := X"92440004";
        ram_buffer(24677) := X"0C031190";
        ram_buffer(24678) := X"2484FF80";
        ram_buffer(24679) := X"AFA200E0";
        ram_buffer(24680) := X"92440005";
        ram_buffer(24681) := X"0C031190";
        ram_buffer(24682) := X"2484FF80";
        ram_buffer(24683) := X"AFA200E4";
        ram_buffer(24684) := X"92440006";
        ram_buffer(24685) := X"0C031190";
        ram_buffer(24686) := X"2484FF80";
        ram_buffer(24687) := X"AFA200E8";
        ram_buffer(24688) := X"92440007";
        ram_buffer(24689) := X"0C031190";
        ram_buffer(24690) := X"2484FF80";
        ram_buffer(24691) := X"8FA30130";
        ram_buffer(24692) := X"AFA200EC";
        ram_buffer(24693) := X"8C720000";
        ram_buffer(24694) := X"00000000";
        ram_buffer(24695) := X"02539021";
        ram_buffer(24696) := X"92440000";
        ram_buffer(24697) := X"0C031190";
        ram_buffer(24698) := X"2484FF80";
        ram_buffer(24699) := X"AFA200F0";
        ram_buffer(24700) := X"92440001";
        ram_buffer(24701) := X"0C031190";
        ram_buffer(24702) := X"2484FF80";
        ram_buffer(24703) := X"AFA200F4";
        ram_buffer(24704) := X"92440002";
        ram_buffer(24705) := X"0C031190";
        ram_buffer(24706) := X"2484FF80";
        ram_buffer(24707) := X"AFA200F8";
        ram_buffer(24708) := X"92440003";
        ram_buffer(24709) := X"0C031190";
        ram_buffer(24710) := X"2484FF80";
        ram_buffer(24711) := X"AFA200FC";
        ram_buffer(24712) := X"92440004";
        ram_buffer(24713) := X"0C031190";
        ram_buffer(24714) := X"2484FF80";
        ram_buffer(24715) := X"AFA20100";
        ram_buffer(24716) := X"92440005";
        ram_buffer(24717) := X"0C031190";
        ram_buffer(24718) := X"2484FF80";
        ram_buffer(24719) := X"AFA20104";
        ram_buffer(24720) := X"92440006";
        ram_buffer(24721) := X"0C031190";
        ram_buffer(24722) := X"2484FF80";
        ram_buffer(24723) := X"AFA20108";
        ram_buffer(24724) := X"92440007";
        ram_buffer(24725) := X"27B20010";
        ram_buffer(24726) := X"0C031190";
        ram_buffer(24727) := X"2484FF80";
        ram_buffer(24728) := X"AFA2010C";
        ram_buffer(24729) := X"8FA20110";
        ram_buffer(24730) := X"00000000";
        ram_buffer(24731) := X"0040F809";
        ram_buffer(24732) := X"27A40010";
        ram_buffer(24733) := X"8FB70114";
        ram_buffer(24734) := X"00000000";
        ram_buffer(24735) := X"8EE50000";
        ram_buffer(24736) := X"8E440000";
        ram_buffer(24737) := X"0C030EFE";
        ram_buffer(24738) := X"26520004";
        ram_buffer(24739) := X"00402021";
        ram_buffer(24740) := X"0C030D91";
        ram_buffer(24741) := X"02002821";
        ram_buffer(24742) := X"0C031171";
        ram_buffer(24743) := X"00402021";
        ram_buffer(24744) := X"2442C000";
        ram_buffer(24745) := X"A6C20000";
        ram_buffer(24746) := X"26F70004";
        ram_buffer(24747) := X"1632FFF3";
        ram_buffer(24748) := X"26D60002";
        ram_buffer(24749) := X"8FA20178";
        ram_buffer(24750) := X"26B50001";
        ram_buffer(24751) := X"26730008";
        ram_buffer(24752) := X"1455FEC8";
        ram_buffer(24753) := X"26940080";
        ram_buffer(24754) := X"8FBF015C";
        ram_buffer(24755) := X"8FBE0158";
        ram_buffer(24756) := X"8FB70154";
        ram_buffer(24757) := X"8FB60150";
        ram_buffer(24758) := X"8FB5014C";
        ram_buffer(24759) := X"8FB40148";
        ram_buffer(24760) := X"8FB30144";
        ram_buffer(24761) := X"8FB20140";
        ram_buffer(24762) := X"8FB1013C";
        ram_buffer(24763) := X"8FB00138";
        ram_buffer(24764) := X"03E00008";
        ram_buffer(24765) := X"27BD0160";
        ram_buffer(24766) := X"8C820004";
        ram_buffer(24767) := X"27BDFFE0";
        ram_buffer(24768) := X"8C420000";
        ram_buffer(24769) := X"24060030";
        ram_buffer(24770) := X"AFB10018";
        ram_buffer(24771) := X"AFB00014";
        ram_buffer(24772) := X"AFBF001C";
        ram_buffer(24773) := X"24050001";
        ram_buffer(24774) := X"0040F809";
        ram_buffer(24775) := X"00808821";
        ram_buffer(24776) := X"00408021";
        ram_buffer(24777) := X"AE220160";
        ram_buffer(24778) := X"3C021009";
        ram_buffer(24779) := X"2442707C";
        ram_buffer(24780) := X"8E2300BC";
        ram_buffer(24781) := X"AE020000";
        ram_buffer(24782) := X"24020001";
        ram_buffer(24783) := X"10620024";
        ram_buffer(24784) := X"3C021009";
        ram_buffer(24785) := X"1060001B";
        ram_buffer(24786) := X"24020002";
        ram_buffer(24787) := X"10620013";
        ram_buffer(24788) := X"3C021009";
        ram_buffer(24789) := X"8E220000";
        ram_buffer(24790) := X"2404002F";
        ram_buffer(24791) := X"8C430000";
        ram_buffer(24792) := X"AC440014";
        ram_buffer(24793) := X"0060F809";
        ram_buffer(24794) := X"02202021";
        ram_buffer(24795) := X"2604000C";
        ram_buffer(24796) := X"24060010";
        ram_buffer(24797) := X"0C02801D";
        ram_buffer(24798) := X"00002821";
        ram_buffer(24799) := X"8FBF001C";
        ram_buffer(24800) := X"8FB10018";
        ram_buffer(24801) := X"26040020";
        ram_buffer(24802) := X"8FB00014";
        ram_buffer(24803) := X"24060010";
        ram_buffer(24804) := X"00002821";
        ram_buffer(24805) := X"0802801D";
        ram_buffer(24806) := X"27BD0020";
        ram_buffer(24807) := X"24427D14";
        ram_buffer(24808) := X"AE020004";
        ram_buffer(24809) := X"3C02100A";
        ram_buffer(24810) := X"244286CC";
        ram_buffer(24811) := X"1000FFEF";
        ram_buffer(24812) := X"AE02001C";
        ram_buffer(24813) := X"3C021009";
        ram_buffer(24814) := X"24427750";
        ram_buffer(24815) := X"AE020004";
        ram_buffer(24816) := X"3C02100A";
        ram_buffer(24817) := X"24428BF8";
        ram_buffer(24818) := X"1000FFE8";
        ram_buffer(24819) := X"AE020008";
        ram_buffer(24820) := X"24427750";
        ram_buffer(24821) := X"AE020004";
        ram_buffer(24822) := X"3C02100A";
        ram_buffer(24823) := X"244283E8";
        ram_buffer(24824) := X"1000FFE2";
        ram_buffer(24825) := X"AE020008";
        ram_buffer(24826) := X"27BDFFE0";
        ram_buffer(24827) := X"248C0100";
        ram_buffer(24828) := X"00801021";
        ram_buffer(24829) := X"AFB6001C";
        ram_buffer(24830) := X"AFB50018";
        ram_buffer(24831) := X"AFB40014";
        ram_buffer(24832) := X"AFB30010";
        ram_buffer(24833) := X"AFB2000C";
        ram_buffer(24834) := X"AFB10008";
        ram_buffer(24835) := X"AFB00004";
        ram_buffer(24836) := X"8C4D0000";
        ram_buffer(24837) := X"8C480018";
        ram_buffer(24838) := X"8C46001C";
        ram_buffer(24839) := X"8C4B0004";
        ram_buffer(24840) := X"8C510014";
        ram_buffer(24841) := X"8C43000C";
        ram_buffer(24842) := X"8C470008";
        ram_buffer(24843) := X"8C450010";
        ram_buffer(24844) := X"01A64823";
        ram_buffer(24845) := X"01685023";
        ram_buffer(24846) := X"012AA821";
        ram_buffer(24847) := X"00F17821";
        ram_buffer(24848) := X"0065C021";
        ram_buffer(24849) := X"01685821";
        ram_buffer(24850) := X"00F13823";
        ram_buffer(24851) := X"00652823";
        ram_buffer(24852) := X"01A63021";
        ram_buffer(24853) := X"00A74021";
        ram_buffer(24854) := X"00D86823";
        ram_buffer(24855) := X"01478821";
        ram_buffer(24856) := X"00152940";
        ram_buffer(24857) := X"016F3823";
        ram_buffer(24858) := X"001518C0";
        ram_buffer(24859) := X"00ED8021";
        ram_buffer(24860) := X"00A31823";
        ram_buffer(24861) := X"01159023";
        ram_buffer(24862) := X"00083880";
        ram_buffer(24863) := X"00082900";
        ram_buffer(24864) := X"00115080";
        ram_buffer(24865) := X"00117100";
        ram_buffer(24866) := X"00E5B021";
        ram_buffer(24867) := X"01CAA023";
        ram_buffer(24868) := X"00103880";
        ram_buffer(24869) := X"00105100";
        ram_buffer(24870) := X"0012C840";
        ram_buffer(24871) := X"000328C0";
        ram_buffer(24872) := X"00129100";
        ram_buffer(24873) := X"01479823";
        ram_buffer(24874) := X"0259C823";
        ram_buffer(24875) := X"00A32823";
        ram_buffer(24876) := X"001638C0";
        ram_buffer(24877) := X"00147100";
        ram_buffer(24878) := X"00F63823";
        ram_buffer(24879) := X"00B51823";
        ram_buffer(24880) := X"01D47023";
        ram_buffer(24881) := X"00135100";
        ram_buffer(24882) := X"001990C0";
        ram_buffer(24883) := X"00E82823";
        ram_buffer(24884) := X"01535023";
        ram_buffer(24885) := X"01D14021";
        ram_buffer(24886) := X"0259C823";
        ram_buffer(24887) := X"00031840";
        ram_buffer(24888) := X"00084203";
        ram_buffer(24889) := X"0019CA03";
        ram_buffer(24890) := X"01503821";
        ram_buffer(24891) := X"00052A03";
        ram_buffer(24892) := X"00031A03";
        ram_buffer(24893) := X"01285021";
        ram_buffer(24894) := X"016F5821";
        ram_buffer(24895) := X"00B92821";
        ram_buffer(24896) := X"00D83021";
        ram_buffer(24897) := X"00073A03";
        ram_buffer(24898) := X"00791821";
        ram_buffer(24899) := X"01284823";
        ram_buffer(24900) := X"00CB7021";
        ram_buffer(24901) := X"00A94021";
        ram_buffer(24902) := X"00CB3023";
        ram_buffer(24903) := X"01254823";
        ram_buffer(24904) := X"01A75821";
        ram_buffer(24905) := X"006A2821";
        ram_buffer(24906) := X"01A73823";
        ram_buffer(24907) := X"01431823";
        ram_buffer(24908) := X"AC4E0000";
        ram_buffer(24909) := X"AC460010";
        ram_buffer(24910) := X"AC4B0008";
        ram_buffer(24911) := X"AC470018";
        ram_buffer(24912) := X"AC480014";
        ram_buffer(24913) := X"AC49000C";
        ram_buffer(24914) := X"AC450004";
        ram_buffer(24915) := X"AC43001C";
        ram_buffer(24916) := X"24420020";
        ram_buffer(24917) := X"144CFFAE";
        ram_buffer(24918) := X"24890020";
        ram_buffer(24919) := X"8C8700E0";
        ram_buffer(24920) := X"8C8A00C0";
        ram_buffer(24921) := X"8C8C0000";
        ram_buffer(24922) := X"8C8D0020";
        ram_buffer(24923) := X"8C880040";
        ram_buffer(24924) := X"8C860080";
        ram_buffer(24925) := X"8C8500A0";
        ram_buffer(24926) := X"8C830060";
        ram_buffer(24927) := X"01875823";
        ram_buffer(24928) := X"01AAC023";
        ram_buffer(24929) := X"01781021";
        ram_buffer(24930) := X"01876021";
        ram_buffer(24931) := X"01057021";
        ram_buffer(24932) := X"00667821";
        ram_buffer(24933) := X"01052823";
        ram_buffer(24934) := X"01AA6821";
        ram_buffer(24935) := X"00661823";
        ram_buffer(24936) := X"00653021";
        ram_buffer(24937) := X"018F5023";
        ram_buffer(24938) := X"03058821";
        ram_buffer(24939) := X"000218C0";
        ram_buffer(24940) := X"01AEC823";
        ram_buffer(24941) := X"00028140";
        ram_buffer(24942) := X"032AC821";
        ram_buffer(24943) := X"00C2A823";
        ram_buffer(24944) := X"02038023";
        ram_buffer(24945) := X"00062880";
        ram_buffer(24946) := X"00061900";
        ram_buffer(24947) := X"00113880";
        ram_buffer(24948) := X"00114100";
        ram_buffer(24949) := X"00A3A021";
        ram_buffer(24950) := X"01079823";
        ram_buffer(24951) := X"00192880";
        ram_buffer(24952) := X"00193900";
        ram_buffer(24953) := X"0015C040";
        ram_buffer(24954) := X"001018C0";
        ram_buffer(24955) := X"0015A900";
        ram_buffer(24956) := X"00E59023";
        ram_buffer(24957) := X"00701823";
        ram_buffer(24958) := X"02B8C023";
        ram_buffer(24959) := X"001428C0";
        ram_buffer(24960) := X"00134100";
        ram_buffer(24961) := X"00B42823";
        ram_buffer(24962) := X"00621023";
        ram_buffer(24963) := X"01134023";
        ram_buffer(24964) := X"00123900";
        ram_buffer(24965) := X"001880C0";
        ram_buffer(24966) := X"00A61823";
        ram_buffer(24967) := X"00F23823";
        ram_buffer(24968) := X"01112821";
        ram_buffer(24969) := X"0218C023";
        ram_buffer(24970) := X"00021040";
        ram_buffer(24971) := X"0018C203";
        ram_buffer(24972) := X"00052A03";
        ram_buffer(24973) := X"00F93021";
        ram_buffer(24974) := X"00031A03";
        ram_buffer(24975) := X"00021203";
        ram_buffer(24976) := X"01654021";
        ram_buffer(24977) := X"018F3821";
        ram_buffer(24978) := X"01652823";
        ram_buffer(24979) := X"01AE6821";
        ram_buffer(24980) := X"00063203";
        ram_buffer(24981) := X"00781821";
        ram_buffer(24982) := X"00581021";
        ram_buffer(24983) := X"01465821";
        ram_buffer(24984) := X"00ED6021";
        ram_buffer(24985) := X"01463023";
        ram_buffer(24986) := X"00ED3823";
        ram_buffer(24987) := X"00655021";
        ram_buffer(24988) := X"00A31823";
        ram_buffer(24989) := X"00482821";
        ram_buffer(24990) := X"01021023";
        ram_buffer(24991) := X"AC8C0000";
        ram_buffer(24992) := X"AC870080";
        ram_buffer(24993) := X"AC8B0040";
        ram_buffer(24994) := X"AC8600C0";
        ram_buffer(24995) := X"AC8A00A0";
        ram_buffer(24996) := X"AC830060";
        ram_buffer(24997) := X"AC850020";
        ram_buffer(24998) := X"AC8200E0";
        ram_buffer(24999) := X"24840004";
        ram_buffer(25000) := X"1489FFAE";
        ram_buffer(25001) := X"00000000";
        ram_buffer(25002) := X"8FB6001C";
        ram_buffer(25003) := X"8FB50018";
        ram_buffer(25004) := X"8FB40014";
        ram_buffer(25005) := X"8FB30010";
        ram_buffer(25006) := X"8FB2000C";
        ram_buffer(25007) := X"8FB10008";
        ram_buffer(25008) := X"8FB00004";
        ram_buffer(25009) := X"03E00008";
        ram_buffer(25010) := X"27BD0020";
        ram_buffer(25011) := X"8F838074";
        ram_buffer(25012) := X"27BDFFA0";
        ram_buffer(25013) := X"AFA30020";
        ram_buffer(25014) := X"8F838078";
        ram_buffer(25015) := X"8F828070";
        ram_buffer(25016) := X"AFA30024";
        ram_buffer(25017) := X"8F83807C";
        ram_buffer(25018) := X"AFB1003C";
        ram_buffer(25019) := X"AFA30028";
        ram_buffer(25020) := X"24830100";
        ram_buffer(25021) := X"AFB00038";
        ram_buffer(25022) := X"AFBF005C";
        ram_buffer(25023) := X"AFBE0058";
        ram_buffer(25024) := X"AFB70054";
        ram_buffer(25025) := X"AFB60050";
        ram_buffer(25026) := X"AFB5004C";
        ram_buffer(25027) := X"AFB40048";
        ram_buffer(25028) := X"AFB30044";
        ram_buffer(25029) := X"AFB20040";
        ram_buffer(25030) := X"AFA2001C";
        ram_buffer(25031) := X"00808021";
        ram_buffer(25032) := X"AFA3002C";
        ram_buffer(25033) := X"00808821";
        ram_buffer(25034) := X"AFA20030";
        ram_buffer(25035) := X"8E320000";
        ram_buffer(25036) := X"8E34001C";
        ram_buffer(25037) := X"02402021";
        ram_buffer(25038) := X"0C030D91";
        ram_buffer(25039) := X"02802821";
        ram_buffer(25040) := X"02802821";
        ram_buffer(25041) := X"02402021";
        ram_buffer(25042) := X"0C030FF2";
        ram_buffer(25043) := X"00409821";
        ram_buffer(25044) := X"8E350018";
        ram_buffer(25045) := X"8E340004";
        ram_buffer(25046) := X"02A02821";
        ram_buffer(25047) := X"02802021";
        ram_buffer(25048) := X"0C030D91";
        ram_buffer(25049) := X"00409021";
        ram_buffer(25050) := X"02A02821";
        ram_buffer(25051) := X"02802021";
        ram_buffer(25052) := X"0C030FF2";
        ram_buffer(25053) := X"0040B021";
        ram_buffer(25054) := X"8E350008";
        ram_buffer(25055) := X"8E3E0014";
        ram_buffer(25056) := X"02A02021";
        ram_buffer(25057) := X"03C02821";
        ram_buffer(25058) := X"0C030D91";
        ram_buffer(25059) := X"0040A021";
        ram_buffer(25060) := X"03C02821";
        ram_buffer(25061) := X"02A02021";
        ram_buffer(25062) := X"0C030FF2";
        ram_buffer(25063) := X"0040B821";
        ram_buffer(25064) := X"8E260010";
        ram_buffer(25065) := X"8E23000C";
        ram_buffer(25066) := X"00C02821";
        ram_buffer(25067) := X"00602021";
        ram_buffer(25068) := X"AFA60018";
        ram_buffer(25069) := X"AFA30014";
        ram_buffer(25070) := X"0C030D91";
        ram_buffer(25071) := X"0040A821";
        ram_buffer(25072) := X"00402821";
        ram_buffer(25073) := X"02602021";
        ram_buffer(25074) := X"0C030D91";
        ram_buffer(25075) := X"AFA20010";
        ram_buffer(25076) := X"8FA70010";
        ram_buffer(25077) := X"02602021";
        ram_buffer(25078) := X"00E02821";
        ram_buffer(25079) := X"0C030FF2";
        ram_buffer(25080) := X"0040F021";
        ram_buffer(25081) := X"02E02821";
        ram_buffer(25082) := X"02C02021";
        ram_buffer(25083) := X"0C030D91";
        ram_buffer(25084) := X"00409821";
        ram_buffer(25085) := X"00402821";
        ram_buffer(25086) := X"03C02021";
        ram_buffer(25087) := X"0C030D91";
        ram_buffer(25088) := X"AFA20010";
        ram_buffer(25089) := X"8FA70010";
        ram_buffer(25090) := X"AE220000";
        ram_buffer(25091) := X"00E02821";
        ram_buffer(25092) := X"0C030FF2";
        ram_buffer(25093) := X"03C02021";
        ram_buffer(25094) := X"AE220010";
        ram_buffer(25095) := X"02E02821";
        ram_buffer(25096) := X"0C030FF2";
        ram_buffer(25097) := X"02C02021";
        ram_buffer(25098) := X"00402021";
        ram_buffer(25099) := X"0C030D91";
        ram_buffer(25100) := X"02602821";
        ram_buffer(25101) := X"8FA5001C";
        ram_buffer(25102) := X"0C030EFE";
        ram_buffer(25103) := X"00402021";
        ram_buffer(25104) := X"00402821";
        ram_buffer(25105) := X"02602021";
        ram_buffer(25106) := X"0C030D91";
        ram_buffer(25107) := X"0040B021";
        ram_buffer(25108) := X"AE220008";
        ram_buffer(25109) := X"02C02821";
        ram_buffer(25110) := X"0C030FF2";
        ram_buffer(25111) := X"02602021";
        ram_buffer(25112) := X"8FA60018";
        ram_buffer(25113) := X"8FA30014";
        ram_buffer(25114) := X"00C02821";
        ram_buffer(25115) := X"00602021";
        ram_buffer(25116) := X"0C030FF2";
        ram_buffer(25117) := X"AE220018";
        ram_buffer(25118) := X"00402021";
        ram_buffer(25119) := X"0C030D91";
        ram_buffer(25120) := X"02A02821";
        ram_buffer(25121) := X"02802821";
        ram_buffer(25122) := X"02402021";
        ram_buffer(25123) := X"0C030D91";
        ram_buffer(25124) := X"0040B021";
        ram_buffer(25125) := X"00402821";
        ram_buffer(25126) := X"02C02021";
        ram_buffer(25127) := X"0C030FF2";
        ram_buffer(25128) := X"0040B821";
        ram_buffer(25129) := X"8FA50020";
        ram_buffer(25130) := X"0C030EFE";
        ram_buffer(25131) := X"00402021";
        ram_buffer(25132) := X"8FA50024";
        ram_buffer(25133) := X"02C02021";
        ram_buffer(25134) := X"0C030EFE";
        ram_buffer(25135) := X"00409821";
        ram_buffer(25136) := X"00402021";
        ram_buffer(25137) := X"0C030D91";
        ram_buffer(25138) := X"02602821";
        ram_buffer(25139) := X"8FA50028";
        ram_buffer(25140) := X"02E02021";
        ram_buffer(25141) := X"0C030EFE";
        ram_buffer(25142) := X"0040B021";
        ram_buffer(25143) := X"00402021";
        ram_buffer(25144) := X"0C030D91";
        ram_buffer(25145) := X"02602821";
        ram_buffer(25146) := X"02A02821";
        ram_buffer(25147) := X"02802021";
        ram_buffer(25148) := X"0C030D91";
        ram_buffer(25149) := X"00409821";
        ram_buffer(25150) := X"8FA50030";
        ram_buffer(25151) := X"0C030EFE";
        ram_buffer(25152) := X"00402021";
        ram_buffer(25153) := X"0040A821";
        ram_buffer(25154) := X"02402021";
        ram_buffer(25155) := X"0C030D91";
        ram_buffer(25156) := X"00402821";
        ram_buffer(25157) := X"02402021";
        ram_buffer(25158) := X"02A02821";
        ram_buffer(25159) := X"0C030FF2";
        ram_buffer(25160) := X"0040A021";
        ram_buffer(25161) := X"00402821";
        ram_buffer(25162) := X"02C02021";
        ram_buffer(25163) := X"0C030D91";
        ram_buffer(25164) := X"00409021";
        ram_buffer(25165) := X"AE220014";
        ram_buffer(25166) := X"02C02821";
        ram_buffer(25167) := X"0C030FF2";
        ram_buffer(25168) := X"02402021";
        ram_buffer(25169) := X"AE22000C";
        ram_buffer(25170) := X"02802821";
        ram_buffer(25171) := X"0C030D91";
        ram_buffer(25172) := X"02602021";
        ram_buffer(25173) := X"AE220004";
        ram_buffer(25174) := X"02602821";
        ram_buffer(25175) := X"0C030FF2";
        ram_buffer(25176) := X"02802021";
        ram_buffer(25177) := X"AE22001C";
        ram_buffer(25178) := X"8FA2002C";
        ram_buffer(25179) := X"26310020";
        ram_buffer(25180) := X"1622FF6E";
        ram_buffer(25181) := X"26030020";
        ram_buffer(25182) := X"8FA2001C";
        ram_buffer(25183) := X"AFA30018";
        ram_buffer(25184) := X"AFA2002C";
        ram_buffer(25185) := X"8E110000";
        ram_buffer(25186) := X"8E1300E0";
        ram_buffer(25187) := X"02202021";
        ram_buffer(25188) := X"0C030D91";
        ram_buffer(25189) := X"02602821";
        ram_buffer(25190) := X"02602821";
        ram_buffer(25191) := X"02202021";
        ram_buffer(25192) := X"0C030FF2";
        ram_buffer(25193) := X"00409021";
        ram_buffer(25194) := X"8E1400C0";
        ram_buffer(25195) := X"8E130020";
        ram_buffer(25196) := X"02802821";
        ram_buffer(25197) := X"02602021";
        ram_buffer(25198) := X"0C030D91";
        ram_buffer(25199) := X"00408821";
        ram_buffer(25200) := X"02802821";
        ram_buffer(25201) := X"02602021";
        ram_buffer(25202) := X"0C030FF2";
        ram_buffer(25203) := X"0040B021";
        ram_buffer(25204) := X"8E140040";
        ram_buffer(25205) := X"8E1E00A0";
        ram_buffer(25206) := X"02802021";
        ram_buffer(25207) := X"03C02821";
        ram_buffer(25208) := X"0C030D91";
        ram_buffer(25209) := X"00409821";
        ram_buffer(25210) := X"03C02821";
        ram_buffer(25211) := X"02802021";
        ram_buffer(25212) := X"0C030FF2";
        ram_buffer(25213) := X"0040B821";
        ram_buffer(25214) := X"8E060080";
        ram_buffer(25215) := X"8E150060";
        ram_buffer(25216) := X"00C02821";
        ram_buffer(25217) := X"02A02021";
        ram_buffer(25218) := X"AFA60014";
        ram_buffer(25219) := X"0C030D91";
        ram_buffer(25220) := X"0040A021";
        ram_buffer(25221) := X"00402821";
        ram_buffer(25222) := X"02402021";
        ram_buffer(25223) := X"0C030D91";
        ram_buffer(25224) := X"AFA20010";
        ram_buffer(25225) := X"8FA70010";
        ram_buffer(25226) := X"02402021";
        ram_buffer(25227) := X"00E02821";
        ram_buffer(25228) := X"0C030FF2";
        ram_buffer(25229) := X"0040F021";
        ram_buffer(25230) := X"02E02821";
        ram_buffer(25231) := X"02C02021";
        ram_buffer(25232) := X"0C030D91";
        ram_buffer(25233) := X"00409021";
        ram_buffer(25234) := X"00402821";
        ram_buffer(25235) := X"03C02021";
        ram_buffer(25236) := X"0C030D91";
        ram_buffer(25237) := X"AFA20010";
        ram_buffer(25238) := X"8FA70010";
        ram_buffer(25239) := X"AE020000";
        ram_buffer(25240) := X"00E02821";
        ram_buffer(25241) := X"0C030FF2";
        ram_buffer(25242) := X"03C02021";
        ram_buffer(25243) := X"AE020080";
        ram_buffer(25244) := X"02E02821";
        ram_buffer(25245) := X"0C030FF2";
        ram_buffer(25246) := X"02C02021";
        ram_buffer(25247) := X"00402021";
        ram_buffer(25248) := X"0C030D91";
        ram_buffer(25249) := X"02402821";
        ram_buffer(25250) := X"8FA5001C";
        ram_buffer(25251) := X"0C030EFE";
        ram_buffer(25252) := X"00402021";
        ram_buffer(25253) := X"00402821";
        ram_buffer(25254) := X"02402021";
        ram_buffer(25255) := X"0C030D91";
        ram_buffer(25256) := X"0040B021";
        ram_buffer(25257) := X"AE020040";
        ram_buffer(25258) := X"02C02821";
        ram_buffer(25259) := X"0C030FF2";
        ram_buffer(25260) := X"02402021";
        ram_buffer(25261) := X"8FA60014";
        ram_buffer(25262) := X"AE0200C0";
        ram_buffer(25263) := X"00C02821";
        ram_buffer(25264) := X"0C030FF2";
        ram_buffer(25265) := X"02A02021";
        ram_buffer(25266) := X"00402021";
        ram_buffer(25267) := X"0C030D91";
        ram_buffer(25268) := X"02802821";
        ram_buffer(25269) := X"02602821";
        ram_buffer(25270) := X"02202021";
        ram_buffer(25271) := X"0C030D91";
        ram_buffer(25272) := X"0040B021";
        ram_buffer(25273) := X"00402821";
        ram_buffer(25274) := X"02C02021";
        ram_buffer(25275) := X"0C030FF2";
        ram_buffer(25276) := X"0040B821";
        ram_buffer(25277) := X"8FA50020";
        ram_buffer(25278) := X"0C030EFE";
        ram_buffer(25279) := X"00402021";
        ram_buffer(25280) := X"8FA50024";
        ram_buffer(25281) := X"02C02021";
        ram_buffer(25282) := X"0C030EFE";
        ram_buffer(25283) := X"00409021";
        ram_buffer(25284) := X"00402021";
        ram_buffer(25285) := X"0C030D91";
        ram_buffer(25286) := X"02402821";
        ram_buffer(25287) := X"8FA50028";
        ram_buffer(25288) := X"02E02021";
        ram_buffer(25289) := X"0C030EFE";
        ram_buffer(25290) := X"0040B021";
        ram_buffer(25291) := X"00402021";
        ram_buffer(25292) := X"0C030D91";
        ram_buffer(25293) := X"02402821";
        ram_buffer(25294) := X"02802821";
        ram_buffer(25295) := X"02602021";
        ram_buffer(25296) := X"0C030D91";
        ram_buffer(25297) := X"00409021";
        ram_buffer(25298) := X"8FA5002C";
        ram_buffer(25299) := X"0C030EFE";
        ram_buffer(25300) := X"00402021";
        ram_buffer(25301) := X"0040A021";
        ram_buffer(25302) := X"02202021";
        ram_buffer(25303) := X"0C030D91";
        ram_buffer(25304) := X"00402821";
        ram_buffer(25305) := X"02202021";
        ram_buffer(25306) := X"02802821";
        ram_buffer(25307) := X"0C030FF2";
        ram_buffer(25308) := X"00409821";
        ram_buffer(25309) := X"00402821";
        ram_buffer(25310) := X"02C02021";
        ram_buffer(25311) := X"0C030D91";
        ram_buffer(25312) := X"00408821";
        ram_buffer(25313) := X"AE0200A0";
        ram_buffer(25314) := X"02C02821";
        ram_buffer(25315) := X"0C030FF2";
        ram_buffer(25316) := X"02202021";
        ram_buffer(25317) := X"AE020060";
        ram_buffer(25318) := X"02602821";
        ram_buffer(25319) := X"0C030D91";
        ram_buffer(25320) := X"02402021";
        ram_buffer(25321) := X"AE020020";
        ram_buffer(25322) := X"02402821";
        ram_buffer(25323) := X"0C030FF2";
        ram_buffer(25324) := X"02602021";
        ram_buffer(25325) := X"AE0200E0";
        ram_buffer(25326) := X"8FA20018";
        ram_buffer(25327) := X"26100004";
        ram_buffer(25328) := X"1602FF70";
        ram_buffer(25329) := X"00000000";
        ram_buffer(25330) := X"8FBF005C";
        ram_buffer(25331) := X"8FBE0058";
        ram_buffer(25332) := X"8FB70054";
        ram_buffer(25333) := X"8FB60050";
        ram_buffer(25334) := X"8FB5004C";
        ram_buffer(25335) := X"8FB40048";
        ram_buffer(25336) := X"8FB30044";
        ram_buffer(25337) := X"8FB20040";
        ram_buffer(25338) := X"8FB1003C";
        ram_buffer(25339) := X"8FB00038";
        ram_buffer(25340) := X"03E00008";
        ram_buffer(25341) := X"27BD0060";
        ram_buffer(25342) := X"27BDFFC0";
        ram_buffer(25343) := X"24820100";
        ram_buffer(25344) := X"00805821";
        ram_buffer(25345) := X"AFBE003C";
        ram_buffer(25346) := X"AFB70038";
        ram_buffer(25347) := X"AFB60034";
        ram_buffer(25348) := X"AFB50030";
        ram_buffer(25349) := X"AFB4002C";
        ram_buffer(25350) := X"AFB30028";
        ram_buffer(25351) := X"AFB20024";
        ram_buffer(25352) := X"AFB10020";
        ram_buffer(25353) := X"AFB0001C";
        ram_buffer(25354) := X"AFA20014";
        ram_buffer(25355) := X"AFA40040";
        ram_buffer(25356) := X"8D6C0000";
        ram_buffer(25357) := X"8D65000C";
        ram_buffer(25358) := X"8D66001C";
        ram_buffer(25359) := X"8D630010";
        ram_buffer(25360) := X"0186C823";
        ram_buffer(25361) := X"00A38023";
        ram_buffer(25362) := X"03301021";
        ram_buffer(25363) := X"2407E333";
        ram_buffer(25364) := X"00470018";
        ram_buffer(25365) := X"8D6A0004";
        ram_buffer(25366) := X"8D680008";
        ram_buffer(25367) := X"8D690018";
        ram_buffer(25368) := X"8D640014";
        ram_buffer(25369) := X"01497023";
        ram_buffer(25370) := X"01047823";
        ram_buffer(25371) := X"01D0C021";
        ram_buffer(25372) := X"032F3821";
        ram_buffer(25373) := X"01CFF021";
        ram_buffer(25374) := X"000F6980";
        ram_buffer(25375) := X"01494821";
        ram_buffer(25376) := X"01042021";
        ram_buffer(25377) := X"00A31821";
        ram_buffer(25378) := X"000F10C0";
        ram_buffer(25379) := X"01863021";
        ram_buffer(25380) := X"03078821";
        ram_buffer(25381) := X"01209021";
        ram_buffer(25382) := X"00809821";
        ram_buffer(25383) := X"0060A021";
        ram_buffer(25384) := X"01A21023";
        ram_buffer(25385) := X"001E4140";
        ram_buffer(25386) := X"000E2080";
        ram_buffer(25387) := X"00C06021";
        ram_buffer(25388) := X"001E5080";
        ram_buffer(25389) := X"000E4900";
        ram_buffer(25390) := X"02536823";
        ram_buffer(25391) := X"01244823";
        ram_buffer(25392) := X"01485021";
        ram_buffer(25393) := X"00113100";
        ram_buffer(25394) := X"00182A00";
        ram_buffer(25395) := X"00022100";
        ram_buffer(25396) := X"AFAC0000";
        ram_buffer(25397) := X"00114080";
        ram_buffer(25398) := X"01946023";
        ram_buffer(25399) := X"00181880";
        ram_buffer(25400) := X"01064021";
        ram_buffer(25401) := X"AFB20004";
        ram_buffer(25402) := X"AFB30008";
        ram_buffer(25403) := X"01809021";
        ram_buffer(25404) := X"000799C0";
        ram_buffer(25405) := X"000D6180";
        ram_buffer(25406) := X"AFB4000C";
        ram_buffer(25407) := X"000D3080";
        ram_buffer(25408) := X"000AB0C0";
        ram_buffer(25409) := X"00A31823";
        ram_buffer(25410) := X"0007A940";
        ram_buffer(25411) := X"00102980";
        ram_buffer(25412) := X"00821023";
        ram_buffer(25413) := X"0010A0C0";
        ram_buffer(25414) := X"00092100";
        ram_buffer(25415) := X"024DB821";
        ram_buffer(25416) := X"0285A021";
        ram_buffer(25417) := X"02B3A821";
        ram_buffer(25418) := X"004F1021";
        ram_buffer(25419) := X"00122980";
        ram_buffer(25420) := X"AFB20010";
        ram_buffer(25421) := X"00129A40";
        ram_buffer(25422) := X"01863023";
        ram_buffer(25423) := X"01565021";
        ram_buffer(25424) := X"00086100";
        ram_buffer(25425) := X"0019B080";
        ram_buffer(25426) := X"01242021";
        ram_buffer(25427) := X"00199100";
        ram_buffer(25428) := X"00781823";
        ram_buffer(25429) := X"008E4823";
        ram_buffer(25430) := X"015E5023";
        ram_buffer(25431) := X"02569023";
        ram_buffer(25432) := X"00CD3023";
        ram_buffer(25433) := X"01884023";
        ram_buffer(25434) := X"0015B080";
        ram_buffer(25435) := X"00142100";
        ram_buffer(25436) := X"00031900";
        ram_buffer(25437) := X"0002F080";
        ram_buffer(25438) := X"02659823";
        ram_buffer(25439) := X"00177100";
        ram_buffer(25440) := X"001729C0";
        ram_buffer(25441) := X"000A6180";
        ram_buffer(25442) := X"02B6A821";
        ram_buffer(25443) := X"02842021";
        ram_buffer(25444) := X"000630C0";
        ram_buffer(25445) := X"0012A280";
        ram_buffer(25446) := X"01114021";
        ram_buffer(25447) := X"00781821";
        ram_buffer(25448) := X"005E1021";
        ram_buffer(25449) := X"01C57021";
        ram_buffer(25450) := X"00CD3021";
        ram_buffer(25451) := X"001328C0";
        ram_buffer(25452) := X"014C5021";
        ram_buffer(25453) := X"00F5A823";
        ram_buffer(25454) := X"00021080";
        ram_buffer(25455) := X"02549021";
        ram_buffer(25456) := X"8FAC0010";
        ram_buffer(25457) := X"0009B140";
        ram_buffer(25458) := X"00084140";
        ram_buffer(25459) := X"00031880";
        ram_buffer(25460) := X"01D77023";
        ram_buffer(25461) := X"00B32823";
        ram_buffer(25462) := X"01114021";
        ram_buffer(25463) := X"004F7823";
        ram_buffer(25464) := X"00902023";
        ram_buffer(25465) := X"00001012";
        ram_buffer(25466) := X"02C94823";
        ram_buffer(25467) := X"00063140";
        ram_buffer(25468) := X"00781821";
        ram_buffer(25469) := X"0015A880";
        ram_buffer(25470) := X"02599023";
        ram_buffer(25471) := X"000A5023";
        ram_buffer(25472) := X"01031823";
        ram_buffer(25473) := X"00CD3021";
        ram_buffer(25474) := X"00AC2823";
        ram_buffer(25475) := X"00042040";
        ram_buffer(25476) := X"01154021";
        ram_buffer(25477) := X"8FAC0000";
        ram_buffer(25478) := X"000EB940";
        ram_buffer(25479) := X"00094880";
        ram_buffer(25480) := X"0242C821";
        ram_buffer(25481) := X"8FB4000C";
        ram_buffer(25482) := X"8FAD0004";
        ram_buffer(25483) := X"8FB30008";
        ram_buffer(25484) := X"00823821";
        ram_buffer(25485) := X"02EE7023";
        ram_buffer(25486) := X"01EA2021";
        ram_buffer(25487) := X"012A4821";
        ram_buffer(25488) := X"00052840";
        ram_buffer(25489) := X"03281021";
        ram_buffer(25490) := X"01945021";
        ram_buffer(25491) := X"00AE2821";
        ram_buffer(25492) := X"01B36021";
        ram_buffer(25493) := X"01C67023";
        ram_buffer(25494) := X"00E33821";
        ram_buffer(25495) := X"00882021";
        ram_buffer(25496) := X"01231821";
        ram_buffer(25497) := X"24420400";
        ram_buffer(25498) := X"014C3021";
        ram_buffer(25499) := X"000212C3";
        ram_buffer(25500) := X"014C5023";
        ram_buffer(25501) := X"24A50400";
        ram_buffer(25502) := X"25CE0400";
        ram_buffer(25503) := X"24E70400";
        ram_buffer(25504) := X"24840400";
        ram_buffer(25505) := X"24630400";
        ram_buffer(25506) := X"AD620004";
        ram_buffer(25507) := X"00063080";
        ram_buffer(25508) := X"000A5080";
        ram_buffer(25509) := X"00052AC3";
        ram_buffer(25510) := X"000E72C3";
        ram_buffer(25511) := X"00073AC3";
        ram_buffer(25512) := X"000422C3";
        ram_buffer(25513) := X"00031AC3";
        ram_buffer(25514) := X"8FA20014";
        ram_buffer(25515) := X"AD660000";
        ram_buffer(25516) := X"AD6A0010";
        ram_buffer(25517) := X"AD650008";
        ram_buffer(25518) := X"AD6E0018";
        ram_buffer(25519) := X"AD67001C";
        ram_buffer(25520) := X"AD640014";
        ram_buffer(25521) := X"AD63000C";
        ram_buffer(25522) := X"256B0020";
        ram_buffer(25523) := X"1562FF58";
        ram_buffer(25524) := X"00000000";
        ram_buffer(25525) := X"8FAD0040";
        ram_buffer(25526) := X"00000000";
        ram_buffer(25527) := X"25A20020";
        ram_buffer(25528) := X"AFA20014";
        ram_buffer(25529) := X"8DB00000";
        ram_buffer(25530) := X"8DA70060";
        ram_buffer(25531) := X"8DAA00E0";
        ram_buffer(25532) := X"8DA50080";
        ram_buffer(25533) := X"020AC023";
        ram_buffer(25534) := X"00E5C823";
        ram_buffer(25535) := X"8DAB0020";
        ram_buffer(25536) := X"8DA80040";
        ram_buffer(25537) := X"8DA900C0";
        ram_buffer(25538) := X"8DA300A0";
        ram_buffer(25539) := X"03191021";
        ram_buffer(25540) := X"2404E333";
        ram_buffer(25541) := X"01037023";
        ram_buffer(25542) := X"01696023";
        ram_buffer(25543) := X"00440018";
        ram_buffer(25544) := X"018EF021";
        ram_buffer(25545) := X"000E10C0";
        ram_buffer(25546) := X"01031821";
        ram_buffer(25547) := X"000E2180";
        ram_buffer(25548) := X"01694821";
        ram_buffer(25549) := X"01997821";
        ram_buffer(25550) := X"030E3021";
        ram_buffer(25551) := X"00609021";
        ram_buffer(25552) := X"01205821";
        ram_buffer(25553) := X"00822023";
        ram_buffer(25554) := X"001E1940";
        ram_buffer(25555) := X"001E4880";
        ram_buffer(25556) := X"01E68821";
        ram_buffer(25557) := X"000C1080";
        ram_buffer(25558) := X"00E52821";
        ram_buffer(25559) := X"01234821";
        ram_buffer(25560) := X"000C4100";
        ram_buffer(25561) := X"00041900";
        ram_buffer(25562) := X"020A5021";
        ram_buffer(25563) := X"01024023";
        ram_buffer(25564) := X"00A08021";
        ram_buffer(25565) := X"000F9A00";
        ram_buffer(25566) := X"AFAB0008";
        ram_buffer(25567) := X"00112900";
        ram_buffer(25568) := X"01725823";
        ram_buffer(25569) := X"000F1080";
        ram_buffer(25570) := X"00642023";
        ram_buffer(25571) := X"00113880";
        ram_buffer(25572) := X"00E53821";
        ram_buffer(25573) := X"008E2021";
        ram_buffer(25574) := X"AFAA0004";
        ram_buffer(25575) := X"AFB00010";
        ram_buffer(25576) := X"000B2880";
        ram_buffer(25577) := X"01508023";
        ram_buffer(25578) := X"0009B0C0";
        ram_buffer(25579) := X"000B5180";
        ram_buffer(25580) := X"02621023";
        ram_buffer(25581) := X"0019A0C0";
        ram_buffer(25582) := X"00199980";
        ram_buffer(25583) := X"00081900";
        ram_buffer(25584) := X"0293A021";
        ram_buffer(25585) := X"AFA40000";
        ram_buffer(25586) := X"01452823";
        ram_buffer(25587) := X"01364821";
        ram_buffer(25588) := X"004F1023";
        ram_buffer(25589) := X"01031821";
        ram_buffer(25590) := X"006C4023";
        ram_buffer(25591) := X"013E4823";
        ram_buffer(25592) := X"AFB2000C";
        ram_buffer(25593) := X"0006A9C0";
        ram_buffer(25594) := X"00069140";
        ram_buffer(25595) := X"00AB2823";
        ram_buffer(25596) := X"00141900";
        ram_buffer(25597) := X"00021100";
        ram_buffer(25598) := X"8FBE0000";
        ram_buffer(25599) := X"020BB821";
        ram_buffer(25600) := X"0255A821";
        ram_buffer(25601) := X"00102180";
        ram_buffer(25602) := X"0018B080";
        ram_buffer(25603) := X"00109A40";
        ram_buffer(25604) := X"00075100";
        ram_buffer(25605) := X"00189100";
        ram_buffer(25606) := X"004F1021";
        ram_buffer(25607) := X"02831821";
        ram_buffer(25608) := X"000528C0";
        ram_buffer(25609) := X"8FB40000";
        ram_buffer(25610) := X"02649823";
        ram_buffer(25611) := X"02569023";
        ram_buffer(25612) := X"001721C0";
        ram_buffer(25613) := X"00AB2821";
        ram_buffer(25614) := X"00791823";
        ram_buffer(25615) := X"00176100";
        ram_buffer(25616) := X"01473823";
        ram_buffer(25617) := X"0015B080";
        ram_buffer(25618) := X"00095180";
        ram_buffer(25619) := X"00021080";
        ram_buffer(25620) := X"001EF080";
        ram_buffer(25621) := X"01846021";
        ram_buffer(25622) := X"02B6A821";
        ram_buffer(25623) := X"029EF021";
        ram_buffer(25624) := X"012A4821";
        ram_buffer(25625) := X"004F7821";
        ram_buffer(25626) := X"00055140";
        ram_buffer(25627) := X"8FA20008";
        ram_buffer(25628) := X"00032840";
        ram_buffer(25629) := X"001320C0";
        ram_buffer(25630) := X"8FA3000C";
        ram_buffer(25631) := X"00F13821";
        ram_buffer(25632) := X"0012A280";
        ram_buffer(25633) := X"00D5A823";
        ram_buffer(25634) := X"0008B140";
        ram_buffer(25635) := X"00932023";
        ram_buffer(25636) := X"00073940";
        ram_buffer(25637) := X"02549021";
        ram_buffer(25638) := X"0043C821";
        ram_buffer(25639) := X"00F13821";
        ram_buffer(25640) := X"00902023";
        ram_buffer(25641) := X"00001012";
        ram_buffer(25642) := X"01976023";
        ram_buffer(25643) := X"8FA60004";
        ram_buffer(25644) := X"001EF080";
        ram_buffer(25645) := X"02C84023";
        ram_buffer(25646) := X"0015A880";
        ram_buffer(25647) := X"02589023";
        ram_buffer(25648) := X"8FB00010";
        ram_buffer(25649) := X"00F5A821";
        ram_buffer(25650) := X"00094823";
        ram_buffer(25651) := X"03CEF023";
        ram_buffer(25652) := X"000CB940";
        ram_buffer(25653) := X"00084080";
        ram_buffer(25654) := X"0242C021";
        ram_buffer(25655) := X"00D07021";
        ram_buffer(25656) := X"00EF1823";
        ram_buffer(25657) := X"02EC6023";
        ram_buffer(25658) := X"00043040";
        ram_buffer(25659) := X"00A22821";
        ram_buffer(25660) := X"014B5821";
        ram_buffer(25661) := X"03C92021";
        ram_buffer(25662) := X"01094021";
        ram_buffer(25663) := X"03151021";
        ram_buffer(25664) := X"01D93821";
        ram_buffer(25665) := X"00CC3021";
        ram_buffer(25666) := X"00A32821";
        ram_buffer(25667) := X"01D97023";
        ram_buffer(25668) := X"018B6023";
        ram_buffer(25669) := X"00952021";
        ram_buffer(25670) := X"01031821";
        ram_buffer(25671) := X"24424000";
        ram_buffer(25672) := X"000213C3";
        ram_buffer(25673) := X"24E70002";
        ram_buffer(25674) := X"25CE0002";
        ram_buffer(25675) := X"24C64000";
        ram_buffer(25676) := X"258C4000";
        ram_buffer(25677) := X"24A54000";
        ram_buffer(25678) := X"24844000";
        ram_buffer(25679) := X"24634000";
        ram_buffer(25680) := X"ADA20020";
        ram_buffer(25681) := X"00073883";
        ram_buffer(25682) := X"000E7083";
        ram_buffer(25683) := X"000633C3";
        ram_buffer(25684) := X"000C63C3";
        ram_buffer(25685) := X"00052BC3";
        ram_buffer(25686) := X"000423C3";
        ram_buffer(25687) := X"00031BC3";
        ram_buffer(25688) := X"8FA20014";
        ram_buffer(25689) := X"ADA70000";
        ram_buffer(25690) := X"ADAE0080";
        ram_buffer(25691) := X"ADA60040";
        ram_buffer(25692) := X"ADAC00C0";
        ram_buffer(25693) := X"ADA500E0";
        ram_buffer(25694) := X"ADA400A0";
        ram_buffer(25695) := X"ADA30060";
        ram_buffer(25696) := X"25AD0004";
        ram_buffer(25697) := X"15A2FF57";
        ram_buffer(25698) := X"00000000";
        ram_buffer(25699) := X"8FBE003C";
        ram_buffer(25700) := X"8FB70038";
        ram_buffer(25701) := X"8FB60034";
        ram_buffer(25702) := X"8FB50030";
        ram_buffer(25703) := X"8FB4002C";
        ram_buffer(25704) := X"8FB30028";
        ram_buffer(25705) := X"8FB20024";
        ram_buffer(25706) := X"8FB10020";
        ram_buffer(25707) := X"8FB0001C";
        ram_buffer(25708) := X"03E00008";
        ram_buffer(25709) := X"27BD0040";
        ram_buffer(25710) := X"8C820004";
        ram_buffer(25711) := X"27BDFFE8";
        ram_buffer(25712) := X"8C420024";
        ram_buffer(25713) := X"24050001";
        ram_buffer(25714) := X"AFB00010";
        ram_buffer(25715) := X"AFBF0014";
        ram_buffer(25716) := X"0040F809";
        ram_buffer(25717) := X"00808021";
        ram_buffer(25718) := X"8E02000C";
        ram_buffer(25719) := X"00000000";
        ram_buffer(25720) := X"14400006";
        ram_buffer(25721) := X"24020064";
        ram_buffer(25722) := X"8FBF0014";
        ram_buffer(25723) := X"AE020010";
        ram_buffer(25724) := X"8FB00010";
        ram_buffer(25725) := X"03E00008";
        ram_buffer(25726) := X"27BD0018";
        ram_buffer(25727) := X"8FBF0014";
        ram_buffer(25728) := X"240200C8";
        ram_buffer(25729) := X"AE020010";
        ram_buffer(25730) := X"8FB00010";
        ram_buffer(25731) := X"03E00008";
        ram_buffer(25732) := X"27BD0018";
        ram_buffer(25733) := X"8C820004";
        ram_buffer(25734) := X"27BDFFE8";
        ram_buffer(25735) := X"AFB00010";
        ram_buffer(25736) := X"AFBF0014";
        ram_buffer(25737) := X"10400005";
        ram_buffer(25738) := X"00808021";
        ram_buffer(25739) := X"8C420028";
        ram_buffer(25740) := X"00000000";
        ram_buffer(25741) := X"0040F809";
        ram_buffer(25742) := X"00000000";
        ram_buffer(25743) := X"8FBF0014";
        ram_buffer(25744) := X"AE000004";
        ram_buffer(25745) := X"AE000010";
        ram_buffer(25746) := X"8FB00010";
        ram_buffer(25747) := X"03E00008";
        ram_buffer(25748) := X"27BD0018";
        ram_buffer(25749) := X"8C820004";
        ram_buffer(25750) := X"27BDFFE8";
        ram_buffer(25751) := X"8C420000";
        ram_buffer(25752) := X"24060084";
        ram_buffer(25753) := X"AFBF0014";
        ram_buffer(25754) := X"0040F809";
        ram_buffer(25755) := X"00002821";
        ram_buffer(25756) := X"8FBF0014";
        ram_buffer(25757) := X"AC400080";
        ram_buffer(25758) := X"03E00008";
        ram_buffer(25759) := X"27BD0018";
        ram_buffer(25760) := X"8C820004";
        ram_buffer(25761) := X"27BDFFE8";
        ram_buffer(25762) := X"8C420000";
        ram_buffer(25763) := X"24060118";
        ram_buffer(25764) := X"AFBF0014";
        ram_buffer(25765) := X"0040F809";
        ram_buffer(25766) := X"00002821";
        ram_buffer(25767) := X"8FBF0014";
        ram_buffer(25768) := X"AC400114";
        ram_buffer(25769) := X"03E00008";
        ram_buffer(25770) := X"27BD0018";
        ram_buffer(25771) := X"00852021";
        ram_buffer(25772) := X"2482FFFF";
        ram_buffer(25773) := X"14A00002";
        ram_buffer(25774) := X"0045001A";
        ram_buffer(25775) := X"0007000D";
        ram_buffer(25776) := X"00001012";
        ram_buffer(25777) := X"03E00008";
        ram_buffer(25778) := X"00000000";
        ram_buffer(25779) := X"24A3FFFF";
        ram_buffer(25780) := X"00642021";
        ram_buffer(25781) := X"14A00002";
        ram_buffer(25782) := X"0085001A";
        ram_buffer(25783) := X"0007000D";
        ram_buffer(25784) := X"00001010";
        ram_buffer(25785) := X"03E00008";
        ram_buffer(25786) := X"00821023";
        ram_buffer(25787) := X"27BDFFD8";
        ram_buffer(25788) := X"AFB2001C";
        ram_buffer(25789) := X"8FB20038";
        ram_buffer(25790) := X"00052880";
        ram_buffer(25791) := X"00073880";
        ram_buffer(25792) := X"AFB30020";
        ram_buffer(25793) := X"AFB10018";
        ram_buffer(25794) := X"AFB00014";
        ram_buffer(25795) := X"AFBF0024";
        ram_buffer(25796) := X"8FB3003C";
        ram_buffer(25797) := X"00858821";
        ram_buffer(25798) := X"1A40000A";
        ram_buffer(25799) := X"00C78021";
        ram_buffer(25800) := X"26310004";
        ram_buffer(25801) := X"26100004";
        ram_buffer(25802) := X"8E25FFFC";
        ram_buffer(25803) := X"8E04FFFC";
        ram_buffer(25804) := X"2652FFFF";
        ram_buffer(25805) := X"0C027F93";
        ram_buffer(25806) := X"02603021";
        ram_buffer(25807) := X"1640FFF9";
        ram_buffer(25808) := X"26310004";
        ram_buffer(25809) := X"8FBF0024";
        ram_buffer(25810) := X"8FB30020";
        ram_buffer(25811) := X"8FB2001C";
        ram_buffer(25812) := X"8FB10018";
        ram_buffer(25813) := X"8FB00014";
        ram_buffer(25814) := X"03E00008";
        ram_buffer(25815) := X"27BD0028";
        ram_buffer(25816) := X"00A01021";
        ram_buffer(25817) := X"000631C0";
        ram_buffer(25818) := X"00802821";
        ram_buffer(25819) := X"08027F93";
        ram_buffer(25820) := X"00402021";
        ram_buffer(25821) := X"00A03021";
        ram_buffer(25822) := X"0802801D";
        ram_buffer(25823) := X"00002821";
        ram_buffer(25824) := X"27BDFFE8";
        ram_buffer(25825) := X"AFB00010";
        ram_buffer(25826) := X"AFBF0014";
        ram_buffer(25827) := X"8C900000";
        ram_buffer(25828) := X"04A0000F";
        ram_buffer(25829) := X"00000000";
        ram_buffer(25830) := X"8E020068";
        ram_buffer(25831) := X"00000000";
        ram_buffer(25832) := X"0045282A";
        ram_buffer(25833) := X"10A00005";
        ram_buffer(25834) := X"00000000";
        ram_buffer(25835) := X"8FBF0014";
        ram_buffer(25836) := X"8FB00010";
        ram_buffer(25837) := X"03E00008";
        ram_buffer(25838) := X"27BD0018";
        ram_buffer(25839) := X"8E190008";
        ram_buffer(25840) := X"8FBF0014";
        ram_buffer(25841) := X"8FB00010";
        ram_buffer(25842) := X"03200008";
        ram_buffer(25843) := X"27BD0018";
        ram_buffer(25844) := X"8E03006C";
        ram_buffer(25845) := X"00000000";
        ram_buffer(25846) := X"10600006";
        ram_buffer(25847) := X"00801021";
        ram_buffer(25848) := X"8E040068";
        ram_buffer(25849) := X"00000000";
        ram_buffer(25850) := X"28840003";
        ram_buffer(25851) := X"14800007";
        ram_buffer(25852) := X"00000000";
        ram_buffer(25853) := X"00402021";
        ram_buffer(25854) := X"8E020008";
        ram_buffer(25855) := X"00000000";
        ram_buffer(25856) := X"0040F809";
        ram_buffer(25857) := X"00000000";
        ram_buffer(25858) := X"8E03006C";
        ram_buffer(25859) := X"8FBF0014";
        ram_buffer(25860) := X"24630001";
        ram_buffer(25861) := X"AE03006C";
        ram_buffer(25862) := X"8FB00010";
        ram_buffer(25863) := X"03E00008";
        ram_buffer(25864) := X"27BD0018";
        ram_buffer(25865) := X"8C820000";
        ram_buffer(25866) := X"00000000";
        ram_buffer(25867) := X"AC40006C";
        ram_buffer(25868) := X"03E00008";
        ram_buffer(25869) := X"AC400014";
        ram_buffer(25870) := X"8C880000";
        ram_buffer(25871) := X"27BDFFD0";
        ram_buffer(25872) := X"8D020014";
        ram_buffer(25873) := X"00A02021";
        ram_buffer(25874) := X"18400006";
        ram_buffer(25875) := X"AFBF002C";
        ram_buffer(25876) := X"8D030074";
        ram_buffer(25877) := X"00000000";
        ram_buffer(25878) := X"0062182A";
        ram_buffer(25879) := X"10600037";
        ram_buffer(25880) := X"00022880";
        ram_buffer(25881) := X"8D050078";
        ram_buffer(25882) := X"00000000";
        ram_buffer(25883) := X"10A00043";
        ram_buffer(25884) := X"00000000";
        ram_buffer(25885) := X"8D03007C";
        ram_buffer(25886) := X"00000000";
        ram_buffer(25887) := X"0043302A";
        ram_buffer(25888) := X"14C0003E";
        ram_buffer(25889) := X"00000000";
        ram_buffer(25890) := X"8D060080";
        ram_buffer(25891) := X"00000000";
        ram_buffer(25892) := X"00C2302A";
        ram_buffer(25893) := X"14C00039";
        ram_buffer(25894) := X"00431823";
        ram_buffer(25895) := X"00031880";
        ram_buffer(25896) := X"00A31821";
        ram_buffer(25897) := X"8C650000";
        ram_buffer(25898) := X"00000000";
        ram_buffer(25899) := X"10A00033";
        ram_buffer(25900) := X"00000000";
        ram_buffer(25901) := X"00A03021";
        ram_buffer(25902) := X"10000004";
        ram_buffer(25903) := X"24070025";
        ram_buffer(25904) := X"10470027";
        ram_buffer(25905) := X"24020073";
        ram_buffer(25906) := X"00603021";
        ram_buffer(25907) := X"24C30001";
        ram_buffer(25908) := X"8062FFFF";
        ram_buffer(25909) := X"00000000";
        ram_buffer(25910) := X"1440FFF9";
        ram_buffer(25911) := X"00000000";
        ram_buffer(25912) := X"8D020034";
        ram_buffer(25913) := X"8D07001C";
        ram_buffer(25914) := X"8D060018";
        ram_buffer(25915) := X"AFA20024";
        ram_buffer(25916) := X"8D020030";
        ram_buffer(25917) := X"00000000";
        ram_buffer(25918) := X"AFA20020";
        ram_buffer(25919) := X"8D02002C";
        ram_buffer(25920) := X"00000000";
        ram_buffer(25921) := X"AFA2001C";
        ram_buffer(25922) := X"8D020028";
        ram_buffer(25923) := X"00000000";
        ram_buffer(25924) := X"AFA20018";
        ram_buffer(25925) := X"8D020024";
        ram_buffer(25926) := X"00000000";
        ram_buffer(25927) := X"AFA20014";
        ram_buffer(25928) := X"8D020020";
        ram_buffer(25929) := X"0C0283DB";
        ram_buffer(25930) := X"AFA20010";
        ram_buffer(25931) := X"8FBF002C";
        ram_buffer(25932) := X"00000000";
        ram_buffer(25933) := X"03E00008";
        ram_buffer(25934) := X"27BD0030";
        ram_buffer(25935) := X"8D030070";
        ram_buffer(25936) := X"00000000";
        ram_buffer(25937) := X"00651821";
        ram_buffer(25938) := X"8C650000";
        ram_buffer(25939) := X"00000000";
        ram_buffer(25940) := X"14A0FFD8";
        ram_buffer(25941) := X"00000000";
        ram_buffer(25942) := X"10000008";
        ram_buffer(25943) := X"00000000";
        ram_buffer(25944) := X"80C30001";
        ram_buffer(25945) := X"00000000";
        ram_buffer(25946) := X"1462FFDD";
        ram_buffer(25947) := X"25060018";
        ram_buffer(25948) := X"8FBF002C";
        ram_buffer(25949) := X"080283DB";
        ram_buffer(25950) := X"27BD0030";
        ram_buffer(25951) := X"8D030070";
        ram_buffer(25952) := X"AD020018";
        ram_buffer(25953) := X"8C650000";
        ram_buffer(25954) := X"1000FFCB";
        ram_buffer(25955) := X"00A03021";
        ram_buffer(25956) := X"8C820000";
        ram_buffer(25957) := X"27BDFF20";
        ram_buffer(25958) := X"8C42000C";
        ram_buffer(25959) := X"AFBF00DC";
        ram_buffer(25960) := X"0040F809";
        ram_buffer(25961) := X"27A50010";
        ram_buffer(25962) := X"8F828098";
        ram_buffer(25963) := X"3C05100D";
        ram_buffer(25964) := X"8C44000C";
        ram_buffer(25965) := X"27A60010";
        ram_buffer(25966) := X"0C027196";
        ram_buffer(25967) := X"24A5B410";
        ram_buffer(25968) := X"8FBF00DC";
        ram_buffer(25969) := X"00000000";
        ram_buffer(25970) := X"03E00008";
        ram_buffer(25971) := X"27BD00E0";
        ram_buffer(25972) := X"8C820000";
        ram_buffer(25973) := X"27BDFFE8";
        ram_buffer(25974) := X"8C420008";
        ram_buffer(25975) := X"AFBF0014";
        ram_buffer(25976) := X"AFB00010";
        ram_buffer(25977) := X"0040F809";
        ram_buffer(25978) := X"00808021";
        ram_buffer(25979) := X"0C026485";
        ram_buffer(25980) := X"02002021";
        ram_buffer(25981) := X"0C026D37";
        ram_buffer(25982) := X"24040001";
        ram_buffer(25983) := X"3C03100A";
        ram_buffer(25984) := X"246395D0";
        ram_buffer(25985) := X"AC830000";
        ram_buffer(25986) := X"3C03100A";
        ram_buffer(25987) := X"24639380";
        ram_buffer(25988) := X"AC830004";
        ram_buffer(25989) := X"3C03100A";
        ram_buffer(25990) := X"24639590";
        ram_buffer(25991) := X"AC830008";
        ram_buffer(25992) := X"3C03100A";
        ram_buffer(25993) := X"24639438";
        ram_buffer(25994) := X"AC83000C";
        ram_buffer(25995) := X"3C03100A";
        ram_buffer(25996) := X"24639424";
        ram_buffer(25997) := X"AC830010";
        ram_buffer(25998) := X"3C03100D";
        ram_buffer(25999) := X"24639C00";
        ram_buffer(26000) := X"AC830070";
        ram_buffer(26001) := X"24030077";
        ram_buffer(26002) := X"00801021";
        ram_buffer(26003) := X"AC800068";
        ram_buffer(26004) := X"AC80006C";
        ram_buffer(26005) := X"AC800014";
        ram_buffer(26006) := X"AC830074";
        ram_buffer(26007) := X"AC800078";
        ram_buffer(26008) := X"AC80007C";
        ram_buffer(26009) := X"03E00008";
        ram_buffer(26010) := X"AC800080";
        ram_buffer(26011) := X"3C023B9A";
        ram_buffer(26012) := X"3442C9F1";
        ram_buffer(26013) := X"27BDFFC8";
        ram_buffer(26014) := X"00C2102B";
        ram_buffer(26015) := X"AFBE0030";
        ram_buffer(26016) := X"AFB3001C";
        ram_buffer(26017) := X"AFB20018";
        ram_buffer(26018) := X"AFB00010";
        ram_buffer(26019) := X"AFBF0034";
        ram_buffer(26020) := X"AFB7002C";
        ram_buffer(26021) := X"AFB60028";
        ram_buffer(26022) := X"AFB50024";
        ram_buffer(26023) := X"AFB40020";
        ram_buffer(26024) := X"AFB10014";
        ram_buffer(26025) := X"00C09021";
        ram_buffer(26026) := X"0080F021";
        ram_buffer(26027) := X"8C930004";
        ram_buffer(26028) := X"10400069";
        ram_buffer(26029) := X"00A08021";
        ram_buffer(26030) := X"32420007";
        ram_buffer(26031) := X"10400002";
        ram_buffer(26032) := X"26430008";
        ram_buffer(26033) := X"00629023";
        ram_buffer(26034) := X"2E020002";
        ram_buffer(26035) := X"1440000A";
        ram_buffer(26036) := X"00000000";
        ram_buffer(26037) := X"8FC20000";
        ram_buffer(26038) := X"2404000C";
        ram_buffer(26039) := X"AC500018";
        ram_buffer(26040) := X"8FC30000";
        ram_buffer(26041) := X"AC440014";
        ram_buffer(26042) := X"8C620000";
        ram_buffer(26043) := X"00000000";
        ram_buffer(26044) := X"0040F809";
        ram_buffer(26045) := X"03C02021";
        ram_buffer(26046) := X"00108080";
        ram_buffer(26047) := X"0270A021";
        ram_buffer(26048) := X"8E910030";
        ram_buffer(26049) := X"00000000";
        ram_buffer(26050) := X"12200064";
        ram_buffer(26051) := X"27828088";
        ram_buffer(26052) := X"8E230008";
        ram_buffer(26053) := X"00000000";
        ram_buffer(26054) := X"0072102B";
        ram_buffer(26055) := X"14400008";
        ram_buffer(26056) := X"02201021";
        ram_buffer(26057) := X"10000061";
        ram_buffer(26058) := X"00000000";
        ram_buffer(26059) := X"8C430008";
        ram_buffer(26060) := X"00000000";
        ram_buffer(26061) := X"0072202B";
        ram_buffer(26062) := X"10800033";
        ram_buffer(26063) := X"00408821";
        ram_buffer(26064) := X"8E220000";
        ram_buffer(26065) := X"00000000";
        ram_buffer(26066) := X"1440FFF8";
        ram_buffer(26067) := X"26550010";
        ram_buffer(26068) := X"27828080";
        ram_buffer(26069) := X"00508021";
        ram_buffer(26070) := X"8E100000";
        ram_buffer(26071) := X"3C023B9A";
        ram_buffer(26072) := X"3442CA00";
        ram_buffer(26073) := X"00551023";
        ram_buffer(26074) := X"0050182B";
        ram_buffer(26075) := X"14600045";
        ram_buffer(26076) := X"00000000";
        ram_buffer(26077) := X"24170035";
        ram_buffer(26078) := X"0215B021";
        ram_buffer(26079) := X"02C02821";
        ram_buffer(26080) := X"0C026D23";
        ram_buffer(26081) := X"03C02021";
        ram_buffer(26082) := X"14400013";
        ram_buffer(26083) := X"00000000";
        ram_buffer(26084) := X"00108042";
        ram_buffer(26085) := X"2E020032";
        ram_buffer(26086) := X"1040FFF7";
        ram_buffer(26087) := X"24030002";
        ram_buffer(26088) := X"8FC20000";
        ram_buffer(26089) := X"00000000";
        ram_buffer(26090) := X"AC430018";
        ram_buffer(26091) := X"8FC30000";
        ram_buffer(26092) := X"AC570014";
        ram_buffer(26093) := X"8C620000";
        ram_buffer(26094) := X"03C02021";
        ram_buffer(26095) := X"0040F809";
        ram_buffer(26096) := X"0215B021";
        ram_buffer(26097) := X"02C02821";
        ram_buffer(26098) := X"0C026D23";
        ram_buffer(26099) := X"03C02021";
        ram_buffer(26100) := X"1040FFEF";
        ram_buffer(26101) := X"00000000";
        ram_buffer(26102) := X"8E640048";
        ram_buffer(26103) := X"02501821";
        ram_buffer(26104) := X"00963021";
        ram_buffer(26105) := X"AE660048";
        ram_buffer(26106) := X"AC400000";
        ram_buffer(26107) := X"AC400004";
        ram_buffer(26108) := X"12200026";
        ram_buffer(26109) := X"AC430008";
        ram_buffer(26110) := X"AE220000";
        ram_buffer(26111) := X"24050010";
        ram_buffer(26112) := X"10000004";
        ram_buffer(26113) := X"00002021";
        ram_buffer(26114) := X"8C440004";
        ram_buffer(26115) := X"00000000";
        ram_buffer(26116) := X"24850010";
        ram_buffer(26117) := X"02442021";
        ram_buffer(26118) := X"00721823";
        ram_buffer(26119) := X"AC440004";
        ram_buffer(26120) := X"AC430008";
        ram_buffer(26121) := X"8FBF0034";
        ram_buffer(26122) := X"8FBE0030";
        ram_buffer(26123) := X"8FB7002C";
        ram_buffer(26124) := X"8FB60028";
        ram_buffer(26125) := X"8FB50024";
        ram_buffer(26126) := X"8FB40020";
        ram_buffer(26127) := X"8FB3001C";
        ram_buffer(26128) := X"8FB20018";
        ram_buffer(26129) := X"8FB10014";
        ram_buffer(26130) := X"8FB00010";
        ram_buffer(26131) := X"00451021";
        ram_buffer(26132) := X"03E00008";
        ram_buffer(26133) := X"27BD0038";
        ram_buffer(26134) := X"8C820000";
        ram_buffer(26135) := X"24030001";
        ram_buffer(26136) := X"AC430018";
        ram_buffer(26137) := X"8C830000";
        ram_buffer(26138) := X"24050035";
        ram_buffer(26139) := X"8C630000";
        ram_buffer(26140) := X"00000000";
        ram_buffer(26141) := X"0060F809";
        ram_buffer(26142) := X"AC450014";
        ram_buffer(26143) := X"1000FF8F";
        ram_buffer(26144) := X"32420007";
        ram_buffer(26145) := X"1000FFBB";
        ram_buffer(26146) := X"00408021";
        ram_buffer(26147) := X"AE820030";
        ram_buffer(26148) := X"24050010";
        ram_buffer(26149) := X"1000FFDF";
        ram_buffer(26150) := X"00002021";
        ram_buffer(26151) := X"00508021";
        ram_buffer(26152) := X"8E100000";
        ram_buffer(26153) := X"1000FFAD";
        ram_buffer(26154) := X"26550010";
        ram_buffer(26155) := X"8E240004";
        ram_buffer(26156) := X"1000FFD8";
        ram_buffer(26157) := X"24850010";
        ram_buffer(26158) := X"27BDFFD8";
        ram_buffer(26159) := X"2CA20002";
        ram_buffer(26160) := X"AFB40020";
        ram_buffer(26161) := X"AFB3001C";
        ram_buffer(26162) := X"AFB20018";
        ram_buffer(26163) := X"AFBF0024";
        ram_buffer(26164) := X"AFB10014";
        ram_buffer(26165) := X"AFB00010";
        ram_buffer(26166) := X"00A0A021";
        ram_buffer(26167) := X"8C930004";
        ram_buffer(26168) := X"14400039";
        ram_buffer(26169) := X"00809021";
        ram_buffer(26170) := X"8C820000";
        ram_buffer(26171) := X"00000000";
        ram_buffer(26172) := X"AC450018";
        ram_buffer(26173) := X"8C830000";
        ram_buffer(26174) := X"2405000C";
        ram_buffer(26175) := X"AC450014";
        ram_buffer(26176) := X"8C620000";
        ram_buffer(26177) := X"00000000";
        ram_buffer(26178) := X"0040F809";
        ram_buffer(26179) := X"00000000";
        ram_buffer(26180) := X"0014A080";
        ram_buffer(26181) := X"0274A021";
        ram_buffer(26182) := X"8E820038";
        ram_buffer(26183) := X"00000000";
        ram_buffer(26184) := X"1040000F";
        ram_buffer(26185) := X"AE800038";
        ram_buffer(26186) := X"8C430004";
        ram_buffer(26187) := X"8C510008";
        ram_buffer(26188) := X"00402821";
        ram_buffer(26189) := X"00718821";
        ram_buffer(26190) := X"26310010";
        ram_buffer(26191) := X"02203021";
        ram_buffer(26192) := X"8C500000";
        ram_buffer(26193) := X"0C026D29";
        ram_buffer(26194) := X"02402021";
        ram_buffer(26195) := X"8E630048";
        ram_buffer(26196) := X"02001021";
        ram_buffer(26197) := X"00718823";
        ram_buffer(26198) := X"1600FFF3";
        ram_buffer(26199) := X"AE710048";
        ram_buffer(26200) := X"8E820030";
        ram_buffer(26201) := X"00000000";
        ram_buffer(26202) := X"1040000F";
        ram_buffer(26203) := X"AE800030";
        ram_buffer(26204) := X"8C430004";
        ram_buffer(26205) := X"8C510008";
        ram_buffer(26206) := X"00402821";
        ram_buffer(26207) := X"00718821";
        ram_buffer(26208) := X"26310010";
        ram_buffer(26209) := X"02203021";
        ram_buffer(26210) := X"8C500000";
        ram_buffer(26211) := X"0C026D25";
        ram_buffer(26212) := X"02402021";
        ram_buffer(26213) := X"8E630048";
        ram_buffer(26214) := X"02001021";
        ram_buffer(26215) := X"00718823";
        ram_buffer(26216) := X"1600FFF3";
        ram_buffer(26217) := X"AE710048";
        ram_buffer(26218) := X"8FBF0024";
        ram_buffer(26219) := X"8FB40020";
        ram_buffer(26220) := X"8FB3001C";
        ram_buffer(26221) := X"8FB20018";
        ram_buffer(26222) := X"8FB10014";
        ram_buffer(26223) := X"8FB00010";
        ram_buffer(26224) := X"03E00008";
        ram_buffer(26225) := X"27BD0028";
        ram_buffer(26226) := X"24020001";
        ram_buffer(26227) := X"14A2FFD0";
        ram_buffer(26228) := X"00000000";
        ram_buffer(26229) := X"8E700040";
        ram_buffer(26230) := X"00000000";
        ram_buffer(26231) := X"16000007";
        ram_buffer(26232) := X"00000000";
        ram_buffer(26233) := X"10000011";
        ram_buffer(26234) := X"00000000";
        ram_buffer(26235) := X"8E10002C";
        ram_buffer(26236) := X"00000000";
        ram_buffer(26237) := X"1200000D";
        ram_buffer(26238) := X"00000000";
        ram_buffer(26239) := X"8E020028";
        ram_buffer(26240) := X"00000000";
        ram_buffer(26241) := X"1040FFF9";
        ram_buffer(26242) := X"26050030";
        ram_buffer(26243) := X"8E020038";
        ram_buffer(26244) := X"AE000028";
        ram_buffer(26245) := X"0040F809";
        ram_buffer(26246) := X"02402021";
        ram_buffer(26247) := X"8E10002C";
        ram_buffer(26248) := X"00000000";
        ram_buffer(26249) := X"1600FFF5";
        ram_buffer(26250) := X"00000000";
        ram_buffer(26251) := X"8E700044";
        ram_buffer(26252) := X"00000000";
        ram_buffer(26253) := X"16000007";
        ram_buffer(26254) := X"AE600040";
        ram_buffer(26255) := X"1000FFB4";
        ram_buffer(26256) := X"AE600044";
        ram_buffer(26257) := X"8E10002C";
        ram_buffer(26258) := X"00000000";
        ram_buffer(26259) := X"1200000D";
        ram_buffer(26260) := X"00000000";
        ram_buffer(26261) := X"8E020028";
        ram_buffer(26262) := X"00000000";
        ram_buffer(26263) := X"1040FFF9";
        ram_buffer(26264) := X"26050030";
        ram_buffer(26265) := X"8E020038";
        ram_buffer(26266) := X"AE000028";
        ram_buffer(26267) := X"0040F809";
        ram_buffer(26268) := X"02402021";
        ram_buffer(26269) := X"8E10002C";
        ram_buffer(26270) := X"00000000";
        ram_buffer(26271) := X"1600FFF5";
        ram_buffer(26272) := X"00000000";
        ram_buffer(26273) := X"1000FFA2";
        ram_buffer(26274) := X"AE600044";
        ram_buffer(26275) := X"27BDFFE8";
        ram_buffer(26276) := X"24050001";
        ram_buffer(26277) := X"AFB00010";
        ram_buffer(26278) := X"AFBF0014";
        ram_buffer(26279) := X"0C02662E";
        ram_buffer(26280) := X"00808021";
        ram_buffer(26281) := X"02002021";
        ram_buffer(26282) := X"0C02662E";
        ram_buffer(26283) := X"00002821";
        ram_buffer(26284) := X"8E050004";
        ram_buffer(26285) := X"02002021";
        ram_buffer(26286) := X"0C026D25";
        ram_buffer(26287) := X"24060050";
        ram_buffer(26288) := X"AE000004";
        ram_buffer(26289) := X"8FBF0014";
        ram_buffer(26290) := X"02002021";
        ram_buffer(26291) := X"8FB00010";
        ram_buffer(26292) := X"08026D35";
        ram_buffer(26293) := X"27BD0018";
        ram_buffer(26294) := X"3C023B9A";
        ram_buffer(26295) := X"3442C9F1";
        ram_buffer(26296) := X"27BDFFD8";
        ram_buffer(26297) := X"00C2102B";
        ram_buffer(26298) := X"AFB40020";
        ram_buffer(26299) := X"AFB3001C";
        ram_buffer(26300) := X"AFB10014";
        ram_buffer(26301) := X"AFB00010";
        ram_buffer(26302) := X"AFBF0024";
        ram_buffer(26303) := X"AFB20018";
        ram_buffer(26304) := X"00C08021";
        ram_buffer(26305) := X"0080A021";
        ram_buffer(26306) := X"8C910004";
        ram_buffer(26307) := X"1040002B";
        ram_buffer(26308) := X"00A09821";
        ram_buffer(26309) := X"32020007";
        ram_buffer(26310) := X"10400003";
        ram_buffer(26311) := X"00000000";
        ram_buffer(26312) := X"26100008";
        ram_buffer(26313) := X"02028023";
        ram_buffer(26314) := X"2E620002";
        ram_buffer(26315) := X"1440000A";
        ram_buffer(26316) := X"2404000C";
        ram_buffer(26317) := X"8E820000";
        ram_buffer(26318) := X"00000000";
        ram_buffer(26319) := X"AC530018";
        ram_buffer(26320) := X"8E830000";
        ram_buffer(26321) := X"AC440014";
        ram_buffer(26322) := X"8C620000";
        ram_buffer(26323) := X"00000000";
        ram_buffer(26324) := X"0040F809";
        ram_buffer(26325) := X"02802021";
        ram_buffer(26326) := X"26050010";
        ram_buffer(26327) := X"0C026D27";
        ram_buffer(26328) := X"02802021";
        ram_buffer(26329) := X"10400020";
        ram_buffer(26330) := X"00409021";
        ram_buffer(26331) := X"8E220048";
        ram_buffer(26332) := X"00139880";
        ram_buffer(26333) := X"24420010";
        ram_buffer(26334) := X"00501021";
        ram_buffer(26335) := X"AE220048";
        ram_buffer(26336) := X"02338821";
        ram_buffer(26337) := X"8E230038";
        ram_buffer(26338) := X"AE500004";
        ram_buffer(26339) := X"AE430000";
        ram_buffer(26340) := X"AE400008";
        ram_buffer(26341) := X"8FBF0024";
        ram_buffer(26342) := X"AE320038";
        ram_buffer(26343) := X"26420010";
        ram_buffer(26344) := X"8FB40020";
        ram_buffer(26345) := X"8FB3001C";
        ram_buffer(26346) := X"8FB20018";
        ram_buffer(26347) := X"8FB10014";
        ram_buffer(26348) := X"8FB00010";
        ram_buffer(26349) := X"03E00008";
        ram_buffer(26350) := X"27BD0028";
        ram_buffer(26351) := X"8C820000";
        ram_buffer(26352) := X"24030003";
        ram_buffer(26353) := X"AC430018";
        ram_buffer(26354) := X"8C830000";
        ram_buffer(26355) := X"24050035";
        ram_buffer(26356) := X"8C630000";
        ram_buffer(26357) := X"00000000";
        ram_buffer(26358) := X"0060F809";
        ram_buffer(26359) := X"AC450014";
        ram_buffer(26360) := X"1000FFCD";
        ram_buffer(26361) := X"32020007";
        ram_buffer(26362) := X"8E820000";
        ram_buffer(26363) := X"24030004";
        ram_buffer(26364) := X"AC430018";
        ram_buffer(26365) := X"8E830000";
        ram_buffer(26366) := X"24040035";
        ram_buffer(26367) := X"8C630000";
        ram_buffer(26368) := X"AC440014";
        ram_buffer(26369) := X"0060F809";
        ram_buffer(26370) := X"02802021";
        ram_buffer(26371) := X"1000FFD7";
        ram_buffer(26372) := X"00000000";
        ram_buffer(26373) := X"27BDFFC0";
        ram_buffer(26374) := X"8CA20004";
        ram_buffer(26375) := X"AFB5002C";
        ram_buffer(26376) := X"00C7A821";
        ram_buffer(26377) := X"0055102B";
        ram_buffer(26378) := X"AFB60030";
        ram_buffer(26379) := X"AFB30024";
        ram_buffer(26380) := X"AFB00018";
        ram_buffer(26381) := X"AFBF003C";
        ram_buffer(26382) := X"AFBE0038";
        ram_buffer(26383) := X"AFB70034";
        ram_buffer(26384) := X"AFB40028";
        ram_buffer(26385) := X"AFB20020";
        ram_buffer(26386) := X"AFB1001C";
        ram_buffer(26387) := X"00A08021";
        ram_buffer(26388) := X"00C0B021";
        ram_buffer(26389) := X"14400006";
        ram_buffer(26390) := X"00809821";
        ram_buffer(26391) := X"8CA2000C";
        ram_buffer(26392) := X"00000000";
        ram_buffer(26393) := X"0047382B";
        ram_buffer(26394) := X"10E0009F";
        ram_buffer(26395) := X"00000000";
        ram_buffer(26396) := X"8E620000";
        ram_buffer(26397) := X"24040014";
        ram_buffer(26398) := X"8C430000";
        ram_buffer(26399) := X"AC440014";
        ram_buffer(26400) := X"0060F809";
        ram_buffer(26401) := X"02602021";
        ram_buffer(26402) := X"8E050018";
        ram_buffer(26403) := X"00000000";
        ram_buffer(26404) := X"02C5102B";
        ram_buffer(26405) := X"14400007";
        ram_buffer(26406) := X"00000000";
        ram_buffer(26407) := X"8E020010";
        ram_buffer(26408) := X"00000000";
        ram_buffer(26409) := X"00A21021";
        ram_buffer(26410) := X"0055102B";
        ram_buffer(26411) := X"10400053";
        ram_buffer(26412) := X"00000000";
        ram_buffer(26413) := X"8E020028";
        ram_buffer(26414) := X"00000000";
        ram_buffer(26415) := X"1040009B";
        ram_buffer(26416) := X"00000000";
        ram_buffer(26417) := X"8E120008";
        ram_buffer(26418) := X"8E020024";
        ram_buffer(26419) := X"8E030010";
        ram_buffer(26420) := X"144000A2";
        ram_buffer(26421) := X"001291C0";
        ram_buffer(26422) := X"8E04001C";
        ram_buffer(26423) := X"00B6282B";
        ram_buffer(26424) := X"10A0007D";
        ram_buffer(26425) := X"02A32823";
        ram_buffer(26426) := X"AE160018";
        ram_buffer(26427) := X"02C02821";
        ram_buffer(26428) := X"00B20018";
        ram_buffer(26429) := X"0000B812";
        ram_buffer(26430) := X"18600043";
        ram_buffer(26431) := X"0095102B";
        ram_buffer(26432) := X"8E020014";
        ram_buffer(26433) := X"00000000";
        ram_buffer(26434) := X"0062302A";
        ram_buffer(26435) := X"10C00002";
        ram_buffer(26436) := X"00000000";
        ram_buffer(26437) := X"00601021";
        ram_buffer(26438) := X"00851823";
        ram_buffer(26439) := X"0043302A";
        ram_buffer(26440) := X"10C00002";
        ram_buffer(26441) := X"00000000";
        ram_buffer(26442) := X"00401821";
        ram_buffer(26443) := X"8E020004";
        ram_buffer(26444) := X"00000000";
        ram_buffer(26445) := X"00451023";
        ram_buffer(26446) := X"0062282A";
        ram_buffer(26447) := X"10A00002";
        ram_buffer(26448) := X"00000000";
        ram_buffer(26449) := X"00601021";
        ram_buffer(26450) := X"1840002E";
        ram_buffer(26451) := X"26140030";
        ram_buffer(26452) := X"0000F021";
        ram_buffer(26453) := X"00520018";
        ram_buffer(26454) := X"8E020000";
        ram_buffer(26455) := X"001E1880";
        ram_buffer(26456) := X"00431021";
        ram_buffer(26457) := X"8C460000";
        ram_buffer(26458) := X"8E020030";
        ram_buffer(26459) := X"02E03821";
        ram_buffer(26460) := X"02802821";
        ram_buffer(26461) := X"02602021";
        ram_buffer(26462) := X"00008812";
        ram_buffer(26463) := X"0040F809";
        ram_buffer(26464) := X"AFB10010";
        ram_buffer(26465) := X"8E030014";
        ram_buffer(26466) := X"8E020010";
        ram_buffer(26467) := X"03C3F021";
        ram_buffer(26468) := X"005E2823";
        ram_buffer(26469) := X"03C2102A";
        ram_buffer(26470) := X"0065202A";
        ram_buffer(26471) := X"10400017";
        ram_buffer(26472) := X"02F1B821";
        ram_buffer(26473) := X"10800002";
        ram_buffer(26474) := X"00000000";
        ram_buffer(26475) := X"00602821";
        ram_buffer(26476) := X"8E020018";
        ram_buffer(26477) := X"8E04001C";
        ram_buffer(26478) := X"03C21821";
        ram_buffer(26479) := X"00833023";
        ram_buffer(26480) := X"00A6102A";
        ram_buffer(26481) := X"10400002";
        ram_buffer(26482) := X"00000000";
        ram_buffer(26483) := X"00A03021";
        ram_buffer(26484) := X"8E020004";
        ram_buffer(26485) := X"00000000";
        ram_buffer(26486) := X"00431023";
        ram_buffer(26487) := X"00C2182A";
        ram_buffer(26488) := X"10600002";
        ram_buffer(26489) := X"00000000";
        ram_buffer(26490) := X"00C01021";
        ram_buffer(26491) := X"1C40FFDA";
        ram_buffer(26492) := X"00520018";
        ram_buffer(26493) := X"10000004";
        ram_buffer(26494) := X"0095102B";
        ram_buffer(26495) := X"8E04001C";
        ram_buffer(26496) := X"00000000";
        ram_buffer(26497) := X"0095102B";
        ram_buffer(26498) := X"1040001D";
        ram_buffer(26499) := X"0096102B";
        ram_buffer(26500) := X"1040003B";
        ram_buffer(26501) := X"00000000";
        ram_buffer(26502) := X"8FA20050";
        ram_buffer(26503) := X"00000000";
        ram_buffer(26504) := X"144000AD";
        ram_buffer(26505) := X"24040014";
        ram_buffer(26506) := X"02C02021";
        ram_buffer(26507) := X"8E020020";
        ram_buffer(26508) := X"00000000";
        ram_buffer(26509) := X"104000B0";
        ram_buffer(26510) := X"00000000";
        ram_buffer(26511) := X"8E020018";
        ram_buffer(26512) := X"8E130008";
        ram_buffer(26513) := X"00828823";
        ram_buffer(26514) := X"02A2A823";
        ram_buffer(26515) := X"0235182B";
        ram_buffer(26516) := X"1060000C";
        ram_buffer(26517) := X"001399C0";
        ram_buffer(26518) := X"00119080";
        ram_buffer(26519) := X"8E020000";
        ram_buffer(26520) := X"02602821";
        ram_buffer(26521) := X"00521021";
        ram_buffer(26522) := X"8C440000";
        ram_buffer(26523) := X"0C0264DD";
        ram_buffer(26524) := X"26310001";
        ram_buffer(26525) := X"0235102B";
        ram_buffer(26526) := X"1440FFF8";
        ram_buffer(26527) := X"26520004";
        ram_buffer(26528) := X"8E020018";
        ram_buffer(26529) := X"8FA30050";
        ram_buffer(26530) := X"00000000";
        ram_buffer(26531) := X"10600002";
        ram_buffer(26532) := X"24030001";
        ram_buffer(26533) := X"AE030024";
        ram_buffer(26534) := X"02C2B023";
        ram_buffer(26535) := X"8FBF003C";
        ram_buffer(26536) := X"8E020000";
        ram_buffer(26537) := X"0016B080";
        ram_buffer(26538) := X"00561021";
        ram_buffer(26539) := X"8FBE0038";
        ram_buffer(26540) := X"8FB70034";
        ram_buffer(26541) := X"8FB60030";
        ram_buffer(26542) := X"8FB5002C";
        ram_buffer(26543) := X"8FB40028";
        ram_buffer(26544) := X"8FB30024";
        ram_buffer(26545) := X"8FB20020";
        ram_buffer(26546) := X"8FB1001C";
        ram_buffer(26547) := X"8FB00018";
        ram_buffer(26548) := X"03E00008";
        ram_buffer(26549) := X"27BD0040";
        ram_buffer(26550) := X"04A0007C";
        ram_buffer(26551) := X"00000000";
        ram_buffer(26552) := X"1000FF83";
        ram_buffer(26553) := X"AE050018";
        ram_buffer(26554) := X"8CA20000";
        ram_buffer(26555) := X"00000000";
        ram_buffer(26556) := X"1440FF65";
        ram_buffer(26557) := X"00000000";
        ram_buffer(26558) := X"1000FF5D";
        ram_buffer(26559) := X"00000000";
        ram_buffer(26560) := X"8FA20050";
        ram_buffer(26561) := X"00000000";
        ram_buffer(26562) := X"1040FFC8";
        ram_buffer(26563) := X"00000000";
        ram_buffer(26564) := X"8E020020";
        ram_buffer(26565) := X"00000000";
        ram_buffer(26566) := X"1440FFC8";
        ram_buffer(26567) := X"AE15001C";
        ram_buffer(26568) := X"8E020018";
        ram_buffer(26569) := X"1000FFDB";
        ram_buffer(26570) := X"24030001";
        ram_buffer(26571) := X"8E620000";
        ram_buffer(26572) := X"24040044";
        ram_buffer(26573) := X"8C430000";
        ram_buffer(26574) := X"AC440014";
        ram_buffer(26575) := X"0060F809";
        ram_buffer(26576) := X"02602021";
        ram_buffer(26577) := X"8E120008";
        ram_buffer(26578) := X"8E020024";
        ram_buffer(26579) := X"8E050018";
        ram_buffer(26580) := X"8E030010";
        ram_buffer(26581) := X"1040FF60";
        ram_buffer(26582) := X"001291C0";
        ram_buffer(26583) := X"02450018";
        ram_buffer(26584) := X"0000B812";
        ram_buffer(26585) := X"18600073";
        ram_buffer(26586) := X"00000000";
        ram_buffer(26587) := X"8E020014";
        ram_buffer(26588) := X"00000000";
        ram_buffer(26589) := X"0062202A";
        ram_buffer(26590) := X"1480004C";
        ram_buffer(26591) := X"00000000";
        ram_buffer(26592) := X"8E04001C";
        ram_buffer(26593) := X"00000000";
        ram_buffer(26594) := X"00853023";
        ram_buffer(26595) := X"0046382A";
        ram_buffer(26596) := X"14E0003D";
        ram_buffer(26597) := X"00000000";
        ram_buffer(26598) := X"8E020004";
        ram_buffer(26599) := X"00000000";
        ram_buffer(26600) := X"00451023";
        ram_buffer(26601) := X"00C2382A";
        ram_buffer(26602) := X"14E00032";
        ram_buffer(26603) := X"00000000";
        ram_buffer(26604) := X"1840002E";
        ram_buffer(26605) := X"00000000";
        ram_buffer(26606) := X"26110030";
        ram_buffer(26607) := X"0000F021";
        ram_buffer(26608) := X"02420018";
        ram_buffer(26609) := X"8E020000";
        ram_buffer(26610) := X"001E1880";
        ram_buffer(26611) := X"00431021";
        ram_buffer(26612) := X"8C460000";
        ram_buffer(26613) := X"8E020034";
        ram_buffer(26614) := X"02E03821";
        ram_buffer(26615) := X"02202821";
        ram_buffer(26616) := X"02602021";
        ram_buffer(26617) := X"0000A012";
        ram_buffer(26618) := X"0040F809";
        ram_buffer(26619) := X"AFB40010";
        ram_buffer(26620) := X"8E020014";
        ram_buffer(26621) := X"8E030010";
        ram_buffer(26622) := X"03C2F021";
        ram_buffer(26623) := X"007E3023";
        ram_buffer(26624) := X"03C3202A";
        ram_buffer(26625) := X"0046282A";
        ram_buffer(26626) := X"10800044";
        ram_buffer(26627) := X"02F4B821";
        ram_buffer(26628) := X"10A00002";
        ram_buffer(26629) := X"00000000";
        ram_buffer(26630) := X"00403021";
        ram_buffer(26631) := X"8E050018";
        ram_buffer(26632) := X"8E04001C";
        ram_buffer(26633) := X"00BE4821";
        ram_buffer(26634) := X"00893823";
        ram_buffer(26635) := X"00C7102A";
        ram_buffer(26636) := X"10400002";
        ram_buffer(26637) := X"00000000";
        ram_buffer(26638) := X"00C03821";
        ram_buffer(26639) := X"8E020004";
        ram_buffer(26640) := X"00000000";
        ram_buffer(26641) := X"00491023";
        ram_buffer(26642) := X"00E2302A";
        ram_buffer(26643) := X"10C00002";
        ram_buffer(26644) := X"00000000";
        ram_buffer(26645) := X"00E01021";
        ram_buffer(26646) := X"1C40FFDA";
        ram_buffer(26647) := X"02420018";
        ram_buffer(26648) := X"8E120008";
        ram_buffer(26649) := X"00000000";
        ram_buffer(26650) := X"001291C0";
        ram_buffer(26651) := X"1000FF1B";
        ram_buffer(26652) := X"AE000024";
        ram_buffer(26653) := X"00C01021";
        ram_buffer(26654) := X"1C40FFD0";
        ram_buffer(26655) := X"26110030";
        ram_buffer(26656) := X"1000FF16";
        ram_buffer(26657) := X"AE000024";
        ram_buffer(26658) := X"00403021";
        ram_buffer(26659) := X"8E020004";
        ram_buffer(26660) := X"00000000";
        ram_buffer(26661) := X"00451023";
        ram_buffer(26662) := X"00C2382A";
        ram_buffer(26663) := X"10E0FFC4";
        ram_buffer(26664) := X"00000000";
        ram_buffer(26665) := X"1000FFF4";
        ram_buffer(26666) := X"00C01021";
        ram_buffer(26667) := X"8E04001C";
        ram_buffer(26668) := X"00601021";
        ram_buffer(26669) := X"00853023";
        ram_buffer(26670) := X"0046382A";
        ram_buffer(26671) := X"10E0FFB6";
        ram_buffer(26672) := X"00000000";
        ram_buffer(26673) := X"1000FFF1";
        ram_buffer(26674) := X"00403021";
        ram_buffer(26675) := X"00002821";
        ram_buffer(26676) := X"1000FF07";
        ram_buffer(26677) := X"AE050018";
        ram_buffer(26678) := X"8E620000";
        ram_buffer(26679) := X"00000000";
        ram_buffer(26680) := X"8C430000";
        ram_buffer(26681) := X"AC440014";
        ram_buffer(26682) := X"0060F809";
        ram_buffer(26683) := X"02602021";
        ram_buffer(26684) := X"1000FF87";
        ram_buffer(26685) := X"02C02021";
        ram_buffer(26686) := X"8E620000";
        ram_buffer(26687) := X"24040014";
        ram_buffer(26688) := X"8C430000";
        ram_buffer(26689) := X"AC440014";
        ram_buffer(26690) := X"0060F809";
        ram_buffer(26691) := X"02602021";
        ram_buffer(26692) := X"8E020018";
        ram_buffer(26693) := X"1000FF61";
        ram_buffer(26694) := X"02C2B023";
        ram_buffer(26695) := X"8E120008";
        ram_buffer(26696) := X"8E050018";
        ram_buffer(26697) := X"8E04001C";
        ram_buffer(26698) := X"001291C0";
        ram_buffer(26699) := X"1000FEEB";
        ram_buffer(26700) := X"AE000024";
        ram_buffer(26701) := X"8E04001C";
        ram_buffer(26702) := X"1000FEE8";
        ram_buffer(26703) := X"AE000024";
        ram_buffer(26704) := X"27BDFFC0";
        ram_buffer(26705) := X"8CA20004";
        ram_buffer(26706) := X"AFB5002C";
        ram_buffer(26707) := X"00C7A821";
        ram_buffer(26708) := X"0055102B";
        ram_buffer(26709) := X"AFB60030";
        ram_buffer(26710) := X"AFB20020";
        ram_buffer(26711) := X"AFB00018";
        ram_buffer(26712) := X"AFBF003C";
        ram_buffer(26713) := X"AFBE0038";
        ram_buffer(26714) := X"AFB70034";
        ram_buffer(26715) := X"AFB40028";
        ram_buffer(26716) := X"AFB30024";
        ram_buffer(26717) := X"AFB1001C";
        ram_buffer(26718) := X"00A08021";
        ram_buffer(26719) := X"00C0B021";
        ram_buffer(26720) := X"14400006";
        ram_buffer(26721) := X"00809021";
        ram_buffer(26722) := X"8CA2000C";
        ram_buffer(26723) := X"00000000";
        ram_buffer(26724) := X"0047382B";
        ram_buffer(26725) := X"10E0009E";
        ram_buffer(26726) := X"00000000";
        ram_buffer(26727) := X"8E420000";
        ram_buffer(26728) := X"24040014";
        ram_buffer(26729) := X"8C430000";
        ram_buffer(26730) := X"AC440014";
        ram_buffer(26731) := X"0060F809";
        ram_buffer(26732) := X"02402021";
        ram_buffer(26733) := X"8E050018";
        ram_buffer(26734) := X"00000000";
        ram_buffer(26735) := X"02C5102B";
        ram_buffer(26736) := X"14400007";
        ram_buffer(26737) := X"00000000";
        ram_buffer(26738) := X"8E020010";
        ram_buffer(26739) := X"00000000";
        ram_buffer(26740) := X"00A21021";
        ram_buffer(26741) := X"0055102B";
        ram_buffer(26742) := X"10400053";
        ram_buffer(26743) := X"00000000";
        ram_buffer(26744) := X"8E020028";
        ram_buffer(26745) := X"00000000";
        ram_buffer(26746) := X"1040009A";
        ram_buffer(26747) := X"00000000";
        ram_buffer(26748) := X"8E020024";
        ram_buffer(26749) := X"8E130008";
        ram_buffer(26750) := X"8E030010";
        ram_buffer(26751) := X"144000A1";
        ram_buffer(26752) := X"02650018";
        ram_buffer(26753) := X"8E04001C";
        ram_buffer(26754) := X"00B6282B";
        ram_buffer(26755) := X"10A0007C";
        ram_buffer(26756) := X"02A32823";
        ram_buffer(26757) := X"AE160018";
        ram_buffer(26758) := X"02C02821";
        ram_buffer(26759) := X"00B30018";
        ram_buffer(26760) := X"0000B812";
        ram_buffer(26761) := X"18600043";
        ram_buffer(26762) := X"0095102B";
        ram_buffer(26763) := X"8E020014";
        ram_buffer(26764) := X"00000000";
        ram_buffer(26765) := X"0062302A";
        ram_buffer(26766) := X"10C00002";
        ram_buffer(26767) := X"00000000";
        ram_buffer(26768) := X"00601021";
        ram_buffer(26769) := X"00851823";
        ram_buffer(26770) := X"0043302A";
        ram_buffer(26771) := X"10C00002";
        ram_buffer(26772) := X"00000000";
        ram_buffer(26773) := X"00401821";
        ram_buffer(26774) := X"8E020004";
        ram_buffer(26775) := X"00000000";
        ram_buffer(26776) := X"00451023";
        ram_buffer(26777) := X"0062282A";
        ram_buffer(26778) := X"10A00002";
        ram_buffer(26779) := X"00000000";
        ram_buffer(26780) := X"00601021";
        ram_buffer(26781) := X"1840002E";
        ram_buffer(26782) := X"26140030";
        ram_buffer(26783) := X"0000F021";
        ram_buffer(26784) := X"00530018";
        ram_buffer(26785) := X"8E020000";
        ram_buffer(26786) := X"001E1880";
        ram_buffer(26787) := X"00431021";
        ram_buffer(26788) := X"8C460000";
        ram_buffer(26789) := X"8E020030";
        ram_buffer(26790) := X"02E03821";
        ram_buffer(26791) := X"02802821";
        ram_buffer(26792) := X"02402021";
        ram_buffer(26793) := X"00008812";
        ram_buffer(26794) := X"0040F809";
        ram_buffer(26795) := X"AFB10010";
        ram_buffer(26796) := X"8E030014";
        ram_buffer(26797) := X"8E020010";
        ram_buffer(26798) := X"03C3F021";
        ram_buffer(26799) := X"005E2823";
        ram_buffer(26800) := X"03C2102A";
        ram_buffer(26801) := X"0065202A";
        ram_buffer(26802) := X"10400017";
        ram_buffer(26803) := X"02F1B821";
        ram_buffer(26804) := X"10800002";
        ram_buffer(26805) := X"00000000";
        ram_buffer(26806) := X"00602821";
        ram_buffer(26807) := X"8E020018";
        ram_buffer(26808) := X"8E04001C";
        ram_buffer(26809) := X"03C21821";
        ram_buffer(26810) := X"00833023";
        ram_buffer(26811) := X"00A6102A";
        ram_buffer(26812) := X"10400002";
        ram_buffer(26813) := X"00000000";
        ram_buffer(26814) := X"00A03021";
        ram_buffer(26815) := X"8E020004";
        ram_buffer(26816) := X"00000000";
        ram_buffer(26817) := X"00431023";
        ram_buffer(26818) := X"00C2182A";
        ram_buffer(26819) := X"10600002";
        ram_buffer(26820) := X"00000000";
        ram_buffer(26821) := X"00C01021";
        ram_buffer(26822) := X"1C40FFDA";
        ram_buffer(26823) := X"00530018";
        ram_buffer(26824) := X"10000004";
        ram_buffer(26825) := X"0095102B";
        ram_buffer(26826) := X"8E04001C";
        ram_buffer(26827) := X"00000000";
        ram_buffer(26828) := X"0095102B";
        ram_buffer(26829) := X"1040001C";
        ram_buffer(26830) := X"0096102B";
        ram_buffer(26831) := X"1040003A";
        ram_buffer(26832) := X"00000000";
        ram_buffer(26833) := X"8FA20050";
        ram_buffer(26834) := X"00000000";
        ram_buffer(26835) := X"144000A9";
        ram_buffer(26836) := X"24040014";
        ram_buffer(26837) := X"02C02021";
        ram_buffer(26838) := X"8E020020";
        ram_buffer(26839) := X"00000000";
        ram_buffer(26840) := X"104000AC";
        ram_buffer(26841) := X"00000000";
        ram_buffer(26842) := X"8E020018";
        ram_buffer(26843) := X"8E120008";
        ram_buffer(26844) := X"00828823";
        ram_buffer(26845) := X"02A2A823";
        ram_buffer(26846) := X"0235182B";
        ram_buffer(26847) := X"1060000B";
        ram_buffer(26848) := X"00119880";
        ram_buffer(26849) := X"8E020000";
        ram_buffer(26850) := X"02402821";
        ram_buffer(26851) := X"00531021";
        ram_buffer(26852) := X"8C440000";
        ram_buffer(26853) := X"0C0264DD";
        ram_buffer(26854) := X"26310001";
        ram_buffer(26855) := X"0235102B";
        ram_buffer(26856) := X"1440FFF8";
        ram_buffer(26857) := X"26730004";
        ram_buffer(26858) := X"8E020018";
        ram_buffer(26859) := X"8FA30050";
        ram_buffer(26860) := X"00000000";
        ram_buffer(26861) := X"10600002";
        ram_buffer(26862) := X"24030001";
        ram_buffer(26863) := X"AE030024";
        ram_buffer(26864) := X"02C2B023";
        ram_buffer(26865) := X"8FBF003C";
        ram_buffer(26866) := X"8E020000";
        ram_buffer(26867) := X"0016B080";
        ram_buffer(26868) := X"00561021";
        ram_buffer(26869) := X"8FBE0038";
        ram_buffer(26870) := X"8FB70034";
        ram_buffer(26871) := X"8FB60030";
        ram_buffer(26872) := X"8FB5002C";
        ram_buffer(26873) := X"8FB40028";
        ram_buffer(26874) := X"8FB30024";
        ram_buffer(26875) := X"8FB20020";
        ram_buffer(26876) := X"8FB1001C";
        ram_buffer(26877) := X"8FB00018";
        ram_buffer(26878) := X"03E00008";
        ram_buffer(26879) := X"27BD0040";
        ram_buffer(26880) := X"04A00079";
        ram_buffer(26881) := X"00000000";
        ram_buffer(26882) := X"1000FF84";
        ram_buffer(26883) := X"AE050018";
        ram_buffer(26884) := X"8CA20000";
        ram_buffer(26885) := X"00000000";
        ram_buffer(26886) := X"1440FF66";
        ram_buffer(26887) := X"00000000";
        ram_buffer(26888) := X"1000FF5E";
        ram_buffer(26889) := X"00000000";
        ram_buffer(26890) := X"8FA20050";
        ram_buffer(26891) := X"00000000";
        ram_buffer(26892) := X"1040FFC9";
        ram_buffer(26893) := X"00000000";
        ram_buffer(26894) := X"8E020020";
        ram_buffer(26895) := X"00000000";
        ram_buffer(26896) := X"1440FFC9";
        ram_buffer(26897) := X"AE15001C";
        ram_buffer(26898) := X"8E020018";
        ram_buffer(26899) := X"1000FFDB";
        ram_buffer(26900) := X"24030001";
        ram_buffer(26901) := X"8E420000";
        ram_buffer(26902) := X"24040044";
        ram_buffer(26903) := X"8C430000";
        ram_buffer(26904) := X"AC440014";
        ram_buffer(26905) := X"0060F809";
        ram_buffer(26906) := X"02402021";
        ram_buffer(26907) := X"8E020024";
        ram_buffer(26908) := X"8E050018";
        ram_buffer(26909) := X"8E130008";
        ram_buffer(26910) := X"8E030010";
        ram_buffer(26911) := X"1040FF61";
        ram_buffer(26912) := X"02650018";
        ram_buffer(26913) := X"0000B812";
        ram_buffer(26914) := X"1860006D";
        ram_buffer(26915) := X"00000000";
        ram_buffer(26916) := X"8E020014";
        ram_buffer(26917) := X"00000000";
        ram_buffer(26918) := X"0062202A";
        ram_buffer(26919) := X"1480004A";
        ram_buffer(26920) := X"00000000";
        ram_buffer(26921) := X"8E04001C";
        ram_buffer(26922) := X"00000000";
        ram_buffer(26923) := X"00853023";
        ram_buffer(26924) := X"0046382A";
        ram_buffer(26925) := X"14E0003B";
        ram_buffer(26926) := X"00000000";
        ram_buffer(26927) := X"8E020004";
        ram_buffer(26928) := X"00000000";
        ram_buffer(26929) := X"00451023";
        ram_buffer(26930) := X"00C2382A";
        ram_buffer(26931) := X"14E00030";
        ram_buffer(26932) := X"00000000";
        ram_buffer(26933) := X"1840002C";
        ram_buffer(26934) := X"00000000";
        ram_buffer(26935) := X"26110030";
        ram_buffer(26936) := X"0000F021";
        ram_buffer(26937) := X"02620018";
        ram_buffer(26938) := X"8E020000";
        ram_buffer(26939) := X"001E1880";
        ram_buffer(26940) := X"00431021";
        ram_buffer(26941) := X"8C460000";
        ram_buffer(26942) := X"8E020034";
        ram_buffer(26943) := X"02E03821";
        ram_buffer(26944) := X"02202821";
        ram_buffer(26945) := X"02402021";
        ram_buffer(26946) := X"0000A012";
        ram_buffer(26947) := X"0040F809";
        ram_buffer(26948) := X"AFB40010";
        ram_buffer(26949) := X"8E020014";
        ram_buffer(26950) := X"8E030010";
        ram_buffer(26951) := X"03C2F021";
        ram_buffer(26952) := X"007E3023";
        ram_buffer(26953) := X"03C3202A";
        ram_buffer(26954) := X"0046282A";
        ram_buffer(26955) := X"10800042";
        ram_buffer(26956) := X"02F4B821";
        ram_buffer(26957) := X"10A00002";
        ram_buffer(26958) := X"00000000";
        ram_buffer(26959) := X"00403021";
        ram_buffer(26960) := X"8E050018";
        ram_buffer(26961) := X"8E04001C";
        ram_buffer(26962) := X"00BE4821";
        ram_buffer(26963) := X"00893823";
        ram_buffer(26964) := X"00C7102A";
        ram_buffer(26965) := X"10400002";
        ram_buffer(26966) := X"00000000";
        ram_buffer(26967) := X"00C03821";
        ram_buffer(26968) := X"8E020004";
        ram_buffer(26969) := X"00000000";
        ram_buffer(26970) := X"00491023";
        ram_buffer(26971) := X"00E2302A";
        ram_buffer(26972) := X"10C00002";
        ram_buffer(26973) := X"00000000";
        ram_buffer(26974) := X"00E01021";
        ram_buffer(26975) := X"1C40FFDA";
        ram_buffer(26976) := X"02620018";
        ram_buffer(26977) := X"8E130008";
        ram_buffer(26978) := X"1000FF1F";
        ram_buffer(26979) := X"AE000024";
        ram_buffer(26980) := X"00C01021";
        ram_buffer(26981) := X"1C40FFD2";
        ram_buffer(26982) := X"26110030";
        ram_buffer(26983) := X"1000FF1A";
        ram_buffer(26984) := X"AE000024";
        ram_buffer(26985) := X"00403021";
        ram_buffer(26986) := X"8E020004";
        ram_buffer(26987) := X"00000000";
        ram_buffer(26988) := X"00451023";
        ram_buffer(26989) := X"00C2382A";
        ram_buffer(26990) := X"10E0FFC6";
        ram_buffer(26991) := X"00000000";
        ram_buffer(26992) := X"1000FFF4";
        ram_buffer(26993) := X"00C01021";
        ram_buffer(26994) := X"8E04001C";
        ram_buffer(26995) := X"00601021";
        ram_buffer(26996) := X"00853023";
        ram_buffer(26997) := X"0046382A";
        ram_buffer(26998) := X"10E0FFB8";
        ram_buffer(26999) := X"00000000";
        ram_buffer(27000) := X"1000FFF1";
        ram_buffer(27001) := X"00403021";
        ram_buffer(27002) := X"00002821";
        ram_buffer(27003) := X"1000FF0B";
        ram_buffer(27004) := X"AE050018";
        ram_buffer(27005) := X"8E420000";
        ram_buffer(27006) := X"00000000";
        ram_buffer(27007) := X"8C430000";
        ram_buffer(27008) := X"AC440014";
        ram_buffer(27009) := X"0060F809";
        ram_buffer(27010) := X"02402021";
        ram_buffer(27011) := X"1000FF8A";
        ram_buffer(27012) := X"02C02021";
        ram_buffer(27013) := X"8E420000";
        ram_buffer(27014) := X"24040014";
        ram_buffer(27015) := X"8C430000";
        ram_buffer(27016) := X"AC440014";
        ram_buffer(27017) := X"0060F809";
        ram_buffer(27018) := X"02402021";
        ram_buffer(27019) := X"8E020018";
        ram_buffer(27020) := X"1000FF64";
        ram_buffer(27021) := X"02C2B023";
        ram_buffer(27022) := X"8E130008";
        ram_buffer(27023) := X"8E050018";
        ram_buffer(27024) := X"8E04001C";
        ram_buffer(27025) := X"1000FEF0";
        ram_buffer(27026) := X"AE000024";
        ram_buffer(27027) := X"27BDFFB8";
        ram_buffer(27028) := X"AFB10024";
        ram_buffer(27029) := X"3C113B9A";
        ram_buffer(27030) := X"3631C9F0";
        ram_buffer(27031) := X"14C00002";
        ram_buffer(27032) := X"0226001B";
        ram_buffer(27033) := X"0007000D";
        ram_buffer(27034) := X"AFB7003C";
        ram_buffer(27035) := X"AFB60038";
        ram_buffer(27036) := X"AFB50034";
        ram_buffer(27037) := X"AFB20028";
        ram_buffer(27038) := X"AFB00020";
        ram_buffer(27039) := X"AFBF0044";
        ram_buffer(27040) := X"AFBE0040";
        ram_buffer(27041) := X"AFB40030";
        ram_buffer(27042) := X"AFB3002C";
        ram_buffer(27043) := X"00C0A821";
        ram_buffer(27044) := X"0080B021";
        ram_buffer(27045) := X"AFA5004C";
        ram_buffer(27046) := X"8C920004";
        ram_buffer(27047) := X"00008812";
        ram_buffer(27048) := X"0000B812";
        ram_buffer(27049) := X"12200075";
        ram_buffer(27050) := X"00E08021";
        ram_buffer(27051) := X"0230882A";
        ram_buffer(27052) := X"16200002";
        ram_buffer(27053) := X"00000000";
        ram_buffer(27054) := X"0200B821";
        ram_buffer(27055) := X"8FA5004C";
        ram_buffer(27056) := X"AE57004C";
        ram_buffer(27057) := X"00103080";
        ram_buffer(27058) := X"0C02659B";
        ram_buffer(27059) := X"02C02021";
        ram_buffer(27060) := X"12000043";
        ram_buffer(27061) := X"00408821";
        ram_buffer(27062) := X"8FA2004C";
        ram_buffer(27063) := X"3C123B9A";
        ram_buffer(27064) := X"2C540002";
        ram_buffer(27065) := X"00021080";
        ram_buffer(27066) := X"AFA20010";
        ram_buffer(27067) := X"3642C9F1";
        ram_buffer(27068) := X"0000F021";
        ram_buffer(27069) := X"AFA20014";
        ram_buffer(27070) := X"021E1023";
        ram_buffer(27071) := X"0057182B";
        ram_buffer(27072) := X"10600003";
        ram_buffer(27073) := X"02B70018";
        ram_buffer(27074) := X"0040B821";
        ram_buffer(27075) := X"02B70018";
        ram_buffer(27076) := X"8FA20014";
        ram_buffer(27077) := X"8ED30004";
        ram_buffer(27078) := X"00009012";
        ram_buffer(27079) := X"0242102B";
        ram_buffer(27080) := X"1040003C";
        ram_buffer(27081) := X"24030003";
        ram_buffer(27082) := X"32420007";
        ram_buffer(27083) := X"10400002";
        ram_buffer(27084) := X"26460008";
        ram_buffer(27085) := X"00C29023";
        ram_buffer(27086) := X"1680000B";
        ram_buffer(27087) := X"2405000C";
        ram_buffer(27088) := X"8EC20000";
        ram_buffer(27089) := X"8FA3004C";
        ram_buffer(27090) := X"00000000";
        ram_buffer(27091) := X"AC430018";
        ram_buffer(27092) := X"8EC30000";
        ram_buffer(27093) := X"AC450014";
        ram_buffer(27094) := X"8C620000";
        ram_buffer(27095) := X"00000000";
        ram_buffer(27096) := X"0040F809";
        ram_buffer(27097) := X"02C02021";
        ram_buffer(27098) := X"26450010";
        ram_buffer(27099) := X"0C026D27";
        ram_buffer(27100) := X"02C02021";
        ram_buffer(27101) := X"10400033";
        ram_buffer(27102) := X"00000000";
        ram_buffer(27103) := X"8E630048";
        ram_buffer(27104) := X"8FA40010";
        ram_buffer(27105) := X"24630010";
        ram_buffer(27106) := X"00721821";
        ram_buffer(27107) := X"AE630048";
        ram_buffer(27108) := X"02642021";
        ram_buffer(27109) := X"8C850038";
        ram_buffer(27110) := X"24430010";
        ram_buffer(27111) := X"AC450000";
        ram_buffer(27112) := X"AC520004";
        ram_buffer(27113) := X"AC400008";
        ram_buffer(27114) := X"12E0000A";
        ram_buffer(27115) := X"AC820038";
        ram_buffer(27116) := X"001E1080";
        ram_buffer(27117) := X"03D7F021";
        ram_buffer(27118) := X"001E2080";
        ram_buffer(27119) := X"02221021";
        ram_buffer(27120) := X"02242021";
        ram_buffer(27121) := X"AC430000";
        ram_buffer(27122) := X"24420004";
        ram_buffer(27123) := X"1444FFFD";
        ram_buffer(27124) := X"00751821";
        ram_buffer(27125) := X"03D0102B";
        ram_buffer(27126) := X"1440FFC8";
        ram_buffer(27127) := X"021E1023";
        ram_buffer(27128) := X"8FBF0044";
        ram_buffer(27129) := X"02201021";
        ram_buffer(27130) := X"8FBE0040";
        ram_buffer(27131) := X"8FB7003C";
        ram_buffer(27132) := X"8FB60038";
        ram_buffer(27133) := X"8FB50034";
        ram_buffer(27134) := X"8FB40030";
        ram_buffer(27135) := X"8FB3002C";
        ram_buffer(27136) := X"8FB20028";
        ram_buffer(27137) := X"8FB10024";
        ram_buffer(27138) := X"8FB00020";
        ram_buffer(27139) := X"03E00008";
        ram_buffer(27140) := X"27BD0048";
        ram_buffer(27141) := X"8EC20000";
        ram_buffer(27142) := X"00000000";
        ram_buffer(27143) := X"AC430018";
        ram_buffer(27144) := X"8EC30000";
        ram_buffer(27145) := X"24050035";
        ram_buffer(27146) := X"AC450014";
        ram_buffer(27147) := X"8C620000";
        ram_buffer(27148) := X"00000000";
        ram_buffer(27149) := X"0040F809";
        ram_buffer(27150) := X"02C02021";
        ram_buffer(27151) := X"1000FFBB";
        ram_buffer(27152) := X"32420007";
        ram_buffer(27153) := X"8EC30000";
        ram_buffer(27154) := X"AFA20018";
        ram_buffer(27155) := X"24020004";
        ram_buffer(27156) := X"AC620018";
        ram_buffer(27157) := X"8EC50000";
        ram_buffer(27158) := X"24020035";
        ram_buffer(27159) := X"AC620014";
        ram_buffer(27160) := X"8CA30000";
        ram_buffer(27161) := X"00000000";
        ram_buffer(27162) := X"0060F809";
        ram_buffer(27163) := X"02C02021";
        ram_buffer(27164) := X"8FA20018";
        ram_buffer(27165) := X"1000FFC1";
        ram_buffer(27166) := X"00000000";
        ram_buffer(27167) := X"8C820000";
        ram_buffer(27168) := X"24050045";
        ram_buffer(27169) := X"8C430000";
        ram_buffer(27170) := X"00000000";
        ram_buffer(27171) := X"0060F809";
        ram_buffer(27172) := X"AC450014";
        ram_buffer(27173) := X"1000FF86";
        ram_buffer(27174) := X"0230882A";
        ram_buffer(27175) := X"27BDFFB8";
        ram_buffer(27176) := X"AFB10024";
        ram_buffer(27177) := X"3C113B9A";
        ram_buffer(27178) := X"3631C9F0";
        ram_buffer(27179) := X"AFB7003C";
        ram_buffer(27180) := X"0006B9C0";
        ram_buffer(27181) := X"16E00002";
        ram_buffer(27182) := X"0237001B";
        ram_buffer(27183) := X"0007000D";
        ram_buffer(27184) := X"AFB60038";
        ram_buffer(27185) := X"AFB50034";
        ram_buffer(27186) := X"AFB20028";
        ram_buffer(27187) := X"AFB00020";
        ram_buffer(27188) := X"AFBF0044";
        ram_buffer(27189) := X"AFBE0040";
        ram_buffer(27190) := X"AFB40030";
        ram_buffer(27191) := X"AFB3002C";
        ram_buffer(27192) := X"0080A821";
        ram_buffer(27193) := X"AFA5004C";
        ram_buffer(27194) := X"8C920004";
        ram_buffer(27195) := X"00008812";
        ram_buffer(27196) := X"0000B012";
        ram_buffer(27197) := X"12200071";
        ram_buffer(27198) := X"00E08021";
        ram_buffer(27199) := X"0230882A";
        ram_buffer(27200) := X"16200002";
        ram_buffer(27201) := X"00000000";
        ram_buffer(27202) := X"0200B021";
        ram_buffer(27203) := X"8FA5004C";
        ram_buffer(27204) := X"AE56004C";
        ram_buffer(27205) := X"00103080";
        ram_buffer(27206) := X"0C02659B";
        ram_buffer(27207) := X"02A02021";
        ram_buffer(27208) := X"1200003F";
        ram_buffer(27209) := X"00408821";
        ram_buffer(27210) := X"8FA2004C";
        ram_buffer(27211) := X"3C123B9A";
        ram_buffer(27212) := X"2C540002";
        ram_buffer(27213) := X"00021080";
        ram_buffer(27214) := X"AFA20010";
        ram_buffer(27215) := X"3642C9F1";
        ram_buffer(27216) := X"0000F021";
        ram_buffer(27217) := X"AFA20014";
        ram_buffer(27218) := X"021E1023";
        ram_buffer(27219) := X"0056182B";
        ram_buffer(27220) := X"10600003";
        ram_buffer(27221) := X"02F60018";
        ram_buffer(27222) := X"0040B021";
        ram_buffer(27223) := X"02F60018";
        ram_buffer(27224) := X"8FA20014";
        ram_buffer(27225) := X"8EB30004";
        ram_buffer(27226) := X"00009012";
        ram_buffer(27227) := X"0242102B";
        ram_buffer(27228) := X"10400038";
        ram_buffer(27229) := X"24030003";
        ram_buffer(27230) := X"1680000B";
        ram_buffer(27231) := X"2405000C";
        ram_buffer(27232) := X"8EA20000";
        ram_buffer(27233) := X"8FA3004C";
        ram_buffer(27234) := X"00000000";
        ram_buffer(27235) := X"AC430018";
        ram_buffer(27236) := X"8EA30000";
        ram_buffer(27237) := X"AC450014";
        ram_buffer(27238) := X"8C620000";
        ram_buffer(27239) := X"00000000";
        ram_buffer(27240) := X"0040F809";
        ram_buffer(27241) := X"02A02021";
        ram_buffer(27242) := X"26450010";
        ram_buffer(27243) := X"0C026D27";
        ram_buffer(27244) := X"02A02021";
        ram_buffer(27245) := X"10400033";
        ram_buffer(27246) := X"00000000";
        ram_buffer(27247) := X"8E630048";
        ram_buffer(27248) := X"8FA40010";
        ram_buffer(27249) := X"24630010";
        ram_buffer(27250) := X"00721821";
        ram_buffer(27251) := X"AE630048";
        ram_buffer(27252) := X"02642021";
        ram_buffer(27253) := X"8C850038";
        ram_buffer(27254) := X"24430010";
        ram_buffer(27255) := X"AC450000";
        ram_buffer(27256) := X"AC520004";
        ram_buffer(27257) := X"AC400008";
        ram_buffer(27258) := X"12C0000A";
        ram_buffer(27259) := X"AC820038";
        ram_buffer(27260) := X"001E1080";
        ram_buffer(27261) := X"03D6F021";
        ram_buffer(27262) := X"001E2080";
        ram_buffer(27263) := X"02221021";
        ram_buffer(27264) := X"02242021";
        ram_buffer(27265) := X"AC430000";
        ram_buffer(27266) := X"24420004";
        ram_buffer(27267) := X"1444FFFD";
        ram_buffer(27268) := X"00771821";
        ram_buffer(27269) := X"03D0102B";
        ram_buffer(27270) := X"1440FFCC";
        ram_buffer(27271) := X"021E1023";
        ram_buffer(27272) := X"8FBF0044";
        ram_buffer(27273) := X"02201021";
        ram_buffer(27274) := X"8FBE0040";
        ram_buffer(27275) := X"8FB7003C";
        ram_buffer(27276) := X"8FB60038";
        ram_buffer(27277) := X"8FB50034";
        ram_buffer(27278) := X"8FB40030";
        ram_buffer(27279) := X"8FB3002C";
        ram_buffer(27280) := X"8FB20028";
        ram_buffer(27281) := X"8FB10024";
        ram_buffer(27282) := X"8FB00020";
        ram_buffer(27283) := X"03E00008";
        ram_buffer(27284) := X"27BD0048";
        ram_buffer(27285) := X"8EA20000";
        ram_buffer(27286) := X"00000000";
        ram_buffer(27287) := X"AC430018";
        ram_buffer(27288) := X"8EA30000";
        ram_buffer(27289) := X"24050035";
        ram_buffer(27290) := X"AC450014";
        ram_buffer(27291) := X"8C620000";
        ram_buffer(27292) := X"00000000";
        ram_buffer(27293) := X"0040F809";
        ram_buffer(27294) := X"02A02021";
        ram_buffer(27295) := X"1000FFBE";
        ram_buffer(27296) := X"00000000";
        ram_buffer(27297) := X"8EA30000";
        ram_buffer(27298) := X"AFA20018";
        ram_buffer(27299) := X"24020004";
        ram_buffer(27300) := X"AC620018";
        ram_buffer(27301) := X"8EA50000";
        ram_buffer(27302) := X"24020035";
        ram_buffer(27303) := X"AC620014";
        ram_buffer(27304) := X"8CA30000";
        ram_buffer(27305) := X"00000000";
        ram_buffer(27306) := X"0060F809";
        ram_buffer(27307) := X"02A02021";
        ram_buffer(27308) := X"8FA20018";
        ram_buffer(27309) := X"1000FFC1";
        ram_buffer(27310) := X"00000000";
        ram_buffer(27311) := X"8C820000";
        ram_buffer(27312) := X"24050045";
        ram_buffer(27313) := X"8C430000";
        ram_buffer(27314) := X"00000000";
        ram_buffer(27315) := X"0060F809";
        ram_buffer(27316) := X"AC450014";
        ram_buffer(27317) := X"1000FF8A";
        ram_buffer(27318) := X"0230882A";
        ram_buffer(27319) := X"27BDFFD8";
        ram_buffer(27320) := X"AFB30020";
        ram_buffer(27321) := X"8C930004";
        ram_buffer(27322) := X"AFBF0024";
        ram_buffer(27323) := X"8E620040";
        ram_buffer(27324) := X"AFB2001C";
        ram_buffer(27325) := X"AFB10018";
        ram_buffer(27326) := X"104000B8";
        ram_buffer(27327) := X"AFB00014";
        ram_buffer(27328) := X"00008021";
        ram_buffer(27329) := X"10000005";
        ram_buffer(27330) := X"00008821";
        ram_buffer(27331) := X"8C42002C";
        ram_buffer(27332) := X"00000000";
        ram_buffer(27333) := X"10400011";
        ram_buffer(27334) := X"00000000";
        ram_buffer(27335) := X"8C430000";
        ram_buffer(27336) := X"00000000";
        ram_buffer(27337) := X"1460FFF9";
        ram_buffer(27338) := X"00000000";
        ram_buffer(27339) := X"8C430008";
        ram_buffer(27340) := X"8C45000C";
        ram_buffer(27341) := X"8C460004";
        ram_buffer(27342) := X"00650018";
        ram_buffer(27343) := X"8C42002C";
        ram_buffer(27344) := X"00002812";
        ram_buffer(27345) := X"00B18821";
        ram_buffer(27346) := X"00000000";
        ram_buffer(27347) := X"00660018";
        ram_buffer(27348) := X"00001812";
        ram_buffer(27349) := X"1440FFF1";
        ram_buffer(27350) := X"00708021";
        ram_buffer(27351) := X"8E620044";
        ram_buffer(27352) := X"00000000";
        ram_buffer(27353) := X"14400007";
        ram_buffer(27354) := X"00000000";
        ram_buffer(27355) := X"10000016";
        ram_buffer(27356) := X"00000000";
        ram_buffer(27357) := X"8C42002C";
        ram_buffer(27358) := X"00000000";
        ram_buffer(27359) := X"10400012";
        ram_buffer(27360) := X"00000000";
        ram_buffer(27361) := X"8C430000";
        ram_buffer(27362) := X"00000000";
        ram_buffer(27363) := X"1460FFF9";
        ram_buffer(27364) := X"00000000";
        ram_buffer(27365) := X"8C430008";
        ram_buffer(27366) := X"8C45000C";
        ram_buffer(27367) := X"8C460004";
        ram_buffer(27368) := X"00650018";
        ram_buffer(27369) := X"8C42002C";
        ram_buffer(27370) := X"00002812";
        ram_buffer(27371) := X"000529C0";
        ram_buffer(27372) := X"00B18821";
        ram_buffer(27373) := X"00660018";
        ram_buffer(27374) := X"00001812";
        ram_buffer(27375) := X"000319C0";
        ram_buffer(27376) := X"1440FFF0";
        ram_buffer(27377) := X"00708021";
        ram_buffer(27378) := X"1A20005E";
        ram_buffer(27379) := X"02003021";
        ram_buffer(27380) := X"8E670048";
        ram_buffer(27381) := X"02202821";
        ram_buffer(27382) := X"0C026D2B";
        ram_buffer(27383) := X"00809021";
        ram_buffer(27384) := X"0050802A";
        ram_buffer(27385) := X"1200005E";
        ram_buffer(27386) := X"00000000";
        ram_buffer(27387) := X"16200002";
        ram_buffer(27388) := X"0051001A";
        ram_buffer(27389) := X"0007000D";
        ram_buffer(27390) := X"00008812";
        ram_buffer(27391) := X"1A20007D";
        ram_buffer(27392) := X"00000000";
        ram_buffer(27393) := X"8E700040";
        ram_buffer(27394) := X"00000000";
        ram_buffer(27395) := X"16000007";
        ram_buffer(27396) := X"00000000";
        ram_buffer(27397) := X"10000023";
        ram_buffer(27398) := X"00000000";
        ram_buffer(27399) := X"8E10002C";
        ram_buffer(27400) := X"00000000";
        ram_buffer(27401) := X"1200001F";
        ram_buffer(27402) := X"00000000";
        ram_buffer(27403) := X"8E030000";
        ram_buffer(27404) := X"00000000";
        ram_buffer(27405) := X"1460FFF9";
        ram_buffer(27406) := X"00000000";
        ram_buffer(27407) := X"8E070004";
        ram_buffer(27408) := X"8E03000C";
        ram_buffer(27409) := X"24E2FFFF";
        ram_buffer(27410) := X"14600002";
        ram_buffer(27411) := X"0043001B";
        ram_buffer(27412) := X"0007000D";
        ram_buffer(27413) := X"00001012";
        ram_buffer(27414) := X"24420001";
        ram_buffer(27415) := X"0222102A";
        ram_buffer(27416) := X"14400042";
        ram_buffer(27417) := X"02230018";
        ram_buffer(27418) := X"AE070010";
        ram_buffer(27419) := X"8E060008";
        ram_buffer(27420) := X"24050001";
        ram_buffer(27421) := X"0C026993";
        ram_buffer(27422) := X"02402021";
        ram_buffer(27423) := X"8E63004C";
        ram_buffer(27424) := X"AE020000";
        ram_buffer(27425) := X"AE030014";
        ram_buffer(27426) := X"AE000018";
        ram_buffer(27427) := X"AE00001C";
        ram_buffer(27428) := X"AE000024";
        ram_buffer(27429) := X"8E10002C";
        ram_buffer(27430) := X"00000000";
        ram_buffer(27431) := X"1600FFE3";
        ram_buffer(27432) := X"00000000";
        ram_buffer(27433) := X"8E700044";
        ram_buffer(27434) := X"00000000";
        ram_buffer(27435) := X"16000007";
        ram_buffer(27436) := X"00000000";
        ram_buffer(27437) := X"10000023";
        ram_buffer(27438) := X"00000000";
        ram_buffer(27439) := X"8E10002C";
        ram_buffer(27440) := X"00000000";
        ram_buffer(27441) := X"1200001F";
        ram_buffer(27442) := X"00000000";
        ram_buffer(27443) := X"8E030000";
        ram_buffer(27444) := X"00000000";
        ram_buffer(27445) := X"1460FFF9";
        ram_buffer(27446) := X"00000000";
        ram_buffer(27447) := X"8E070004";
        ram_buffer(27448) := X"8E03000C";
        ram_buffer(27449) := X"24E2FFFF";
        ram_buffer(27450) := X"14600002";
        ram_buffer(27451) := X"0043001B";
        ram_buffer(27452) := X"0007000D";
        ram_buffer(27453) := X"00001012";
        ram_buffer(27454) := X"24420001";
        ram_buffer(27455) := X"0222102A";
        ram_buffer(27456) := X"14400028";
        ram_buffer(27457) := X"02230018";
        ram_buffer(27458) := X"AE070010";
        ram_buffer(27459) := X"8E060008";
        ram_buffer(27460) := X"24050001";
        ram_buffer(27461) := X"0C026A27";
        ram_buffer(27462) := X"02402021";
        ram_buffer(27463) := X"8E63004C";
        ram_buffer(27464) := X"AE020000";
        ram_buffer(27465) := X"AE030014";
        ram_buffer(27466) := X"AE000018";
        ram_buffer(27467) := X"AE00001C";
        ram_buffer(27468) := X"AE000024";
        ram_buffer(27469) := X"8E10002C";
        ram_buffer(27470) := X"00000000";
        ram_buffer(27471) := X"1600FFE3";
        ram_buffer(27472) := X"00000000";
        ram_buffer(27473) := X"8FBF0024";
        ram_buffer(27474) := X"8FB30020";
        ram_buffer(27475) := X"8FB2001C";
        ram_buffer(27476) := X"8FB10018";
        ram_buffer(27477) := X"8FB00014";
        ram_buffer(27478) := X"03E00008";
        ram_buffer(27479) := X"27BD0028";
        ram_buffer(27480) := X"3C113B9A";
        ram_buffer(27481) := X"1000FFA7";
        ram_buffer(27482) := X"3631CA00";
        ram_buffer(27483) := X"8E060008";
        ram_buffer(27484) := X"26050030";
        ram_buffer(27485) := X"02402021";
        ram_buffer(27486) := X"00001812";
        ram_buffer(27487) := X"00000000";
        ram_buffer(27488) := X"00000000";
        ram_buffer(27489) := X"00E60018";
        ram_buffer(27490) := X"00003012";
        ram_buffer(27491) := X"0C026D2D";
        ram_buffer(27492) := X"AE030010";
        ram_buffer(27493) := X"24020001";
        ram_buffer(27494) := X"8E070010";
        ram_buffer(27495) := X"1000FFB3";
        ram_buffer(27496) := X"AE020028";
        ram_buffer(27497) := X"8E060008";
        ram_buffer(27498) := X"26050030";
        ram_buffer(27499) := X"02402021";
        ram_buffer(27500) := X"00001812";
        ram_buffer(27501) := X"AE030010";
        ram_buffer(27502) := X"00000000";
        ram_buffer(27503) := X"00E60018";
        ram_buffer(27504) := X"00003012";
        ram_buffer(27505) := X"0C026D2D";
        ram_buffer(27506) := X"000631C0";
        ram_buffer(27507) := X"24020001";
        ram_buffer(27508) := X"8E070010";
        ram_buffer(27509) := X"1000FFCD";
        ram_buffer(27510) := X"AE020028";
        ram_buffer(27511) := X"8E620044";
        ram_buffer(27512) := X"00000000";
        ram_buffer(27513) := X"1040FFD7";
        ram_buffer(27514) := X"00008021";
        ram_buffer(27515) := X"1000FF65";
        ram_buffer(27516) := X"00008821";
        ram_buffer(27517) := X"1000FF83";
        ram_buffer(27518) := X"24110001";
        ram_buffer(27519) := X"27BDFFC8";
        ram_buffer(27520) := X"24020001";
        ram_buffer(27521) := X"AFB60028";
        ram_buffer(27522) := X"AFB3001C";
        ram_buffer(27523) := X"AFB20018";
        ram_buffer(27524) := X"AFB10014";
        ram_buffer(27525) := X"AFB00010";
        ram_buffer(27526) := X"AFBF0034";
        ram_buffer(27527) := X"AFBE0030";
        ram_buffer(27528) := X"AFB7002C";
        ram_buffer(27529) := X"AFB50024";
        ram_buffer(27530) := X"AFB40020";
        ram_buffer(27531) := X"0080B021";
        ram_buffer(27532) := X"00A08021";
        ram_buffer(27533) := X"00C09021";
        ram_buffer(27534) := X"8C910004";
        ram_buffer(27535) := X"10A2007A";
        ram_buffer(27536) := X"00E09821";
        ram_buffer(27537) := X"8C820000";
        ram_buffer(27538) := X"2415000C";
        ram_buffer(27539) := X"AC450018";
        ram_buffer(27540) := X"8C830000";
        ram_buffer(27541) := X"AC550014";
        ram_buffer(27542) := X"8C620000";
        ram_buffer(27543) := X"00000000";
        ram_buffer(27544) := X"0040F809";
        ram_buffer(27545) := X"00000000";
        ram_buffer(27546) := X"2E020002";
        ram_buffer(27547) := X"8ED40004";
        ram_buffer(27548) := X"1440000A";
        ram_buffer(27549) := X"00000000";
        ram_buffer(27550) := X"8EC20000";
        ram_buffer(27551) := X"00000000";
        ram_buffer(27552) := X"AC500018";
        ram_buffer(27553) := X"8EC30000";
        ram_buffer(27554) := X"AC550014";
        ram_buffer(27555) := X"8C620000";
        ram_buffer(27556) := X"00000000";
        ram_buffer(27557) := X"0040F809";
        ram_buffer(27558) := X"02C02021";
        ram_buffer(27559) := X"00108080";
        ram_buffer(27560) := X"0290A821";
        ram_buffer(27561) := X"8EBE0030";
        ram_buffer(27562) := X"00000000";
        ram_buffer(27563) := X"13C0006B";
        ram_buffer(27564) := X"27828088";
        ram_buffer(27565) := X"8FC30008";
        ram_buffer(27566) := X"00000000";
        ram_buffer(27567) := X"2C620080";
        ram_buffer(27568) := X"14400008";
        ram_buffer(27569) := X"03C01021";
        ram_buffer(27570) := X"1000005F";
        ram_buffer(27571) := X"00000000";
        ram_buffer(27572) := X"8C430008";
        ram_buffer(27573) := X"00000000";
        ram_buffer(27574) := X"2C640080";
        ram_buffer(27575) := X"10800033";
        ram_buffer(27576) := X"0040F021";
        ram_buffer(27577) := X"8FC20000";
        ram_buffer(27578) := X"00000000";
        ram_buffer(27579) := X"1440FFF8";
        ram_buffer(27580) := X"00000000";
        ram_buffer(27581) := X"27828080";
        ram_buffer(27582) := X"00508021";
        ram_buffer(27583) := X"8E030000";
        ram_buffer(27584) := X"3C023B9A";
        ram_buffer(27585) := X"3442C971";
        ram_buffer(27586) := X"00608021";
        ram_buffer(27587) := X"0062182B";
        ram_buffer(27588) := X"10600047";
        ram_buffer(27589) := X"00000000";
        ram_buffer(27590) := X"26170090";
        ram_buffer(27591) := X"02C02021";
        ram_buffer(27592) := X"0C026D23";
        ram_buffer(27593) := X"02E02821";
        ram_buffer(27594) := X"14400014";
        ram_buffer(27595) := X"00000000";
        ram_buffer(27596) := X"00108042";
        ram_buffer(27597) := X"2E020032";
        ram_buffer(27598) := X"1040FFF7";
        ram_buffer(27599) := X"24030002";
        ram_buffer(27600) := X"8EC20000";
        ram_buffer(27601) := X"00000000";
        ram_buffer(27602) := X"AC430018";
        ram_buffer(27603) := X"8EC30000";
        ram_buffer(27604) := X"24050035";
        ram_buffer(27605) := X"AC450014";
        ram_buffer(27606) := X"8C620000";
        ram_buffer(27607) := X"02C02021";
        ram_buffer(27608) := X"0040F809";
        ram_buffer(27609) := X"26170090";
        ram_buffer(27610) := X"02C02021";
        ram_buffer(27611) := X"0C026D23";
        ram_buffer(27612) := X"02E02821";
        ram_buffer(27613) := X"1040FFEE";
        ram_buffer(27614) := X"00000000";
        ram_buffer(27615) := X"8E840048";
        ram_buffer(27616) := X"26030080";
        ram_buffer(27617) := X"00973021";
        ram_buffer(27618) := X"AE860048";
        ram_buffer(27619) := X"AC400000";
        ram_buffer(27620) := X"AC400004";
        ram_buffer(27621) := X"13C00028";
        ram_buffer(27622) := X"AC430008";
        ram_buffer(27623) := X"AFC20000";
        ram_buffer(27624) := X"24040080";
        ram_buffer(27625) := X"10000005";
        ram_buffer(27626) := X"24050010";
        ram_buffer(27627) := X"8C440004";
        ram_buffer(27628) := X"00000000";
        ram_buffer(27629) := X"24850010";
        ram_buffer(27630) := X"24840080";
        ram_buffer(27631) := X"AC440004";
        ram_buffer(27632) := X"2463FF80";
        ram_buffer(27633) := X"8FA40048";
        ram_buffer(27634) := X"AC430008";
        ram_buffer(27635) := X"00451021";
        ram_buffer(27636) := X"8E230040";
        ram_buffer(27637) := X"8FBF0034";
        ram_buffer(27638) := X"AC440004";
        ram_buffer(27639) := X"8FA4004C";
        ram_buffer(27640) := X"AC530008";
        ram_buffer(27641) := X"AC520020";
        ram_buffer(27642) := X"AC400000";
        ram_buffer(27643) := X"AC44000C";
        ram_buffer(27644) := X"AC400028";
        ram_buffer(27645) := X"AC43002C";
        ram_buffer(27646) := X"8FBE0030";
        ram_buffer(27647) := X"AE220040";
        ram_buffer(27648) := X"8FB7002C";
        ram_buffer(27649) := X"8FB60028";
        ram_buffer(27650) := X"8FB50024";
        ram_buffer(27651) := X"8FB40020";
        ram_buffer(27652) := X"8FB3001C";
        ram_buffer(27653) := X"8FB20018";
        ram_buffer(27654) := X"8FB10014";
        ram_buffer(27655) := X"8FB00010";
        ram_buffer(27656) := X"03E00008";
        ram_buffer(27657) := X"27BD0038";
        ram_buffer(27658) := X"1000FF9C";
        ram_buffer(27659) := X"0220A021";
        ram_buffer(27660) := X"1000FFB9";
        ram_buffer(27661) := X"2450FFFF";
        ram_buffer(27662) := X"AEA20030";
        ram_buffer(27663) := X"24040080";
        ram_buffer(27664) := X"1000FFDE";
        ram_buffer(27665) := X"24050010";
        ram_buffer(27666) := X"8FC40004";
        ram_buffer(27667) := X"00000000";
        ram_buffer(27668) := X"24850010";
        ram_buffer(27669) := X"1000FFD9";
        ram_buffer(27670) := X"24840080";
        ram_buffer(27671) := X"00508021";
        ram_buffer(27672) := X"8E030000";
        ram_buffer(27673) := X"1000FFA7";
        ram_buffer(27674) := X"3C023B9A";
        ram_buffer(27675) := X"27BDFFC8";
        ram_buffer(27676) := X"24020001";
        ram_buffer(27677) := X"AFB60028";
        ram_buffer(27678) := X"AFB3001C";
        ram_buffer(27679) := X"AFB20018";
        ram_buffer(27680) := X"AFB10014";
        ram_buffer(27681) := X"AFB00010";
        ram_buffer(27682) := X"AFBF0034";
        ram_buffer(27683) := X"AFBE0030";
        ram_buffer(27684) := X"AFB7002C";
        ram_buffer(27685) := X"AFB50024";
        ram_buffer(27686) := X"AFB40020";
        ram_buffer(27687) := X"0080B021";
        ram_buffer(27688) := X"00A08021";
        ram_buffer(27689) := X"00C09021";
        ram_buffer(27690) := X"8C910004";
        ram_buffer(27691) := X"10A2007A";
        ram_buffer(27692) := X"00E09821";
        ram_buffer(27693) := X"8C820000";
        ram_buffer(27694) := X"2415000C";
        ram_buffer(27695) := X"AC450018";
        ram_buffer(27696) := X"8C830000";
        ram_buffer(27697) := X"AC550014";
        ram_buffer(27698) := X"8C620000";
        ram_buffer(27699) := X"00000000";
        ram_buffer(27700) := X"0040F809";
        ram_buffer(27701) := X"00000000";
        ram_buffer(27702) := X"2E020002";
        ram_buffer(27703) := X"8ED40004";
        ram_buffer(27704) := X"1440000A";
        ram_buffer(27705) := X"00000000";
        ram_buffer(27706) := X"8EC20000";
        ram_buffer(27707) := X"00000000";
        ram_buffer(27708) := X"AC500018";
        ram_buffer(27709) := X"8EC30000";
        ram_buffer(27710) := X"AC550014";
        ram_buffer(27711) := X"8C620000";
        ram_buffer(27712) := X"00000000";
        ram_buffer(27713) := X"0040F809";
        ram_buffer(27714) := X"02C02021";
        ram_buffer(27715) := X"00108080";
        ram_buffer(27716) := X"0290A821";
        ram_buffer(27717) := X"8EBE0030";
        ram_buffer(27718) := X"00000000";
        ram_buffer(27719) := X"13C0006B";
        ram_buffer(27720) := X"27828088";
        ram_buffer(27721) := X"8FC30008";
        ram_buffer(27722) := X"00000000";
        ram_buffer(27723) := X"2C620080";
        ram_buffer(27724) := X"14400008";
        ram_buffer(27725) := X"03C01021";
        ram_buffer(27726) := X"1000005F";
        ram_buffer(27727) := X"00000000";
        ram_buffer(27728) := X"8C430008";
        ram_buffer(27729) := X"00000000";
        ram_buffer(27730) := X"2C640080";
        ram_buffer(27731) := X"10800033";
        ram_buffer(27732) := X"0040F021";
        ram_buffer(27733) := X"8FC20000";
        ram_buffer(27734) := X"00000000";
        ram_buffer(27735) := X"1440FFF8";
        ram_buffer(27736) := X"00000000";
        ram_buffer(27737) := X"27828080";
        ram_buffer(27738) := X"00508021";
        ram_buffer(27739) := X"8E030000";
        ram_buffer(27740) := X"3C023B9A";
        ram_buffer(27741) := X"3442C971";
        ram_buffer(27742) := X"00608021";
        ram_buffer(27743) := X"0062182B";
        ram_buffer(27744) := X"10600047";
        ram_buffer(27745) := X"00000000";
        ram_buffer(27746) := X"26170090";
        ram_buffer(27747) := X"02C02021";
        ram_buffer(27748) := X"0C026D23";
        ram_buffer(27749) := X"02E02821";
        ram_buffer(27750) := X"14400014";
        ram_buffer(27751) := X"00000000";
        ram_buffer(27752) := X"00108042";
        ram_buffer(27753) := X"2E020032";
        ram_buffer(27754) := X"1040FFF7";
        ram_buffer(27755) := X"24030002";
        ram_buffer(27756) := X"8EC20000";
        ram_buffer(27757) := X"00000000";
        ram_buffer(27758) := X"AC430018";
        ram_buffer(27759) := X"8EC30000";
        ram_buffer(27760) := X"24050035";
        ram_buffer(27761) := X"AC450014";
        ram_buffer(27762) := X"8C620000";
        ram_buffer(27763) := X"02C02021";
        ram_buffer(27764) := X"0040F809";
        ram_buffer(27765) := X"26170090";
        ram_buffer(27766) := X"02C02021";
        ram_buffer(27767) := X"0C026D23";
        ram_buffer(27768) := X"02E02821";
        ram_buffer(27769) := X"1040FFEE";
        ram_buffer(27770) := X"00000000";
        ram_buffer(27771) := X"8E840048";
        ram_buffer(27772) := X"26030080";
        ram_buffer(27773) := X"00973021";
        ram_buffer(27774) := X"AE860048";
        ram_buffer(27775) := X"AC400000";
        ram_buffer(27776) := X"AC400004";
        ram_buffer(27777) := X"13C00028";
        ram_buffer(27778) := X"AC430008";
        ram_buffer(27779) := X"AFC20000";
        ram_buffer(27780) := X"24040080";
        ram_buffer(27781) := X"10000005";
        ram_buffer(27782) := X"24050010";
        ram_buffer(27783) := X"8C440004";
        ram_buffer(27784) := X"00000000";
        ram_buffer(27785) := X"24850010";
        ram_buffer(27786) := X"24840080";
        ram_buffer(27787) := X"AC440004";
        ram_buffer(27788) := X"2463FF80";
        ram_buffer(27789) := X"8FA40048";
        ram_buffer(27790) := X"AC430008";
        ram_buffer(27791) := X"00451021";
        ram_buffer(27792) := X"8E230044";
        ram_buffer(27793) := X"8FBF0034";
        ram_buffer(27794) := X"AC440004";
        ram_buffer(27795) := X"8FA4004C";
        ram_buffer(27796) := X"AC530008";
        ram_buffer(27797) := X"AC520020";
        ram_buffer(27798) := X"AC400000";
        ram_buffer(27799) := X"AC44000C";
        ram_buffer(27800) := X"AC400028";
        ram_buffer(27801) := X"AC43002C";
        ram_buffer(27802) := X"8FBE0030";
        ram_buffer(27803) := X"AE220044";
        ram_buffer(27804) := X"8FB7002C";
        ram_buffer(27805) := X"8FB60028";
        ram_buffer(27806) := X"8FB50024";
        ram_buffer(27807) := X"8FB40020";
        ram_buffer(27808) := X"8FB3001C";
        ram_buffer(27809) := X"8FB20018";
        ram_buffer(27810) := X"8FB10014";
        ram_buffer(27811) := X"8FB00010";
        ram_buffer(27812) := X"03E00008";
        ram_buffer(27813) := X"27BD0038";
        ram_buffer(27814) := X"1000FF9C";
        ram_buffer(27815) := X"0220A021";
        ram_buffer(27816) := X"1000FFB9";
        ram_buffer(27817) := X"2450FFFF";
        ram_buffer(27818) := X"AEA20030";
        ram_buffer(27819) := X"24040080";
        ram_buffer(27820) := X"1000FFDE";
        ram_buffer(27821) := X"24050010";
        ram_buffer(27822) := X"8FC40004";
        ram_buffer(27823) := X"00000000";
        ram_buffer(27824) := X"24850010";
        ram_buffer(27825) := X"1000FFD9";
        ram_buffer(27826) := X"24840080";
        ram_buffer(27827) := X"00508021";
        ram_buffer(27828) := X"8E030000";
        ram_buffer(27829) := X"1000FFA7";
        ram_buffer(27830) := X"3C023B9A";
        ram_buffer(27831) := X"27BDFFD8";
        ram_buffer(27832) := X"AFBF0024";
        ram_buffer(27833) := X"AFB10020";
        ram_buffer(27834) := X"AFB0001C";
        ram_buffer(27835) := X"00808821";
        ram_buffer(27836) := X"0C026D33";
        ram_buffer(27837) := X"AC800004";
        ram_buffer(27838) := X"24050050";
        ram_buffer(27839) := X"02202021";
        ram_buffer(27840) := X"0C026D23";
        ram_buffer(27841) := X"AFA20010";
        ram_buffer(27842) := X"10400053";
        ram_buffer(27843) := X"00408021";
        ram_buffer(27844) := X"3C02100A";
        ram_buffer(27845) := X"2442966C";
        ram_buffer(27846) := X"8FA30010";
        ram_buffer(27847) := X"AE020000";
        ram_buffer(27848) := X"3C02100A";
        ram_buffer(27849) := X"24429AD8";
        ram_buffer(27850) := X"AE020004";
        ram_buffer(27851) := X"3C02100A";
        ram_buffer(27852) := X"2442A64C";
        ram_buffer(27853) := X"AE020008";
        ram_buffer(27854) := X"3C02100A";
        ram_buffer(27855) := X"2442A89C";
        ram_buffer(27856) := X"AE02000C";
        ram_buffer(27857) := X"3C02100A";
        ram_buffer(27858) := X"2442ADFC";
        ram_buffer(27859) := X"AE020010";
        ram_buffer(27860) := X"3C02100A";
        ram_buffer(27861) := X"2442B06C";
        ram_buffer(27862) := X"AE020014";
        ram_buffer(27863) := X"3C02100A";
        ram_buffer(27864) := X"2442AADC";
        ram_buffer(27865) := X"AE020018";
        ram_buffer(27866) := X"3C02100A";
        ram_buffer(27867) := X"2442A140";
        ram_buffer(27868) := X"AE02001C";
        ram_buffer(27869) := X"3C02100A";
        ram_buffer(27870) := X"24429C14";
        ram_buffer(27871) := X"AE020020";
        ram_buffer(27872) := X"3C02100A";
        ram_buffer(27873) := X"244298B8";
        ram_buffer(27874) := X"AE020024";
        ram_buffer(27875) := X"3C02100A";
        ram_buffer(27876) := X"24429A8C";
        ram_buffer(27877) := X"AE020028";
        ram_buffer(27878) := X"3C04100D";
        ram_buffer(27879) := X"24020050";
        ram_buffer(27880) := X"AE03002C";
        ram_buffer(27881) := X"AE000034";
        ram_buffer(27882) := X"AE00003C";
        ram_buffer(27883) := X"AE000030";
        ram_buffer(27884) := X"AE000038";
        ram_buffer(27885) := X"AE000040";
        ram_buffer(27886) := X"AE000044";
        ram_buffer(27887) := X"AE020048";
        ram_buffer(27888) := X"24849DE4";
        ram_buffer(27889) := X"0C027901";
        ram_buffer(27890) := X"AE300004";
        ram_buffer(27891) := X"10400018";
        ram_buffer(27892) := X"3C05100C";
        ram_buffer(27893) := X"00402021";
        ram_buffer(27894) := X"27A70014";
        ram_buffer(27895) := X"24020078";
        ram_buffer(27896) := X"27A60010";
        ram_buffer(27897) := X"24A57B58";
        ram_buffer(27898) := X"0C028409";
        ram_buffer(27899) := X"A3A20014";
        ram_buffer(27900) := X"1840000F";
        ram_buffer(27901) := X"2403004D";
        ram_buffer(27902) := X"93A20014";
        ram_buffer(27903) := X"00000000";
        ram_buffer(27904) := X"304200DF";
        ram_buffer(27905) := X"00021600";
        ram_buffer(27906) := X"00021603";
        ram_buffer(27907) := X"8FA40010";
        ram_buffer(27908) := X"1043000C";
        ram_buffer(27909) := X"00041080";
        ram_buffer(27910) := X"00041080";
        ram_buffer(27911) := X"000419C0";
        ram_buffer(27912) := X"00621023";
        ram_buffer(27913) := X"00441021";
        ram_buffer(27914) := X"000210C0";
        ram_buffer(27915) := X"AE02002C";
        ram_buffer(27916) := X"8FBF0024";
        ram_buffer(27917) := X"8FB10020";
        ram_buffer(27918) := X"8FB0001C";
        ram_buffer(27919) := X"03E00008";
        ram_buffer(27920) := X"27BD0028";
        ram_buffer(27921) := X"000419C0";
        ram_buffer(27922) := X"00621023";
        ram_buffer(27923) := X"00441021";
        ram_buffer(27924) := X"1000FFF1";
        ram_buffer(27925) := X"000220C0";
        ram_buffer(27926) := X"0C026D35";
        ram_buffer(27927) := X"02202021";
        ram_buffer(27928) := X"8E220000";
        ram_buffer(27929) := X"24040035";
        ram_buffer(27930) := X"AC400018";
        ram_buffer(27931) := X"8E230000";
        ram_buffer(27932) := X"AC440014";
        ram_buffer(27933) := X"8C620000";
        ram_buffer(27934) := X"00000000";
        ram_buffer(27935) := X"0040F809";
        ram_buffer(27936) := X"02202021";
        ram_buffer(27937) := X"1000FFA3";
        ram_buffer(27938) := X"3C02100A";
        ram_buffer(27939) := X"08027A3D";
        ram_buffer(27940) := X"00A02021";
        ram_buffer(27941) := X"08027A4D";
        ram_buffer(27942) := X"00A02021";
        ram_buffer(27943) := X"08027A3D";
        ram_buffer(27944) := X"00A02021";
        ram_buffer(27945) := X"08027A4D";
        ram_buffer(27946) := X"00A02021";
        ram_buffer(27947) := X"03E00008";
        ram_buffer(27948) := X"00C01021";
        ram_buffer(27949) := X"8C820000";
        ram_buffer(27950) := X"24030030";
        ram_buffer(27951) := X"8C590000";
        ram_buffer(27952) := X"00000000";
        ram_buffer(27953) := X"03200008";
        ram_buffer(27954) := X"AC430014";
        ram_buffer(27955) := X"03E00008";
        ram_buffer(27956) := X"00001021";
        ram_buffer(27957) := X"03E00008";
        ram_buffer(27958) := X"00000000";
        ram_buffer(27959) := X"27BDFFE8";
        ram_buffer(27960) := X"AFBF0014";
        ram_buffer(27961) := X"AFBE0010";
        ram_buffer(27962) := X"03A0F021";
        ram_buffer(27963) := X"AFC40018";
        ram_buffer(27964) := X"00002821";
        ram_buffer(27965) := X"8FC40018";
        ram_buffer(27966) := X"0C02AD8C";
        ram_buffer(27967) := X"00000000";
        ram_buffer(27968) := X"8F82809C";
        ram_buffer(27969) := X"00000000";
        ram_buffer(27970) := X"8C42003C";
        ram_buffer(27971) := X"00000000";
        ram_buffer(27972) := X"10400009";
        ram_buffer(27973) := X"00000000";
        ram_buffer(27974) := X"8F82809C";
        ram_buffer(27975) := X"00000000";
        ram_buffer(27976) := X"8C42003C";
        ram_buffer(27977) := X"8F83809C";
        ram_buffer(27978) := X"00000000";
        ram_buffer(27979) := X"00602021";
        ram_buffer(27980) := X"0040F809";
        ram_buffer(27981) := X"00000000";
        ram_buffer(27982) := X"8FC40018";
        ram_buffer(27983) := X"0C02FB62";
        ram_buffer(27984) := X"00000000";
        ram_buffer(27985) := X"27BDFFD8";
        ram_buffer(27986) := X"AFBF0024";
        ram_buffer(27987) := X"AFBE0020";
        ram_buffer(27988) := X"AFB0001C";
        ram_buffer(27989) := X"03A0F021";
        ram_buffer(27990) := X"AFC40028";
        ram_buffer(27991) := X"00A08021";
        ram_buffer(27992) := X"16000004";
        ram_buffer(27993) := X"00000000";
        ram_buffer(27994) := X"00001021";
        ram_buffer(27995) := X"10000058";
        ram_buffer(27996) := X"00000000";
        ram_buffer(27997) := X"8FC20028";
        ram_buffer(27998) := X"00000000";
        ram_buffer(27999) := X"AFC20014";
        ram_buffer(28000) := X"8FC20014";
        ram_buffer(28001) := X"00000000";
        ram_buffer(28002) := X"1040000A";
        ram_buffer(28003) := X"00000000";
        ram_buffer(28004) := X"8FC20014";
        ram_buffer(28005) := X"00000000";
        ram_buffer(28006) := X"8C420038";
        ram_buffer(28007) := X"00000000";
        ram_buffer(28008) := X"14400004";
        ram_buffer(28009) := X"00000000";
        ram_buffer(28010) := X"8FC40014";
        ram_buffer(28011) := X"0C027069";
        ram_buffer(28012) := X"00000000";
        ram_buffer(28013) := X"8602000C";
        ram_buffer(28014) := X"00000000";
        ram_buffer(28015) := X"14400004";
        ram_buffer(28016) := X"00000000";
        ram_buffer(28017) := X"00001021";
        ram_buffer(28018) := X"10000041";
        ram_buffer(28019) := X"00000000";
        ram_buffer(28020) := X"02002821";
        ram_buffer(28021) := X"8FC40028";
        ram_buffer(28022) := X"0C026DCB";
        ram_buffer(28023) := X"00000000";
        ram_buffer(28024) := X"AFC20010";
        ram_buffer(28025) := X"8E02002C";
        ram_buffer(28026) := X"00000000";
        ram_buffer(28027) := X"1040000C";
        ram_buffer(28028) := X"00000000";
        ram_buffer(28029) := X"8E02002C";
        ram_buffer(28030) := X"8E03001C";
        ram_buffer(28031) := X"00000000";
        ram_buffer(28032) := X"00602821";
        ram_buffer(28033) := X"8FC40028";
        ram_buffer(28034) := X"0040F809";
        ram_buffer(28035) := X"00000000";
        ram_buffer(28036) := X"04410003";
        ram_buffer(28037) := X"00000000";
        ram_buffer(28038) := X"2402FFFF";
        ram_buffer(28039) := X"AFC20010";
        ram_buffer(28040) := X"8602000C";
        ram_buffer(28041) := X"00000000";
        ram_buffer(28042) := X"3042FFFF";
        ram_buffer(28043) := X"30420080";
        ram_buffer(28044) := X"10400007";
        ram_buffer(28045) := X"00000000";
        ram_buffer(28046) := X"8E020010";
        ram_buffer(28047) := X"00000000";
        ram_buffer(28048) := X"00402821";
        ram_buffer(28049) := X"8FC40028";
        ram_buffer(28050) := X"0C027301";
        ram_buffer(28051) := X"00000000";
        ram_buffer(28052) := X"8E020030";
        ram_buffer(28053) := X"00000000";
        ram_buffer(28054) := X"1040000C";
        ram_buffer(28055) := X"00000000";
        ram_buffer(28056) := X"8E030030";
        ram_buffer(28057) := X"26020040";
        ram_buffer(28058) := X"10620007";
        ram_buffer(28059) := X"00000000";
        ram_buffer(28060) := X"8E020030";
        ram_buffer(28061) := X"00000000";
        ram_buffer(28062) := X"00402821";
        ram_buffer(28063) := X"8FC40028";
        ram_buffer(28064) := X"0C027301";
        ram_buffer(28065) := X"00000000";
        ram_buffer(28066) := X"AE000030";
        ram_buffer(28067) := X"8E020044";
        ram_buffer(28068) := X"00000000";
        ram_buffer(28069) := X"10400008";
        ram_buffer(28070) := X"00000000";
        ram_buffer(28071) := X"8E020044";
        ram_buffer(28072) := X"00000000";
        ram_buffer(28073) := X"00402821";
        ram_buffer(28074) := X"8FC40028";
        ram_buffer(28075) := X"0C027301";
        ram_buffer(28076) := X"00000000";
        ram_buffer(28077) := X"AE000044";
        ram_buffer(28078) := X"0C0270B0";
        ram_buffer(28079) := X"00000000";
        ram_buffer(28080) := X"A600000C";
        ram_buffer(28081) := X"0C0270B9";
        ram_buffer(28082) := X"00000000";
        ram_buffer(28083) := X"8FC20010";
        ram_buffer(28084) := X"03C0E821";
        ram_buffer(28085) := X"8FBF0024";
        ram_buffer(28086) := X"8FBE0020";
        ram_buffer(28087) := X"8FB0001C";
        ram_buffer(28088) := X"27BD0028";
        ram_buffer(28089) := X"03E00008";
        ram_buffer(28090) := X"00000000";
        ram_buffer(28091) := X"27BDFFE8";
        ram_buffer(28092) := X"AFBF0014";
        ram_buffer(28093) := X"AFBE0010";
        ram_buffer(28094) := X"03A0F021";
        ram_buffer(28095) := X"00801821";
        ram_buffer(28096) := X"8F828098";
        ram_buffer(28097) := X"00602821";
        ram_buffer(28098) := X"00402021";
        ram_buffer(28099) := X"0C026D51";
        ram_buffer(28100) := X"00000000";
        ram_buffer(28101) := X"03C0E821";
        ram_buffer(28102) := X"8FBF0014";
        ram_buffer(28103) := X"8FBE0010";
        ram_buffer(28104) := X"27BD0018";
        ram_buffer(28105) := X"03E00008";
        ram_buffer(28106) := X"00000000";
        ram_buffer(28107) := X"27BDFFC8";
        ram_buffer(28108) := X"AFBF0034";
        ram_buffer(28109) := X"AFBE0030";
        ram_buffer(28110) := X"AFB3002C";
        ram_buffer(28111) := X"AFB20028";
        ram_buffer(28112) := X"AFB10024";
        ram_buffer(28113) := X"AFB00020";
        ram_buffer(28114) := X"03A0F021";
        ram_buffer(28115) := X"AFC40038";
        ram_buffer(28116) := X"00A08021";
        ram_buffer(28117) := X"9602000C";
        ram_buffer(28118) := X"00000000";
        ram_buffer(28119) := X"A7C20018";
        ram_buffer(28120) := X"97C20018";
        ram_buffer(28121) := X"00000000";
        ram_buffer(28122) := X"30420008";
        ram_buffer(28123) := X"144000C8";
        ram_buffer(28124) := X"00000000";
        ram_buffer(28125) := X"8602000C";
        ram_buffer(28126) := X"00000000";
        ram_buffer(28127) := X"34420800";
        ram_buffer(28128) := X"00021400";
        ram_buffer(28129) := X"00021403";
        ram_buffer(28130) := X"A602000C";
        ram_buffer(28131) := X"8E020004";
        ram_buffer(28132) := X"00000000";
        ram_buffer(28133) := X"1C400005";
        ram_buffer(28134) := X"00000000";
        ram_buffer(28135) := X"8E02003C";
        ram_buffer(28136) := X"00000000";
        ram_buffer(28137) := X"184000B7";
        ram_buffer(28138) := X"00000000";
        ram_buffer(28139) := X"8E020028";
        ram_buffer(28140) := X"00000000";
        ram_buffer(28141) := X"104000B3";
        ram_buffer(28142) := X"00000000";
        ram_buffer(28143) := X"8FC20038";
        ram_buffer(28144) := X"00000000";
        ram_buffer(28145) := X"8C420000";
        ram_buffer(28146) := X"00000000";
        ram_buffer(28147) := X"AFC2001C";
        ram_buffer(28148) := X"8FC20038";
        ram_buffer(28149) := X"00000000";
        ram_buffer(28150) := X"AC400000";
        ram_buffer(28151) := X"8602000C";
        ram_buffer(28152) := X"00000000";
        ram_buffer(28153) := X"3042FFFF";
        ram_buffer(28154) := X"30421000";
        ram_buffer(28155) := X"10400006";
        ram_buffer(28156) := X"00000000";
        ram_buffer(28157) := X"8E020050";
        ram_buffer(28158) := X"00000000";
        ram_buffer(28159) := X"AFC20010";
        ram_buffer(28160) := X"10000032";
        ram_buffer(28161) := X"00000000";
        ram_buffer(28162) := X"8E020028";
        ram_buffer(28163) := X"8E03001C";
        ram_buffer(28164) := X"24070001";
        ram_buffer(28165) := X"00003021";
        ram_buffer(28166) := X"00602821";
        ram_buffer(28167) := X"8FC40038";
        ram_buffer(28168) := X"0040F809";
        ram_buffer(28169) := X"00000000";
        ram_buffer(28170) := X"AFC20010";
        ram_buffer(28171) := X"8FC30010";
        ram_buffer(28172) := X"2402FFFF";
        ram_buffer(28173) := X"14620025";
        ram_buffer(28174) := X"00000000";
        ram_buffer(28175) := X"8FC20038";
        ram_buffer(28176) := X"00000000";
        ram_buffer(28177) := X"8C420000";
        ram_buffer(28178) := X"00000000";
        ram_buffer(28179) := X"1040001F";
        ram_buffer(28180) := X"00000000";
        ram_buffer(28181) := X"2402FFFF";
        ram_buffer(28182) := X"AFC20014";
        ram_buffer(28183) := X"8FC20038";
        ram_buffer(28184) := X"00000000";
        ram_buffer(28185) := X"8C430000";
        ram_buffer(28186) := X"2402001D";
        ram_buffer(28187) := X"10620007";
        ram_buffer(28188) := X"00000000";
        ram_buffer(28189) := X"8FC20038";
        ram_buffer(28190) := X"00000000";
        ram_buffer(28191) := X"8C430000";
        ram_buffer(28192) := X"24020016";
        ram_buffer(28193) := X"14620008";
        ram_buffer(28194) := X"00000000";
        ram_buffer(28195) := X"AFC00014";
        ram_buffer(28196) := X"8FC20038";
        ram_buffer(28197) := X"8FC3001C";
        ram_buffer(28198) := X"00000000";
        ram_buffer(28199) := X"AC430000";
        ram_buffer(28200) := X"10000007";
        ram_buffer(28201) := X"00000000";
        ram_buffer(28202) := X"8602000C";
        ram_buffer(28203) := X"00000000";
        ram_buffer(28204) := X"34420040";
        ram_buffer(28205) := X"00021400";
        ram_buffer(28206) := X"00021403";
        ram_buffer(28207) := X"A602000C";
        ram_buffer(28208) := X"8FC20014";
        ram_buffer(28209) := X"100000A5";
        ram_buffer(28210) := X"00000000";
        ram_buffer(28211) := X"8602000C";
        ram_buffer(28212) := X"00000000";
        ram_buffer(28213) := X"3042FFFF";
        ram_buffer(28214) := X"30420004";
        ram_buffer(28215) := X"1040000F";
        ram_buffer(28216) := X"00000000";
        ram_buffer(28217) := X"8E020004";
        ram_buffer(28218) := X"8FC30010";
        ram_buffer(28219) := X"00000000";
        ram_buffer(28220) := X"00621023";
        ram_buffer(28221) := X"AFC20010";
        ram_buffer(28222) := X"8E020030";
        ram_buffer(28223) := X"00000000";
        ram_buffer(28224) := X"10400006";
        ram_buffer(28225) := X"00000000";
        ram_buffer(28226) := X"8E02003C";
        ram_buffer(28227) := X"8FC30010";
        ram_buffer(28228) := X"00000000";
        ram_buffer(28229) := X"00621023";
        ram_buffer(28230) := X"AFC20010";
        ram_buffer(28231) := X"8E020028";
        ram_buffer(28232) := X"8E03001C";
        ram_buffer(28233) := X"00003821";
        ram_buffer(28234) := X"8FC60010";
        ram_buffer(28235) := X"00602821";
        ram_buffer(28236) := X"8FC40038";
        ram_buffer(28237) := X"0040F809";
        ram_buffer(28238) := X"00000000";
        ram_buffer(28239) := X"AFC20010";
        ram_buffer(28240) := X"8FC30010";
        ram_buffer(28241) := X"2402FFFF";
        ram_buffer(28242) := X"14620013";
        ram_buffer(28243) := X"00000000";
        ram_buffer(28244) := X"8FC20038";
        ram_buffer(28245) := X"00000000";
        ram_buffer(28246) := X"8C420000";
        ram_buffer(28247) := X"00000000";
        ram_buffer(28248) := X"1040000D";
        ram_buffer(28249) := X"00000000";
        ram_buffer(28250) := X"8FC20038";
        ram_buffer(28251) := X"00000000";
        ram_buffer(28252) := X"8C430000";
        ram_buffer(28253) := X"2402001D";
        ram_buffer(28254) := X"10620007";
        ram_buffer(28255) := X"00000000";
        ram_buffer(28256) := X"8FC20038";
        ram_buffer(28257) := X"00000000";
        ram_buffer(28258) := X"8C430000";
        ram_buffer(28259) := X"24020016";
        ram_buffer(28260) := X"14620033";
        ram_buffer(28261) := X"00000000";
        ram_buffer(28262) := X"8603000C";
        ram_buffer(28263) := X"2402F7FF";
        ram_buffer(28264) := X"00621024";
        ram_buffer(28265) := X"00021400";
        ram_buffer(28266) := X"00021403";
        ram_buffer(28267) := X"A602000C";
        ram_buffer(28268) := X"AE000004";
        ram_buffer(28269) := X"8E020010";
        ram_buffer(28270) := X"00000000";
        ram_buffer(28271) := X"AE020000";
        ram_buffer(28272) := X"8602000C";
        ram_buffer(28273) := X"00000000";
        ram_buffer(28274) := X"3042FFFF";
        ram_buffer(28275) := X"30421000";
        ram_buffer(28276) := X"1040000E";
        ram_buffer(28277) := X"00000000";
        ram_buffer(28278) := X"8FC30010";
        ram_buffer(28279) := X"2402FFFF";
        ram_buffer(28280) := X"14620007";
        ram_buffer(28281) := X"00000000";
        ram_buffer(28282) := X"8FC20038";
        ram_buffer(28283) := X"00000000";
        ram_buffer(28284) := X"8C420000";
        ram_buffer(28285) := X"00000000";
        ram_buffer(28286) := X"14400004";
        ram_buffer(28287) := X"00000000";
        ram_buffer(28288) := X"8FC20010";
        ram_buffer(28289) := X"00000000";
        ram_buffer(28290) := X"AE020050";
        ram_buffer(28291) := X"8FC20038";
        ram_buffer(28292) := X"8FC3001C";
        ram_buffer(28293) := X"00000000";
        ram_buffer(28294) := X"AC430000";
        ram_buffer(28295) := X"8E020030";
        ram_buffer(28296) := X"00000000";
        ram_buffer(28297) := X"10400017";
        ram_buffer(28298) := X"00000000";
        ram_buffer(28299) := X"8E030030";
        ram_buffer(28300) := X"26020040";
        ram_buffer(28301) := X"10620007";
        ram_buffer(28302) := X"00000000";
        ram_buffer(28303) := X"8E020030";
        ram_buffer(28304) := X"00000000";
        ram_buffer(28305) := X"00402821";
        ram_buffer(28306) := X"8FC40038";
        ram_buffer(28307) := X"0C027301";
        ram_buffer(28308) := X"00000000";
        ram_buffer(28309) := X"AE000030";
        ram_buffer(28310) := X"1000000A";
        ram_buffer(28311) := X"00000000";
        ram_buffer(28312) := X"8602000C";
        ram_buffer(28313) := X"00000000";
        ram_buffer(28314) := X"34420040";
        ram_buffer(28315) := X"00021400";
        ram_buffer(28316) := X"00021403";
        ram_buffer(28317) := X"A602000C";
        ram_buffer(28318) := X"2402FFFF";
        ram_buffer(28319) := X"10000037";
        ram_buffer(28320) := X"00000000";
        ram_buffer(28321) := X"00001021";
        ram_buffer(28322) := X"10000034";
        ram_buffer(28323) := X"00000000";
        ram_buffer(28324) := X"8E110010";
        ram_buffer(28325) := X"00000000";
        ram_buffer(28326) := X"16200004";
        ram_buffer(28327) := X"00000000";
        ram_buffer(28328) := X"00001021";
        ram_buffer(28329) := X"1000002D";
        ram_buffer(28330) := X"00000000";
        ram_buffer(28331) := X"8E020000";
        ram_buffer(28332) := X"00000000";
        ram_buffer(28333) := X"00401821";
        ram_buffer(28334) := X"02201021";
        ram_buffer(28335) := X"00629023";
        ram_buffer(28336) := X"AE110000";
        ram_buffer(28337) := X"97C20018";
        ram_buffer(28338) := X"00000000";
        ram_buffer(28339) := X"30420003";
        ram_buffer(28340) := X"14400004";
        ram_buffer(28341) := X"00000000";
        ram_buffer(28342) := X"8E020014";
        ram_buffer(28343) := X"10000002";
        ram_buffer(28344) := X"00000000";
        ram_buffer(28345) := X"00001021";
        ram_buffer(28346) := X"AE020008";
        ram_buffer(28347) := X"10000018";
        ram_buffer(28348) := X"00000000";
        ram_buffer(28349) := X"8E020024";
        ram_buffer(28350) := X"8E03001C";
        ram_buffer(28351) := X"02403821";
        ram_buffer(28352) := X"02203021";
        ram_buffer(28353) := X"00602821";
        ram_buffer(28354) := X"8FC40038";
        ram_buffer(28355) := X"0040F809";
        ram_buffer(28356) := X"00000000";
        ram_buffer(28357) := X"00409821";
        ram_buffer(28358) := X"1E60000A";
        ram_buffer(28359) := X"00000000";
        ram_buffer(28360) := X"8602000C";
        ram_buffer(28361) := X"00000000";
        ram_buffer(28362) := X"34420040";
        ram_buffer(28363) := X"00021400";
        ram_buffer(28364) := X"00021403";
        ram_buffer(28365) := X"A602000C";
        ram_buffer(28366) := X"2402FFFF";
        ram_buffer(28367) := X"10000007";
        ram_buffer(28368) := X"00000000";
        ram_buffer(28369) := X"02601021";
        ram_buffer(28370) := X"02228821";
        ram_buffer(28371) := X"02539023";
        ram_buffer(28372) := X"1E40FFE8";
        ram_buffer(28373) := X"00000000";
        ram_buffer(28374) := X"00001021";
        ram_buffer(28375) := X"03C0E821";
        ram_buffer(28376) := X"8FBF0034";
        ram_buffer(28377) := X"8FBE0030";
        ram_buffer(28378) := X"8FB3002C";
        ram_buffer(28379) := X"8FB20028";
        ram_buffer(28380) := X"8FB10024";
        ram_buffer(28381) := X"8FB00020";
        ram_buffer(28382) := X"27BD0038";
        ram_buffer(28383) := X"03E00008";
        ram_buffer(28384) := X"00000000";
        ram_buffer(28385) := X"27BDFFD8";
        ram_buffer(28386) := X"AFBF0024";
        ram_buffer(28387) := X"AFBE0020";
        ram_buffer(28388) := X"AFB0001C";
        ram_buffer(28389) := X"03A0F021";
        ram_buffer(28390) := X"AFC40028";
        ram_buffer(28391) := X"00A08021";
        ram_buffer(28392) := X"8FC20028";
        ram_buffer(28393) := X"00000000";
        ram_buffer(28394) := X"AFC20010";
        ram_buffer(28395) := X"8FC20010";
        ram_buffer(28396) := X"00000000";
        ram_buffer(28397) := X"1040000A";
        ram_buffer(28398) := X"00000000";
        ram_buffer(28399) := X"8FC20010";
        ram_buffer(28400) := X"00000000";
        ram_buffer(28401) := X"8C420038";
        ram_buffer(28402) := X"00000000";
        ram_buffer(28403) := X"14400004";
        ram_buffer(28404) := X"00000000";
        ram_buffer(28405) := X"8FC40010";
        ram_buffer(28406) := X"0C027069";
        ram_buffer(28407) := X"00000000";
        ram_buffer(28408) := X"8602000C";
        ram_buffer(28409) := X"00000000";
        ram_buffer(28410) := X"14400004";
        ram_buffer(28411) := X"00000000";
        ram_buffer(28412) := X"00001021";
        ram_buffer(28413) := X"10000007";
        ram_buffer(28414) := X"00000000";
        ram_buffer(28415) := X"02002821";
        ram_buffer(28416) := X"8FC40028";
        ram_buffer(28417) := X"0C026DCB";
        ram_buffer(28418) := X"00000000";
        ram_buffer(28419) := X"AFC20014";
        ram_buffer(28420) := X"8FC20014";
        ram_buffer(28421) := X"03C0E821";
        ram_buffer(28422) := X"8FBF0024";
        ram_buffer(28423) := X"8FBE0020";
        ram_buffer(28424) := X"8FB0001C";
        ram_buffer(28425) := X"27BD0028";
        ram_buffer(28426) := X"03E00008";
        ram_buffer(28427) := X"00000000";
        ram_buffer(28428) := X"27BDFFE8";
        ram_buffer(28429) := X"AFBF0014";
        ram_buffer(28430) := X"AFBE0010";
        ram_buffer(28431) := X"03A0F021";
        ram_buffer(28432) := X"00801021";
        ram_buffer(28433) := X"14400009";
        ram_buffer(28434) := X"00000000";
        ram_buffer(28435) := X"8F83809C";
        ram_buffer(28436) := X"3C02100A";
        ram_buffer(28437) := X"2445BB84";
        ram_buffer(28438) := X"00602021";
        ram_buffer(28439) := X"0C02783C";
        ram_buffer(28440) := X"00000000";
        ram_buffer(28441) := X"10000006";
        ram_buffer(28442) := X"00000000";
        ram_buffer(28443) := X"8F838098";
        ram_buffer(28444) := X"00402821";
        ram_buffer(28445) := X"00602021";
        ram_buffer(28446) := X"0C026EE1";
        ram_buffer(28447) := X"00000000";
        ram_buffer(28448) := X"03C0E821";
        ram_buffer(28449) := X"8FBF0014";
        ram_buffer(28450) := X"8FBE0010";
        ram_buffer(28451) := X"27BD0018";
        ram_buffer(28452) := X"03E00008";
        ram_buffer(28453) := X"00000000";
        ram_buffer(28454) := X"27BDFFE8";
        ram_buffer(28455) := X"AFBF0014";
        ram_buffer(28456) := X"AFBE0010";
        ram_buffer(28457) := X"03A0F021";
        ram_buffer(28458) := X"AFC40018";
        ram_buffer(28459) := X"AFC5001C";
        ram_buffer(28460) := X"AFC60020";
        ram_buffer(28461) := X"AFC70024";
        ram_buffer(28462) := X"8FC20018";
        ram_buffer(28463) := X"00000000";
        ram_buffer(28464) := X"AC400000";
        ram_buffer(28465) := X"8FC20018";
        ram_buffer(28466) := X"00000000";
        ram_buffer(28467) := X"AC400004";
        ram_buffer(28468) := X"8FC20018";
        ram_buffer(28469) := X"00000000";
        ram_buffer(28470) := X"AC400008";
        ram_buffer(28471) := X"8FC2001C";
        ram_buffer(28472) := X"00000000";
        ram_buffer(28473) := X"00021C00";
        ram_buffer(28474) := X"00031C03";
        ram_buffer(28475) := X"8FC20018";
        ram_buffer(28476) := X"00000000";
        ram_buffer(28477) := X"A443000C";
        ram_buffer(28478) := X"8FC20018";
        ram_buffer(28479) := X"00000000";
        ram_buffer(28480) := X"AC400064";
        ram_buffer(28481) := X"8FC20020";
        ram_buffer(28482) := X"00000000";
        ram_buffer(28483) := X"00021C00";
        ram_buffer(28484) := X"00031C03";
        ram_buffer(28485) := X"8FC20018";
        ram_buffer(28486) := X"00000000";
        ram_buffer(28487) := X"A443000E";
        ram_buffer(28488) := X"8FC20018";
        ram_buffer(28489) := X"00000000";
        ram_buffer(28490) := X"AC400010";
        ram_buffer(28491) := X"8FC20018";
        ram_buffer(28492) := X"00000000";
        ram_buffer(28493) := X"AC400014";
        ram_buffer(28494) := X"8FC20018";
        ram_buffer(28495) := X"00000000";
        ram_buffer(28496) := X"AC400018";
        ram_buffer(28497) := X"8FC20018";
        ram_buffer(28498) := X"00000000";
        ram_buffer(28499) := X"2442005C";
        ram_buffer(28500) := X"24060008";
        ram_buffer(28501) := X"00002821";
        ram_buffer(28502) := X"00402021";
        ram_buffer(28503) := X"0C02801D";
        ram_buffer(28504) := X"00000000";
        ram_buffer(28505) := X"8FC20018";
        ram_buffer(28506) := X"8FC30018";
        ram_buffer(28507) := X"00000000";
        ram_buffer(28508) := X"AC43001C";
        ram_buffer(28509) := X"8FC20018";
        ram_buffer(28510) := X"3C03100A";
        ram_buffer(28511) := X"246311A8";
        ram_buffer(28512) := X"AC430020";
        ram_buffer(28513) := X"8FC20018";
        ram_buffer(28514) := X"3C03100A";
        ram_buffer(28515) := X"24631298";
        ram_buffer(28516) := X"AC430024";
        ram_buffer(28517) := X"8FC20018";
        ram_buffer(28518) := X"3C03100A";
        ram_buffer(28519) := X"24631360";
        ram_buffer(28520) := X"AC430028";
        ram_buffer(28521) := X"8FC20018";
        ram_buffer(28522) := X"3C03100A";
        ram_buffer(28523) := X"2463141C";
        ram_buffer(28524) := X"AC43002C";
        ram_buffer(28525) := X"00000000";
        ram_buffer(28526) := X"03C0E821";
        ram_buffer(28527) := X"8FBF0014";
        ram_buffer(28528) := X"8FBE0010";
        ram_buffer(28529) := X"27BD0018";
        ram_buffer(28530) := X"03E00008";
        ram_buffer(28531) := X"00000000";
        ram_buffer(28532) := X"27BDFFD8";
        ram_buffer(28533) := X"AFBF0024";
        ram_buffer(28534) := X"AFBE0020";
        ram_buffer(28535) := X"AFB0001C";
        ram_buffer(28536) := X"03A0F021";
        ram_buffer(28537) := X"AFC40028";
        ram_buffer(28538) := X"00A08021";
        ram_buffer(28539) := X"2602FFFF";
        ram_buffer(28540) := X"00402021";
        ram_buffer(28541) := X"00801821";
        ram_buffer(28542) := X"00031080";
        ram_buffer(28543) := X"00401821";
        ram_buffer(28544) := X"00031080";
        ram_buffer(28545) := X"00431023";
        ram_buffer(28546) := X"00441021";
        ram_buffer(28547) := X"000210C0";
        ram_buffer(28548) := X"24420074";
        ram_buffer(28549) := X"00402821";
        ram_buffer(28550) := X"8FC40028";
        ram_buffer(28551) := X"0C027B8F";
        ram_buffer(28552) := X"00000000";
        ram_buffer(28553) := X"AFC20010";
        ram_buffer(28554) := X"8FC20010";
        ram_buffer(28555) := X"00000000";
        ram_buffer(28556) := X"14400004";
        ram_buffer(28557) := X"00000000";
        ram_buffer(28558) := X"00001021";
        ram_buffer(28559) := X"1000001E";
        ram_buffer(28560) := X"00000000";
        ram_buffer(28561) := X"8FC20010";
        ram_buffer(28562) := X"00000000";
        ram_buffer(28563) := X"AC400000";
        ram_buffer(28564) := X"8FC20010";
        ram_buffer(28565) := X"00000000";
        ram_buffer(28566) := X"AC500004";
        ram_buffer(28567) := X"8FC20010";
        ram_buffer(28568) := X"00000000";
        ram_buffer(28569) := X"2443000C";
        ram_buffer(28570) := X"8FC20010";
        ram_buffer(28571) := X"00000000";
        ram_buffer(28572) := X"AC430008";
        ram_buffer(28573) := X"8FC20010";
        ram_buffer(28574) := X"00000000";
        ram_buffer(28575) := X"2447000C";
        ram_buffer(28576) := X"02002021";
        ram_buffer(28577) := X"00801821";
        ram_buffer(28578) := X"00031080";
        ram_buffer(28579) := X"00401821";
        ram_buffer(28580) := X"00031080";
        ram_buffer(28581) := X"00431023";
        ram_buffer(28582) := X"00441021";
        ram_buffer(28583) := X"000210C0";
        ram_buffer(28584) := X"00403021";
        ram_buffer(28585) := X"00002821";
        ram_buffer(28586) := X"00E02021";
        ram_buffer(28587) := X"0C02801D";
        ram_buffer(28588) := X"00000000";
        ram_buffer(28589) := X"8FC20010";
        ram_buffer(28590) := X"03C0E821";
        ram_buffer(28591) := X"8FBF0024";
        ram_buffer(28592) := X"8FBE0020";
        ram_buffer(28593) := X"8FB0001C";
        ram_buffer(28594) := X"27BD0028";
        ram_buffer(28595) := X"03E00008";
        ram_buffer(28596) := X"00000000";
        ram_buffer(28597) := X"27BDFFD8";
        ram_buffer(28598) := X"AFBF0024";
        ram_buffer(28599) := X"AFBE0020";
        ram_buffer(28600) := X"03A0F021";
        ram_buffer(28601) := X"AFC40028";
        ram_buffer(28602) := X"0C0270B0";
        ram_buffer(28603) := X"00000000";
        ram_buffer(28604) := X"8F82809C";
        ram_buffer(28605) := X"00000000";
        ram_buffer(28606) := X"8C420038";
        ram_buffer(28607) := X"00000000";
        ram_buffer(28608) := X"14400006";
        ram_buffer(28609) := X"00000000";
        ram_buffer(28610) := X"8F82809C";
        ram_buffer(28611) := X"00000000";
        ram_buffer(28612) := X"00402021";
        ram_buffer(28613) := X"0C027069";
        ram_buffer(28614) := X"00000000";
        ram_buffer(28615) := X"8F82809C";
        ram_buffer(28616) := X"00000000";
        ram_buffer(28617) := X"244202E0";
        ram_buffer(28618) := X"AFC20018";
        ram_buffer(28619) := X"8FC20018";
        ram_buffer(28620) := X"00000000";
        ram_buffer(28621) := X"8C420008";
        ram_buffer(28622) := X"00000000";
        ram_buffer(28623) := X"AFC20010";
        ram_buffer(28624) := X"8FC20018";
        ram_buffer(28625) := X"00000000";
        ram_buffer(28626) := X"8C420004";
        ram_buffer(28627) := X"00000000";
        ram_buffer(28628) := X"AFC20014";
        ram_buffer(28629) := X"1000000B";
        ram_buffer(28630) := X"00000000";
        ram_buffer(28631) := X"8FC20010";
        ram_buffer(28632) := X"00000000";
        ram_buffer(28633) := X"8442000C";
        ram_buffer(28634) := X"00000000";
        ram_buffer(28635) := X"10400031";
        ram_buffer(28636) := X"00000000";
        ram_buffer(28637) := X"8FC20010";
        ram_buffer(28638) := X"00000000";
        ram_buffer(28639) := X"24420068";
        ram_buffer(28640) := X"AFC20010";
        ram_buffer(28641) := X"8FC20014";
        ram_buffer(28642) := X"00000000";
        ram_buffer(28643) := X"2442FFFF";
        ram_buffer(28644) := X"AFC20014";
        ram_buffer(28645) := X"8FC20014";
        ram_buffer(28646) := X"00000000";
        ram_buffer(28647) := X"0441FFEF";
        ram_buffer(28648) := X"00000000";
        ram_buffer(28649) := X"8FC20018";
        ram_buffer(28650) := X"00000000";
        ram_buffer(28651) := X"8C420000";
        ram_buffer(28652) := X"00000000";
        ram_buffer(28653) := X"1440000F";
        ram_buffer(28654) := X"00000000";
        ram_buffer(28655) := X"24050004";
        ram_buffer(28656) := X"8FC40028";
        ram_buffer(28657) := X"0C026F74";
        ram_buffer(28658) := X"00000000";
        ram_buffer(28659) := X"00401821";
        ram_buffer(28660) := X"8FC20018";
        ram_buffer(28661) := X"00000000";
        ram_buffer(28662) := X"AC430000";
        ram_buffer(28663) := X"8FC20018";
        ram_buffer(28664) := X"00000000";
        ram_buffer(28665) := X"8C420000";
        ram_buffer(28666) := X"00000000";
        ram_buffer(28667) := X"10400008";
        ram_buffer(28668) := X"00000000";
        ram_buffer(28669) := X"8FC20018";
        ram_buffer(28670) := X"00000000";
        ram_buffer(28671) := X"8C420000";
        ram_buffer(28672) := X"00000000";
        ram_buffer(28673) := X"AFC20018";
        ram_buffer(28674) := X"1000FFC8";
        ram_buffer(28675) := X"00000000";
        ram_buffer(28676) := X"00000000";
        ram_buffer(28677) := X"0C0270B9";
        ram_buffer(28678) := X"00000000";
        ram_buffer(28679) := X"8FC20028";
        ram_buffer(28680) := X"2403000C";
        ram_buffer(28681) := X"AC430000";
        ram_buffer(28682) := X"00001021";
        ram_buffer(28683) := X"10000034";
        ram_buffer(28684) := X"00000000";
        ram_buffer(28685) := X"00000000";
        ram_buffer(28686) := X"8FC20010";
        ram_buffer(28687) := X"2403FFFF";
        ram_buffer(28688) := X"A443000E";
        ram_buffer(28689) := X"8FC20010";
        ram_buffer(28690) := X"24030001";
        ram_buffer(28691) := X"A443000C";
        ram_buffer(28692) := X"8FC20010";
        ram_buffer(28693) := X"00000000";
        ram_buffer(28694) := X"AC400064";
        ram_buffer(28695) := X"0C0270B9";
        ram_buffer(28696) := X"00000000";
        ram_buffer(28697) := X"8FC20010";
        ram_buffer(28698) := X"00000000";
        ram_buffer(28699) := X"AC400000";
        ram_buffer(28700) := X"8FC20010";
        ram_buffer(28701) := X"00000000";
        ram_buffer(28702) := X"AC400008";
        ram_buffer(28703) := X"8FC20010";
        ram_buffer(28704) := X"00000000";
        ram_buffer(28705) := X"AC400004";
        ram_buffer(28706) := X"8FC20010";
        ram_buffer(28707) := X"00000000";
        ram_buffer(28708) := X"AC400010";
        ram_buffer(28709) := X"8FC20010";
        ram_buffer(28710) := X"00000000";
        ram_buffer(28711) := X"AC400014";
        ram_buffer(28712) := X"8FC20010";
        ram_buffer(28713) := X"00000000";
        ram_buffer(28714) := X"AC400018";
        ram_buffer(28715) := X"8FC20010";
        ram_buffer(28716) := X"00000000";
        ram_buffer(28717) := X"2442005C";
        ram_buffer(28718) := X"24060008";
        ram_buffer(28719) := X"00002821";
        ram_buffer(28720) := X"00402021";
        ram_buffer(28721) := X"0C02801D";
        ram_buffer(28722) := X"00000000";
        ram_buffer(28723) := X"8FC20010";
        ram_buffer(28724) := X"00000000";
        ram_buffer(28725) := X"AC400030";
        ram_buffer(28726) := X"8FC20010";
        ram_buffer(28727) := X"00000000";
        ram_buffer(28728) := X"AC400034";
        ram_buffer(28729) := X"8FC20010";
        ram_buffer(28730) := X"00000000";
        ram_buffer(28731) := X"AC400044";
        ram_buffer(28732) := X"8FC20010";
        ram_buffer(28733) := X"00000000";
        ram_buffer(28734) := X"AC400048";
        ram_buffer(28735) := X"8FC20010";
        ram_buffer(28736) := X"03C0E821";
        ram_buffer(28737) := X"8FBF0024";
        ram_buffer(28738) := X"8FBE0020";
        ram_buffer(28739) := X"27BD0028";
        ram_buffer(28740) := X"03E00008";
        ram_buffer(28741) := X"00000000";
        ram_buffer(28742) := X"27BDFFE0";
        ram_buffer(28743) := X"AFBF001C";
        ram_buffer(28744) := X"AFBE0018";
        ram_buffer(28745) := X"03A0F021";
        ram_buffer(28746) := X"AFC40020";
        ram_buffer(28747) := X"3C02100A";
        ram_buffer(28748) := X"2442B544";
        ram_buffer(28749) := X"AFC20010";
        ram_buffer(28750) := X"8FC50010";
        ram_buffer(28751) := X"8FC40020";
        ram_buffer(28752) := X"0C02783C";
        ram_buffer(28753) := X"00000000";
        ram_buffer(28754) := X"00000000";
        ram_buffer(28755) := X"03C0E821";
        ram_buffer(28756) := X"8FBF001C";
        ram_buffer(28757) := X"8FBE0018";
        ram_buffer(28758) := X"27BD0020";
        ram_buffer(28759) := X"03E00008";
        ram_buffer(28760) := X"00000000";
        ram_buffer(28761) := X"27BDFFE8";
        ram_buffer(28762) := X"AFBF0014";
        ram_buffer(28763) := X"AFBE0010";
        ram_buffer(28764) := X"03A0F021";
        ram_buffer(28765) := X"8F82809C";
        ram_buffer(28766) := X"00000000";
        ram_buffer(28767) := X"00402021";
        ram_buffer(28768) := X"0C027046";
        ram_buffer(28769) := X"00000000";
        ram_buffer(28770) := X"00000000";
        ram_buffer(28771) := X"03C0E821";
        ram_buffer(28772) := X"8FBF0014";
        ram_buffer(28773) := X"8FBE0010";
        ram_buffer(28774) := X"27BD0018";
        ram_buffer(28775) := X"03E00008";
        ram_buffer(28776) := X"00000000";
        ram_buffer(28777) := X"27BDFFE8";
        ram_buffer(28778) := X"AFBF0014";
        ram_buffer(28779) := X"AFBE0010";
        ram_buffer(28780) := X"03A0F021";
        ram_buffer(28781) := X"AFC40018";
        ram_buffer(28782) := X"0C0270C2";
        ram_buffer(28783) := X"00000000";
        ram_buffer(28784) := X"8FC20018";
        ram_buffer(28785) := X"00000000";
        ram_buffer(28786) := X"8C420038";
        ram_buffer(28787) := X"00000000";
        ram_buffer(28788) := X"10400005";
        ram_buffer(28789) := X"00000000";
        ram_buffer(28790) := X"0C0270CB";
        ram_buffer(28791) := X"00000000";
        ram_buffer(28792) := X"10000031";
        ram_buffer(28793) := X"00000000";
        ram_buffer(28794) := X"8FC20018";
        ram_buffer(28795) := X"3C03100A";
        ram_buffer(28796) := X"2463C118";
        ram_buffer(28797) := X"AC43003C";
        ram_buffer(28798) := X"8FC20018";
        ram_buffer(28799) := X"00000000";
        ram_buffer(28800) := X"AC4002E0";
        ram_buffer(28801) := X"8FC20018";
        ram_buffer(28802) := X"24030003";
        ram_buffer(28803) := X"AC4302E4";
        ram_buffer(28804) := X"8FC20018";
        ram_buffer(28805) := X"00000000";
        ram_buffer(28806) := X"244302EC";
        ram_buffer(28807) := X"8FC20018";
        ram_buffer(28808) := X"00000000";
        ram_buffer(28809) := X"AC4302E8";
        ram_buffer(28810) := X"8FC20018";
        ram_buffer(28811) := X"00000000";
        ram_buffer(28812) := X"8C420004";
        ram_buffer(28813) := X"8FC70018";
        ram_buffer(28814) := X"00003021";
        ram_buffer(28815) := X"24050004";
        ram_buffer(28816) := X"00402021";
        ram_buffer(28817) := X"0C026F26";
        ram_buffer(28818) := X"00000000";
        ram_buffer(28819) := X"8FC20018";
        ram_buffer(28820) := X"00000000";
        ram_buffer(28821) := X"8C420008";
        ram_buffer(28822) := X"8FC70018";
        ram_buffer(28823) := X"24060001";
        ram_buffer(28824) := X"24050009";
        ram_buffer(28825) := X"00402021";
        ram_buffer(28826) := X"0C026F26";
        ram_buffer(28827) := X"00000000";
        ram_buffer(28828) := X"8FC20018";
        ram_buffer(28829) := X"00000000";
        ram_buffer(28830) := X"8C42000C";
        ram_buffer(28831) := X"8FC70018";
        ram_buffer(28832) := X"24060002";
        ram_buffer(28833) := X"24050012";
        ram_buffer(28834) := X"00402021";
        ram_buffer(28835) := X"0C026F26";
        ram_buffer(28836) := X"00000000";
        ram_buffer(28837) := X"8FC20018";
        ram_buffer(28838) := X"24030001";
        ram_buffer(28839) := X"AC430038";
        ram_buffer(28840) := X"0C0270CB";
        ram_buffer(28841) := X"00000000";
        ram_buffer(28842) := X"03C0E821";
        ram_buffer(28843) := X"8FBF0014";
        ram_buffer(28844) := X"8FBE0010";
        ram_buffer(28845) := X"27BD0018";
        ram_buffer(28846) := X"03E00008";
        ram_buffer(28847) := X"00000000";
        ram_buffer(28848) := X"27BDFFF8";
        ram_buffer(28849) := X"AFBE0004";
        ram_buffer(28850) := X"03A0F021";
        ram_buffer(28851) := X"00000000";
        ram_buffer(28852) := X"03C0E821";
        ram_buffer(28853) := X"8FBE0004";
        ram_buffer(28854) := X"27BD0008";
        ram_buffer(28855) := X"03E00008";
        ram_buffer(28856) := X"00000000";
        ram_buffer(28857) := X"27BDFFF8";
        ram_buffer(28858) := X"AFBE0004";
        ram_buffer(28859) := X"03A0F021";
        ram_buffer(28860) := X"00000000";
        ram_buffer(28861) := X"03C0E821";
        ram_buffer(28862) := X"8FBE0004";
        ram_buffer(28863) := X"27BD0008";
        ram_buffer(28864) := X"03E00008";
        ram_buffer(28865) := X"00000000";
        ram_buffer(28866) := X"27BDFFF8";
        ram_buffer(28867) := X"AFBE0004";
        ram_buffer(28868) := X"03A0F021";
        ram_buffer(28869) := X"00000000";
        ram_buffer(28870) := X"03C0E821";
        ram_buffer(28871) := X"8FBE0004";
        ram_buffer(28872) := X"27BD0008";
        ram_buffer(28873) := X"03E00008";
        ram_buffer(28874) := X"00000000";
        ram_buffer(28875) := X"27BDFFF8";
        ram_buffer(28876) := X"AFBE0004";
        ram_buffer(28877) := X"03A0F021";
        ram_buffer(28878) := X"00000000";
        ram_buffer(28879) := X"03C0E821";
        ram_buffer(28880) := X"8FBE0004";
        ram_buffer(28881) := X"27BD0008";
        ram_buffer(28882) := X"03E00008";
        ram_buffer(28883) := X"00000000";
        ram_buffer(28884) := X"27BDFFF8";
        ram_buffer(28885) := X"AFBE0004";
        ram_buffer(28886) := X"03A0F021";
        ram_buffer(28887) := X"AFC40008";
        ram_buffer(28888) := X"00001021";
        ram_buffer(28889) := X"03C0E821";
        ram_buffer(28890) := X"8FBE0004";
        ram_buffer(28891) := X"27BD0008";
        ram_buffer(28892) := X"03E00008";
        ram_buffer(28893) := X"00000000";
        ram_buffer(28894) := X"27BDFFF8";
        ram_buffer(28895) := X"AFBE0004";
        ram_buffer(28896) := X"03A0F021";
        ram_buffer(28897) := X"AFC40008";
        ram_buffer(28898) := X"00001021";
        ram_buffer(28899) := X"03C0E821";
        ram_buffer(28900) := X"8FBE0004";
        ram_buffer(28901) := X"27BD0008";
        ram_buffer(28902) := X"03E00008";
        ram_buffer(28903) := X"00000000";
        ram_buffer(28904) := X"27BDFFE8";
        ram_buffer(28905) := X"AFBF0014";
        ram_buffer(28906) := X"AFBE0010";
        ram_buffer(28907) := X"03A0F021";
        ram_buffer(28908) := X"0C0270B0";
        ram_buffer(28909) := X"00000000";
        ram_buffer(28910) := X"8F838098";
        ram_buffer(28911) := X"3C02100A";
        ram_buffer(28912) := X"2445C350";
        ram_buffer(28913) := X"00602021";
        ram_buffer(28914) := X"0C027803";
        ram_buffer(28915) := X"00000000";
        ram_buffer(28916) := X"00000000";
        ram_buffer(28917) := X"03C0E821";
        ram_buffer(28918) := X"8FBF0014";
        ram_buffer(28919) := X"8FBE0010";
        ram_buffer(28920) := X"27BD0018";
        ram_buffer(28921) := X"03E00008";
        ram_buffer(28922) := X"00000000";
        ram_buffer(28923) := X"27BDFFE8";
        ram_buffer(28924) := X"AFBF0014";
        ram_buffer(28925) := X"AFBE0010";
        ram_buffer(28926) := X"03A0F021";
        ram_buffer(28927) := X"8F838098";
        ram_buffer(28928) := X"3C02100A";
        ram_buffer(28929) := X"2445C378";
        ram_buffer(28930) := X"00602021";
        ram_buffer(28931) := X"0C027803";
        ram_buffer(28932) := X"00000000";
        ram_buffer(28933) := X"0C0270B9";
        ram_buffer(28934) := X"00000000";
        ram_buffer(28935) := X"00000000";
        ram_buffer(28936) := X"03C0E821";
        ram_buffer(28937) := X"8FBF0014";
        ram_buffer(28938) := X"8FBE0010";
        ram_buffer(28939) := X"27BD0018";
        ram_buffer(28940) := X"03E00008";
        ram_buffer(28941) := X"00000000";
        ram_buffer(28942) := X"27BDFFD8";
        ram_buffer(28943) := X"AFBF0024";
        ram_buffer(28944) := X"AFBE0020";
        ram_buffer(28945) := X"AFB1001C";
        ram_buffer(28946) := X"AFB00018";
        ram_buffer(28947) := X"03A0F021";
        ram_buffer(28948) := X"AFC40028";
        ram_buffer(28949) := X"AFC5002C";
        ram_buffer(28950) := X"AFC60030";
        ram_buffer(28951) := X"27C20014";
        ram_buffer(28952) := X"00403021";
        ram_buffer(28953) := X"8FC50030";
        ram_buffer(28954) := X"8FC40028";
        ram_buffer(28955) := X"0C02B846";
        ram_buffer(28956) := X"00000000";
        ram_buffer(28957) := X"AFC20010";
        ram_buffer(28958) := X"8FC20010";
        ram_buffer(28959) := X"00000000";
        ram_buffer(28960) := X"14400004";
        ram_buffer(28961) := X"00000000";
        ram_buffer(28962) := X"00001021";
        ram_buffer(28963) := X"1000003E";
        ram_buffer(28964) := X"00000000";
        ram_buffer(28965) := X"8FC40028";
        ram_buffer(28966) := X"0C026FB5";
        ram_buffer(28967) := X"00000000";
        ram_buffer(28968) := X"00408021";
        ram_buffer(28969) := X"16000004";
        ram_buffer(28970) := X"00000000";
        ram_buffer(28971) := X"00001021";
        ram_buffer(28972) := X"10000035";
        ram_buffer(28973) := X"00000000";
        ram_buffer(28974) := X"8FC20014";
        ram_buffer(28975) := X"240701B6";
        ram_buffer(28976) := X"00403021";
        ram_buffer(28977) := X"8FC5002C";
        ram_buffer(28978) := X"8FC40028";
        ram_buffer(28979) := X"0C0280D7";
        ram_buffer(28980) := X"00000000";
        ram_buffer(28981) := X"00408821";
        ram_buffer(28982) := X"06210009";
        ram_buffer(28983) := X"00000000";
        ram_buffer(28984) := X"0C0270B0";
        ram_buffer(28985) := X"00000000";
        ram_buffer(28986) := X"A600000C";
        ram_buffer(28987) := X"0C0270B9";
        ram_buffer(28988) := X"00000000";
        ram_buffer(28989) := X"00001021";
        ram_buffer(28990) := X"10000023";
        ram_buffer(28991) := X"00000000";
        ram_buffer(28992) := X"00111400";
        ram_buffer(28993) := X"00021403";
        ram_buffer(28994) := X"A602000E";
        ram_buffer(28995) := X"8FC20010";
        ram_buffer(28996) := X"00000000";
        ram_buffer(28997) := X"00021400";
        ram_buffer(28998) := X"00021403";
        ram_buffer(28999) := X"A602000C";
        ram_buffer(29000) := X"AE10001C";
        ram_buffer(29001) := X"3C02100A";
        ram_buffer(29002) := X"244211A8";
        ram_buffer(29003) := X"AE020020";
        ram_buffer(29004) := X"3C02100A";
        ram_buffer(29005) := X"24421298";
        ram_buffer(29006) := X"AE020024";
        ram_buffer(29007) := X"3C02100A";
        ram_buffer(29008) := X"24421360";
        ram_buffer(29009) := X"AE020028";
        ram_buffer(29010) := X"3C02100A";
        ram_buffer(29011) := X"2442141C";
        ram_buffer(29012) := X"AE02002C";
        ram_buffer(29013) := X"8602000C";
        ram_buffer(29014) := X"00000000";
        ram_buffer(29015) := X"3042FFFF";
        ram_buffer(29016) := X"30420100";
        ram_buffer(29017) := X"10400007";
        ram_buffer(29018) := X"00000000";
        ram_buffer(29019) := X"24070002";
        ram_buffer(29020) := X"00003021";
        ram_buffer(29021) := X"02002821";
        ram_buffer(29022) := X"8FC40028";
        ram_buffer(29023) := X"0C027579";
        ram_buffer(29024) := X"00000000";
        ram_buffer(29025) := X"02001021";
        ram_buffer(29026) := X"03C0E821";
        ram_buffer(29027) := X"8FBF0024";
        ram_buffer(29028) := X"8FBE0020";
        ram_buffer(29029) := X"8FB1001C";
        ram_buffer(29030) := X"8FB00018";
        ram_buffer(29031) := X"27BD0028";
        ram_buffer(29032) := X"03E00008";
        ram_buffer(29033) := X"00000000";
        ram_buffer(29034) := X"27BDFFE8";
        ram_buffer(29035) := X"AFBF0014";
        ram_buffer(29036) := X"AFBE0010";
        ram_buffer(29037) := X"03A0F021";
        ram_buffer(29038) := X"AFC40018";
        ram_buffer(29039) := X"AFC5001C";
        ram_buffer(29040) := X"8F828098";
        ram_buffer(29041) := X"8FC6001C";
        ram_buffer(29042) := X"8FC50018";
        ram_buffer(29043) := X"00402021";
        ram_buffer(29044) := X"0C02710E";
        ram_buffer(29045) := X"00000000";
        ram_buffer(29046) := X"03C0E821";
        ram_buffer(29047) := X"8FBF0014";
        ram_buffer(29048) := X"8FBE0010";
        ram_buffer(29049) := X"27BD0018";
        ram_buffer(29050) := X"03E00008";
        ram_buffer(29051) := X"00000000";
        ram_buffer(29052) := X"27BDFFE0";
        ram_buffer(29053) := X"AFBF001C";
        ram_buffer(29054) := X"AFBE0018";
        ram_buffer(29055) := X"03A0F021";
        ram_buffer(29056) := X"AFC40020";
        ram_buffer(29057) := X"AFC50024";
        ram_buffer(29058) := X"AFC60028";
        ram_buffer(29059) := X"AFC7002C";
        ram_buffer(29060) := X"27C2002C";
        ram_buffer(29061) := X"AFC20014";
        ram_buffer(29062) := X"8FC20014";
        ram_buffer(29063) := X"00000000";
        ram_buffer(29064) := X"00403821";
        ram_buffer(29065) := X"8FC60028";
        ram_buffer(29066) := X"8FC50024";
        ram_buffer(29067) := X"8FC40020";
        ram_buffer(29068) := X"0C029DFA";
        ram_buffer(29069) := X"00000000";
        ram_buffer(29070) := X"AFC20010";
        ram_buffer(29071) := X"8FC20010";
        ram_buffer(29072) := X"03C0E821";
        ram_buffer(29073) := X"8FBF001C";
        ram_buffer(29074) := X"8FBE0018";
        ram_buffer(29075) := X"27BD0020";
        ram_buffer(29076) := X"03E00008";
        ram_buffer(29077) := X"00000000";
        ram_buffer(29078) := X"27BDFFE0";
        ram_buffer(29079) := X"AFBF001C";
        ram_buffer(29080) := X"AFBE0018";
        ram_buffer(29081) := X"03A0F021";
        ram_buffer(29082) := X"AFC40020";
        ram_buffer(29083) := X"AFC50024";
        ram_buffer(29084) := X"AFC60028";
        ram_buffer(29085) := X"AFC7002C";
        ram_buffer(29086) := X"27C20028";
        ram_buffer(29087) := X"AFC20014";
        ram_buffer(29088) := X"8F828098";
        ram_buffer(29089) := X"8FC30014";
        ram_buffer(29090) := X"00000000";
        ram_buffer(29091) := X"00603821";
        ram_buffer(29092) := X"8FC60024";
        ram_buffer(29093) := X"8FC50020";
        ram_buffer(29094) := X"00402021";
        ram_buffer(29095) := X"0C029DFA";
        ram_buffer(29096) := X"00000000";
        ram_buffer(29097) := X"AFC20010";
        ram_buffer(29098) := X"8FC20010";
        ram_buffer(29099) := X"03C0E821";
        ram_buffer(29100) := X"8FBF001C";
        ram_buffer(29101) := X"8FBE0018";
        ram_buffer(29102) := X"27BD0020";
        ram_buffer(29103) := X"03E00008";
        ram_buffer(29104) := X"00000000";
        ram_buffer(29105) := X"27BDFFB8";
        ram_buffer(29106) := X"AFBF0044";
        ram_buffer(29107) := X"AFBE0040";
        ram_buffer(29108) := X"AFB2003C";
        ram_buffer(29109) := X"AFB10038";
        ram_buffer(29110) := X"AFB00034";
        ram_buffer(29111) := X"03A0F021";
        ram_buffer(29112) := X"AFC40048";
        ram_buffer(29113) := X"AFC5004C";
        ram_buffer(29114) := X"AFC60050";
        ram_buffer(29115) := X"AFC70054";
        ram_buffer(29116) := X"8FC30054";
        ram_buffer(29117) := X"8FC20050";
        ram_buffer(29118) := X"00000000";
        ram_buffer(29119) := X"00620018";
        ram_buffer(29120) := X"00008012";
        ram_buffer(29121) := X"16000004";
        ram_buffer(29122) := X"00000000";
        ram_buffer(29123) := X"00001021";
        ram_buffer(29124) := X"1000011B";
        ram_buffer(29125) := X"00000000";
        ram_buffer(29126) := X"8FC20048";
        ram_buffer(29127) := X"00000000";
        ram_buffer(29128) := X"AFC20010";
        ram_buffer(29129) := X"8FC20010";
        ram_buffer(29130) := X"00000000";
        ram_buffer(29131) := X"1040000A";
        ram_buffer(29132) := X"00000000";
        ram_buffer(29133) := X"8FC20010";
        ram_buffer(29134) := X"00000000";
        ram_buffer(29135) := X"8C420038";
        ram_buffer(29136) := X"00000000";
        ram_buffer(29137) := X"14400004";
        ram_buffer(29138) := X"00000000";
        ram_buffer(29139) := X"8FC40010";
        ram_buffer(29140) := X"0C027069";
        ram_buffer(29141) := X"00000000";
        ram_buffer(29142) := X"8FC20058";
        ram_buffer(29143) := X"00000000";
        ram_buffer(29144) := X"8442000C";
        ram_buffer(29145) := X"00000000";
        ram_buffer(29146) := X"3042FFFF";
        ram_buffer(29147) := X"30422000";
        ram_buffer(29148) := X"14400013";
        ram_buffer(29149) := X"00000000";
        ram_buffer(29150) := X"8FC20058";
        ram_buffer(29151) := X"00000000";
        ram_buffer(29152) := X"8442000C";
        ram_buffer(29153) := X"00000000";
        ram_buffer(29154) := X"34422000";
        ram_buffer(29155) := X"00021C00";
        ram_buffer(29156) := X"00031C03";
        ram_buffer(29157) := X"8FC20058";
        ram_buffer(29158) := X"00000000";
        ram_buffer(29159) := X"A443000C";
        ram_buffer(29160) := X"8FC20058";
        ram_buffer(29161) := X"00000000";
        ram_buffer(29162) := X"8C430064";
        ram_buffer(29163) := X"2402DFFF";
        ram_buffer(29164) := X"00621824";
        ram_buffer(29165) := X"8FC20058";
        ram_buffer(29166) := X"00000000";
        ram_buffer(29167) := X"AC430064";
        ram_buffer(29168) := X"8FC20058";
        ram_buffer(29169) := X"00000000";
        ram_buffer(29170) := X"8C420004";
        ram_buffer(29171) := X"00000000";
        ram_buffer(29172) := X"04410004";
        ram_buffer(29173) := X"00000000";
        ram_buffer(29174) := X"8FC20058";
        ram_buffer(29175) := X"00000000";
        ram_buffer(29176) := X"AC400004";
        ram_buffer(29177) := X"AFD00014";
        ram_buffer(29178) := X"8FD1004C";
        ram_buffer(29179) := X"8FC20058";
        ram_buffer(29180) := X"00000000";
        ram_buffer(29181) := X"8442000C";
        ram_buffer(29182) := X"00000000";
        ram_buffer(29183) := X"3042FFFF";
        ram_buffer(29184) := X"30420002";
        ram_buffer(29185) := X"104000BC";
        ram_buffer(29186) := X"00000000";
        ram_buffer(29187) := X"8FC20058";
        ram_buffer(29188) := X"00000000";
        ram_buffer(29189) := X"8C420004";
        ram_buffer(29190) := X"00000000";
        ram_buffer(29191) := X"0202182B";
        ram_buffer(29192) := X"10600002";
        ram_buffer(29193) := X"00000000";
        ram_buffer(29194) := X"02001021";
        ram_buffer(29195) := X"AFC20018";
        ram_buffer(29196) := X"8FC20058";
        ram_buffer(29197) := X"00000000";
        ram_buffer(29198) := X"8C420000";
        ram_buffer(29199) := X"8FC30018";
        ram_buffer(29200) := X"00000000";
        ram_buffer(29201) := X"00603021";
        ram_buffer(29202) := X"00402821";
        ram_buffer(29203) := X"02202021";
        ram_buffer(29204) := X"0C027F93";
        ram_buffer(29205) := X"00000000";
        ram_buffer(29206) := X"8FC20058";
        ram_buffer(29207) := X"00000000";
        ram_buffer(29208) := X"8C430000";
        ram_buffer(29209) := X"8FC20018";
        ram_buffer(29210) := X"00000000";
        ram_buffer(29211) := X"00621821";
        ram_buffer(29212) := X"8FC20058";
        ram_buffer(29213) := X"00000000";
        ram_buffer(29214) := X"AC430000";
        ram_buffer(29215) := X"8FC20058";
        ram_buffer(29216) := X"00000000";
        ram_buffer(29217) := X"8C430004";
        ram_buffer(29218) := X"8FC20018";
        ram_buffer(29219) := X"00000000";
        ram_buffer(29220) := X"00621823";
        ram_buffer(29221) := X"8FC20058";
        ram_buffer(29222) := X"00000000";
        ram_buffer(29223) := X"AC430004";
        ram_buffer(29224) := X"8FC20018";
        ram_buffer(29225) := X"00000000";
        ram_buffer(29226) := X"02228821";
        ram_buffer(29227) := X"8FC20018";
        ram_buffer(29228) := X"00000000";
        ram_buffer(29229) := X"02028023";
        ram_buffer(29230) := X"8FC20058";
        ram_buffer(29231) := X"00000000";
        ram_buffer(29232) := X"8C420030";
        ram_buffer(29233) := X"00000000";
        ram_buffer(29234) := X"10400060";
        ram_buffer(29235) := X"00000000";
        ram_buffer(29236) := X"1200005E";
        ram_buffer(29237) := X"00000000";
        ram_buffer(29238) := X"8FC20058";
        ram_buffer(29239) := X"00000000";
        ram_buffer(29240) := X"8C430030";
        ram_buffer(29241) := X"8FC20058";
        ram_buffer(29242) := X"00000000";
        ram_buffer(29243) := X"24420040";
        ram_buffer(29244) := X"10620009";
        ram_buffer(29245) := X"00000000";
        ram_buffer(29246) := X"8FC20058";
        ram_buffer(29247) := X"00000000";
        ram_buffer(29248) := X"8C420030";
        ram_buffer(29249) := X"00000000";
        ram_buffer(29250) := X"00402821";
        ram_buffer(29251) := X"8FC40048";
        ram_buffer(29252) := X"0C027301";
        ram_buffer(29253) := X"00000000";
        ram_buffer(29254) := X"8FC20058";
        ram_buffer(29255) := X"00000000";
        ram_buffer(29256) := X"AC400030";
        ram_buffer(29257) := X"10000049";
        ram_buffer(29258) := X"00000000";
        ram_buffer(29259) := X"AFC0001C";
        ram_buffer(29260) := X"8FC20058";
        ram_buffer(29261) := X"00000000";
        ram_buffer(29262) := X"8C420010";
        ram_buffer(29263) := X"00000000";
        ram_buffer(29264) := X"AFC20020";
        ram_buffer(29265) := X"8FC20058";
        ram_buffer(29266) := X"00000000";
        ram_buffer(29267) := X"8C420000";
        ram_buffer(29268) := X"00000000";
        ram_buffer(29269) := X"AFC20024";
        ram_buffer(29270) := X"8FC20058";
        ram_buffer(29271) := X"00000000";
        ram_buffer(29272) := X"8C420014";
        ram_buffer(29273) := X"00000000";
        ram_buffer(29274) := X"AFC20028";
        ram_buffer(29275) := X"8FC20058";
        ram_buffer(29276) := X"00000000";
        ram_buffer(29277) := X"AC510010";
        ram_buffer(29278) := X"02001821";
        ram_buffer(29279) := X"8FC20058";
        ram_buffer(29280) := X"00000000";
        ram_buffer(29281) := X"AC430014";
        ram_buffer(29282) := X"8FC20058";
        ram_buffer(29283) := X"00000000";
        ram_buffer(29284) := X"AC510000";
        ram_buffer(29285) := X"8FC50058";
        ram_buffer(29286) := X"8FC40048";
        ram_buffer(29287) := X"0C028274";
        ram_buffer(29288) := X"00000000";
        ram_buffer(29289) := X"AFC2001C";
        ram_buffer(29290) := X"8FC20058";
        ram_buffer(29291) := X"8FC30020";
        ram_buffer(29292) := X"00000000";
        ram_buffer(29293) := X"AC430010";
        ram_buffer(29294) := X"8FC20058";
        ram_buffer(29295) := X"8FC30028";
        ram_buffer(29296) := X"00000000";
        ram_buffer(29297) := X"AC430014";
        ram_buffer(29298) := X"8FC20058";
        ram_buffer(29299) := X"8FC30024";
        ram_buffer(29300) := X"00000000";
        ram_buffer(29301) := X"AC430000";
        ram_buffer(29302) := X"8FC20058";
        ram_buffer(29303) := X"00000000";
        ram_buffer(29304) := X"8C420004";
        ram_buffer(29305) := X"00000000";
        ram_buffer(29306) := X"02028023";
        ram_buffer(29307) := X"8FC20058";
        ram_buffer(29308) := X"00000000";
        ram_buffer(29309) := X"8C420004";
        ram_buffer(29310) := X"00000000";
        ram_buffer(29311) := X"02228821";
        ram_buffer(29312) := X"8FC20058";
        ram_buffer(29313) := X"00000000";
        ram_buffer(29314) := X"AC400004";
        ram_buffer(29315) := X"8FC2001C";
        ram_buffer(29316) := X"00000000";
        ram_buffer(29317) := X"1040000D";
        ram_buffer(29318) := X"00000000";
        ram_buffer(29319) := X"8FC20014";
        ram_buffer(29320) := X"00000000";
        ram_buffer(29321) := X"00501823";
        ram_buffer(29322) := X"8FC20050";
        ram_buffer(29323) := X"00000000";
        ram_buffer(29324) := X"14400002";
        ram_buffer(29325) := X"0062001B";
        ram_buffer(29326) := X"0007000D";
        ram_buffer(29327) := X"00001010";
        ram_buffer(29328) := X"00001012";
        ram_buffer(29329) := X"1000004E";
        ram_buffer(29330) := X"00000000";
        ram_buffer(29331) := X"1600FFB7";
        ram_buffer(29332) := X"00000000";
        ram_buffer(29333) := X"10000049";
        ram_buffer(29334) := X"00000000";
        ram_buffer(29335) := X"8FC20058";
        ram_buffer(29336) := X"00000000";
        ram_buffer(29337) := X"8C420000";
        ram_buffer(29338) := X"02401821";
        ram_buffer(29339) := X"00603021";
        ram_buffer(29340) := X"00402821";
        ram_buffer(29341) := X"02202021";
        ram_buffer(29342) := X"0C027F93";
        ram_buffer(29343) := X"00000000";
        ram_buffer(29344) := X"8FC20058";
        ram_buffer(29345) := X"00000000";
        ram_buffer(29346) := X"8C420000";
        ram_buffer(29347) := X"02401821";
        ram_buffer(29348) := X"00431821";
        ram_buffer(29349) := X"8FC20058";
        ram_buffer(29350) := X"00000000";
        ram_buffer(29351) := X"AC430000";
        ram_buffer(29352) := X"02401021";
        ram_buffer(29353) := X"02228821";
        ram_buffer(29354) := X"02401021";
        ram_buffer(29355) := X"02028023";
        ram_buffer(29356) := X"8FC50058";
        ram_buffer(29357) := X"8FC40048";
        ram_buffer(29358) := X"0C028274";
        ram_buffer(29359) := X"00000000";
        ram_buffer(29360) := X"1040000D";
        ram_buffer(29361) := X"00000000";
        ram_buffer(29362) := X"8FC20014";
        ram_buffer(29363) := X"00000000";
        ram_buffer(29364) := X"00501823";
        ram_buffer(29365) := X"8FC20050";
        ram_buffer(29366) := X"00000000";
        ram_buffer(29367) := X"14400002";
        ram_buffer(29368) := X"0062001B";
        ram_buffer(29369) := X"0007000D";
        ram_buffer(29370) := X"00001010";
        ram_buffer(29371) := X"00001012";
        ram_buffer(29372) := X"10000023";
        ram_buffer(29373) := X"00000000";
        ram_buffer(29374) := X"8FC20058";
        ram_buffer(29375) := X"00000000";
        ram_buffer(29376) := X"8C520004";
        ram_buffer(29377) := X"00000000";
        ram_buffer(29378) := X"02401021";
        ram_buffer(29379) := X"0050102B";
        ram_buffer(29380) := X"1440FFD2";
        ram_buffer(29381) := X"00000000";
        ram_buffer(29382) := X"8FC20058";
        ram_buffer(29383) := X"00000000";
        ram_buffer(29384) := X"8C420000";
        ram_buffer(29385) := X"02003021";
        ram_buffer(29386) := X"00402821";
        ram_buffer(29387) := X"02202021";
        ram_buffer(29388) := X"0C027F93";
        ram_buffer(29389) := X"00000000";
        ram_buffer(29390) := X"8FC20058";
        ram_buffer(29391) := X"00000000";
        ram_buffer(29392) := X"8C420004";
        ram_buffer(29393) := X"00000000";
        ram_buffer(29394) := X"00501023";
        ram_buffer(29395) := X"00401821";
        ram_buffer(29396) := X"8FC20058";
        ram_buffer(29397) := X"00000000";
        ram_buffer(29398) := X"AC430004";
        ram_buffer(29399) := X"8FC20058";
        ram_buffer(29400) := X"00000000";
        ram_buffer(29401) := X"8C420000";
        ram_buffer(29402) := X"00000000";
        ram_buffer(29403) := X"00501821";
        ram_buffer(29404) := X"8FC20058";
        ram_buffer(29405) := X"00000000";
        ram_buffer(29406) := X"AC430000";
        ram_buffer(29407) := X"8FC20054";
        ram_buffer(29408) := X"03C0E821";
        ram_buffer(29409) := X"8FBF0044";
        ram_buffer(29410) := X"8FBE0040";
        ram_buffer(29411) := X"8FB2003C";
        ram_buffer(29412) := X"8FB10038";
        ram_buffer(29413) := X"8FB00034";
        ram_buffer(29414) := X"27BD0048";
        ram_buffer(29415) := X"03E00008";
        ram_buffer(29416) := X"00000000";
        ram_buffer(29417) := X"27BDFFE0";
        ram_buffer(29418) := X"AFBF001C";
        ram_buffer(29419) := X"AFBE0018";
        ram_buffer(29420) := X"03A0F021";
        ram_buffer(29421) := X"AFC40020";
        ram_buffer(29422) := X"AFC50024";
        ram_buffer(29423) := X"AFC60028";
        ram_buffer(29424) := X"AFC7002C";
        ram_buffer(29425) := X"8F838098";
        ram_buffer(29426) := X"8FC2002C";
        ram_buffer(29427) := X"00000000";
        ram_buffer(29428) := X"AFA20010";
        ram_buffer(29429) := X"8FC70028";
        ram_buffer(29430) := X"8FC60024";
        ram_buffer(29431) := X"8FC50020";
        ram_buffer(29432) := X"00602021";
        ram_buffer(29433) := X"0C0271B1";
        ram_buffer(29434) := X"00000000";
        ram_buffer(29435) := X"03C0E821";
        ram_buffer(29436) := X"8FBF001C";
        ram_buffer(29437) := X"8FBE0018";
        ram_buffer(29438) := X"27BD0020";
        ram_buffer(29439) := X"03E00008";
        ram_buffer(29440) := X"00000000";
        ram_buffer(29441) := X"27BDFFC0";
        ram_buffer(29442) := X"AFBF003C";
        ram_buffer(29443) := X"AFBE0038";
        ram_buffer(29444) := X"03A0F021";
        ram_buffer(29445) := X"AFC40040";
        ram_buffer(29446) := X"AFC50044";
        ram_buffer(29447) := X"8FC20044";
        ram_buffer(29448) := X"00000000";
        ram_buffer(29449) := X"104001D3";
        ram_buffer(29450) := X"00000000";
        ram_buffer(29451) := X"8FC40040";
        ram_buffer(29452) := X"0C0280C3";
        ram_buffer(29453) := X"00000000";
        ram_buffer(29454) := X"8FC20044";
        ram_buffer(29455) := X"00000000";
        ram_buffer(29456) := X"2442FFF8";
        ram_buffer(29457) := X"AFC20010";
        ram_buffer(29458) := X"8FC20010";
        ram_buffer(29459) := X"00000000";
        ram_buffer(29460) := X"8C420004";
        ram_buffer(29461) := X"00000000";
        ram_buffer(29462) := X"AFC20024";
        ram_buffer(29463) := X"8FC30024";
        ram_buffer(29464) := X"2402FFFE";
        ram_buffer(29465) := X"00621024";
        ram_buffer(29466) := X"AFC20014";
        ram_buffer(29467) := X"8FC30010";
        ram_buffer(29468) := X"8FC20014";
        ram_buffer(29469) := X"00000000";
        ram_buffer(29470) := X"00621021";
        ram_buffer(29471) := X"AFC20028";
        ram_buffer(29472) := X"8FC20028";
        ram_buffer(29473) := X"00000000";
        ram_buffer(29474) := X"8C430004";
        ram_buffer(29475) := X"2402FFFC";
        ram_buffer(29476) := X"00621024";
        ram_buffer(29477) := X"AFC2002C";
        ram_buffer(29478) := X"3C02100D";
        ram_buffer(29479) := X"2442CBE0";
        ram_buffer(29480) := X"8C430008";
        ram_buffer(29481) := X"8FC20028";
        ram_buffer(29482) := X"00000000";
        ram_buffer(29483) := X"1462004A";
        ram_buffer(29484) := X"00000000";
        ram_buffer(29485) := X"8FC30014";
        ram_buffer(29486) := X"8FC2002C";
        ram_buffer(29487) := X"00000000";
        ram_buffer(29488) := X"00621021";
        ram_buffer(29489) := X"AFC20014";
        ram_buffer(29490) := X"8FC20024";
        ram_buffer(29491) := X"00000000";
        ram_buffer(29492) := X"30420001";
        ram_buffer(29493) := X"14400024";
        ram_buffer(29494) := X"00000000";
        ram_buffer(29495) := X"8FC20010";
        ram_buffer(29496) := X"00000000";
        ram_buffer(29497) := X"8C420000";
        ram_buffer(29498) := X"00000000";
        ram_buffer(29499) := X"AFC20030";
        ram_buffer(29500) := X"8FC20030";
        ram_buffer(29501) := X"00000000";
        ram_buffer(29502) := X"00021023";
        ram_buffer(29503) := X"8FC30010";
        ram_buffer(29504) := X"00000000";
        ram_buffer(29505) := X"00621021";
        ram_buffer(29506) := X"AFC20010";
        ram_buffer(29507) := X"8FC30014";
        ram_buffer(29508) := X"8FC20030";
        ram_buffer(29509) := X"00000000";
        ram_buffer(29510) := X"00621021";
        ram_buffer(29511) := X"AFC20014";
        ram_buffer(29512) := X"8FC20010";
        ram_buffer(29513) := X"00000000";
        ram_buffer(29514) := X"8C42000C";
        ram_buffer(29515) := X"00000000";
        ram_buffer(29516) := X"AFC20018";
        ram_buffer(29517) := X"8FC20010";
        ram_buffer(29518) := X"00000000";
        ram_buffer(29519) := X"8C420008";
        ram_buffer(29520) := X"00000000";
        ram_buffer(29521) := X"AFC2001C";
        ram_buffer(29522) := X"8FC2001C";
        ram_buffer(29523) := X"8FC30018";
        ram_buffer(29524) := X"00000000";
        ram_buffer(29525) := X"AC43000C";
        ram_buffer(29526) := X"8FC20018";
        ram_buffer(29527) := X"8FC3001C";
        ram_buffer(29528) := X"00000000";
        ram_buffer(29529) := X"AC430008";
        ram_buffer(29530) := X"8FC20014";
        ram_buffer(29531) := X"00000000";
        ram_buffer(29532) := X"34430001";
        ram_buffer(29533) := X"8FC20010";
        ram_buffer(29534) := X"00000000";
        ram_buffer(29535) := X"AC430004";
        ram_buffer(29536) := X"3C02100D";
        ram_buffer(29537) := X"2442CBE0";
        ram_buffer(29538) := X"8FC30010";
        ram_buffer(29539) := X"00000000";
        ram_buffer(29540) := X"AC430008";
        ram_buffer(29541) := X"8F8280A0";
        ram_buffer(29542) := X"8FC30014";
        ram_buffer(29543) := X"00000000";
        ram_buffer(29544) := X"0062102B";
        ram_buffer(29545) := X"14400007";
        ram_buffer(29546) := X"00000000";
        ram_buffer(29547) := X"8F8281B4";
        ram_buffer(29548) := X"00000000";
        ram_buffer(29549) := X"00402821";
        ram_buffer(29550) := X"8FC40040";
        ram_buffer(29551) := X"0C0274E4";
        ram_buffer(29552) := X"00000000";
        ram_buffer(29553) := X"8FC40040";
        ram_buffer(29554) := X"0C0280CD";
        ram_buffer(29555) := X"00000000";
        ram_buffer(29556) := X"10000169";
        ram_buffer(29557) := X"00000000";
        ram_buffer(29558) := X"8FC20028";
        ram_buffer(29559) := X"8FC3002C";
        ram_buffer(29560) := X"00000000";
        ram_buffer(29561) := X"AC430004";
        ram_buffer(29562) := X"AFC00020";
        ram_buffer(29563) := X"8FC20024";
        ram_buffer(29564) := X"00000000";
        ram_buffer(29565) := X"30420001";
        ram_buffer(29566) := X"1440002F";
        ram_buffer(29567) := X"00000000";
        ram_buffer(29568) := X"8FC20010";
        ram_buffer(29569) := X"00000000";
        ram_buffer(29570) := X"8C420000";
        ram_buffer(29571) := X"00000000";
        ram_buffer(29572) := X"AFC20030";
        ram_buffer(29573) := X"8FC20030";
        ram_buffer(29574) := X"00000000";
        ram_buffer(29575) := X"00021023";
        ram_buffer(29576) := X"8FC30010";
        ram_buffer(29577) := X"00000000";
        ram_buffer(29578) := X"00621021";
        ram_buffer(29579) := X"AFC20010";
        ram_buffer(29580) := X"8FC30014";
        ram_buffer(29581) := X"8FC20030";
        ram_buffer(29582) := X"00000000";
        ram_buffer(29583) := X"00621021";
        ram_buffer(29584) := X"AFC20014";
        ram_buffer(29585) := X"8FC20010";
        ram_buffer(29586) := X"00000000";
        ram_buffer(29587) := X"8C430008";
        ram_buffer(29588) := X"3C02100D";
        ram_buffer(29589) := X"2442CBE8";
        ram_buffer(29590) := X"14620005";
        ram_buffer(29591) := X"00000000";
        ram_buffer(29592) := X"24020001";
        ram_buffer(29593) := X"AFC20020";
        ram_buffer(29594) := X"10000013";
        ram_buffer(29595) := X"00000000";
        ram_buffer(29596) := X"8FC20010";
        ram_buffer(29597) := X"00000000";
        ram_buffer(29598) := X"8C42000C";
        ram_buffer(29599) := X"00000000";
        ram_buffer(29600) := X"AFC20018";
        ram_buffer(29601) := X"8FC20010";
        ram_buffer(29602) := X"00000000";
        ram_buffer(29603) := X"8C420008";
        ram_buffer(29604) := X"00000000";
        ram_buffer(29605) := X"AFC2001C";
        ram_buffer(29606) := X"8FC2001C";
        ram_buffer(29607) := X"8FC30018";
        ram_buffer(29608) := X"00000000";
        ram_buffer(29609) := X"AC43000C";
        ram_buffer(29610) := X"8FC20018";
        ram_buffer(29611) := X"8FC3001C";
        ram_buffer(29612) := X"00000000";
        ram_buffer(29613) := X"AC430008";
        ram_buffer(29614) := X"8FC30028";
        ram_buffer(29615) := X"8FC2002C";
        ram_buffer(29616) := X"00000000";
        ram_buffer(29617) := X"00621021";
        ram_buffer(29618) := X"8C420004";
        ram_buffer(29619) := X"00000000";
        ram_buffer(29620) := X"30420001";
        ram_buffer(29621) := X"1440003C";
        ram_buffer(29622) := X"00000000";
        ram_buffer(29623) := X"8FC30014";
        ram_buffer(29624) := X"8FC2002C";
        ram_buffer(29625) := X"00000000";
        ram_buffer(29626) := X"00621021";
        ram_buffer(29627) := X"AFC20014";
        ram_buffer(29628) := X"8FC20020";
        ram_buffer(29629) := X"00000000";
        ram_buffer(29630) := X"14400021";
        ram_buffer(29631) := X"00000000";
        ram_buffer(29632) := X"8FC20028";
        ram_buffer(29633) := X"00000000";
        ram_buffer(29634) := X"8C430008";
        ram_buffer(29635) := X"3C02100D";
        ram_buffer(29636) := X"2442CBE8";
        ram_buffer(29637) := X"1462001A";
        ram_buffer(29638) := X"00000000";
        ram_buffer(29639) := X"24020001";
        ram_buffer(29640) := X"AFC20020";
        ram_buffer(29641) := X"3C02100D";
        ram_buffer(29642) := X"2443CBE8";
        ram_buffer(29643) := X"3C02100D";
        ram_buffer(29644) := X"2442CBE8";
        ram_buffer(29645) := X"8FC40010";
        ram_buffer(29646) := X"00000000";
        ram_buffer(29647) := X"AC44000C";
        ram_buffer(29648) := X"8C42000C";
        ram_buffer(29649) := X"00000000";
        ram_buffer(29650) := X"AC620008";
        ram_buffer(29651) := X"3C02100D";
        ram_buffer(29652) := X"2443CBE8";
        ram_buffer(29653) := X"8FC20010";
        ram_buffer(29654) := X"00000000";
        ram_buffer(29655) := X"AC43000C";
        ram_buffer(29656) := X"8FC20010";
        ram_buffer(29657) := X"00000000";
        ram_buffer(29658) := X"8C43000C";
        ram_buffer(29659) := X"8FC20010";
        ram_buffer(29660) := X"00000000";
        ram_buffer(29661) := X"AC430008";
        ram_buffer(29662) := X"10000013";
        ram_buffer(29663) := X"00000000";
        ram_buffer(29664) := X"8FC20028";
        ram_buffer(29665) := X"00000000";
        ram_buffer(29666) := X"8C42000C";
        ram_buffer(29667) := X"00000000";
        ram_buffer(29668) := X"AFC20018";
        ram_buffer(29669) := X"8FC20028";
        ram_buffer(29670) := X"00000000";
        ram_buffer(29671) := X"8C420008";
        ram_buffer(29672) := X"00000000";
        ram_buffer(29673) := X"AFC2001C";
        ram_buffer(29674) := X"8FC2001C";
        ram_buffer(29675) := X"8FC30018";
        ram_buffer(29676) := X"00000000";
        ram_buffer(29677) := X"AC43000C";
        ram_buffer(29678) := X"8FC20018";
        ram_buffer(29679) := X"8FC3001C";
        ram_buffer(29680) := X"00000000";
        ram_buffer(29681) := X"AC430008";
        ram_buffer(29682) := X"8FC20014";
        ram_buffer(29683) := X"00000000";
        ram_buffer(29684) := X"34430001";
        ram_buffer(29685) := X"8FC20010";
        ram_buffer(29686) := X"00000000";
        ram_buffer(29687) := X"AC430004";
        ram_buffer(29688) := X"8FC30010";
        ram_buffer(29689) := X"8FC20014";
        ram_buffer(29690) := X"00000000";
        ram_buffer(29691) := X"00621021";
        ram_buffer(29692) := X"8FC30014";
        ram_buffer(29693) := X"00000000";
        ram_buffer(29694) := X"AC430000";
        ram_buffer(29695) := X"8FC20020";
        ram_buffer(29696) := X"00000000";
        ram_buffer(29697) := X"144000D6";
        ram_buffer(29698) := X"00000000";
        ram_buffer(29699) := X"8FC20014";
        ram_buffer(29700) := X"00000000";
        ram_buffer(29701) := X"2C420200";
        ram_buffer(29702) := X"10400038";
        ram_buffer(29703) := X"00000000";
        ram_buffer(29704) := X"8FC20014";
        ram_buffer(29705) := X"00000000";
        ram_buffer(29706) := X"000210C2";
        ram_buffer(29707) := X"AFC20034";
        ram_buffer(29708) := X"3C02100D";
        ram_buffer(29709) := X"2443CBE0";
        ram_buffer(29710) := X"3C02100D";
        ram_buffer(29711) := X"2442CBE0";
        ram_buffer(29712) := X"8C440004";
        ram_buffer(29713) := X"8FC20034";
        ram_buffer(29714) := X"00000000";
        ram_buffer(29715) := X"04410002";
        ram_buffer(29716) := X"00000000";
        ram_buffer(29717) := X"24420003";
        ram_buffer(29718) := X"00021083";
        ram_buffer(29719) := X"00402821";
        ram_buffer(29720) := X"24020001";
        ram_buffer(29721) := X"00A21004";
        ram_buffer(29722) := X"00821025";
        ram_buffer(29723) := X"AC620004";
        ram_buffer(29724) := X"8FC20034";
        ram_buffer(29725) := X"00000000";
        ram_buffer(29726) := X"24420001";
        ram_buffer(29727) := X"00021040";
        ram_buffer(29728) := X"00021880";
        ram_buffer(29729) := X"3C02100D";
        ram_buffer(29730) := X"2442CBE0";
        ram_buffer(29731) := X"00621021";
        ram_buffer(29732) := X"2442FFF8";
        ram_buffer(29733) := X"AFC20018";
        ram_buffer(29734) := X"8FC20018";
        ram_buffer(29735) := X"00000000";
        ram_buffer(29736) := X"8C420008";
        ram_buffer(29737) := X"00000000";
        ram_buffer(29738) := X"AFC2001C";
        ram_buffer(29739) := X"8FC20010";
        ram_buffer(29740) := X"8FC30018";
        ram_buffer(29741) := X"00000000";
        ram_buffer(29742) := X"AC43000C";
        ram_buffer(29743) := X"8FC20010";
        ram_buffer(29744) := X"8FC3001C";
        ram_buffer(29745) := X"00000000";
        ram_buffer(29746) := X"AC430008";
        ram_buffer(29747) := X"8FC20018";
        ram_buffer(29748) := X"8FC30010";
        ram_buffer(29749) := X"00000000";
        ram_buffer(29750) := X"AC430008";
        ram_buffer(29751) := X"8FC20018";
        ram_buffer(29752) := X"00000000";
        ram_buffer(29753) := X"8C430008";
        ram_buffer(29754) := X"8FC2001C";
        ram_buffer(29755) := X"00000000";
        ram_buffer(29756) := X"AC43000C";
        ram_buffer(29757) := X"1000009A";
        ram_buffer(29758) := X"00000000";
        ram_buffer(29759) := X"8FC20014";
        ram_buffer(29760) := X"00000000";
        ram_buffer(29761) := X"00021242";
        ram_buffer(29762) := X"14400006";
        ram_buffer(29763) := X"00000000";
        ram_buffer(29764) := X"8FC20014";
        ram_buffer(29765) := X"00000000";
        ram_buffer(29766) := X"000210C2";
        ram_buffer(29767) := X"1000003E";
        ram_buffer(29768) := X"00000000";
        ram_buffer(29769) := X"8FC20014";
        ram_buffer(29770) := X"00000000";
        ram_buffer(29771) := X"00021242";
        ram_buffer(29772) := X"2C420005";
        ram_buffer(29773) := X"10400007";
        ram_buffer(29774) := X"00000000";
        ram_buffer(29775) := X"8FC20014";
        ram_buffer(29776) := X"00000000";
        ram_buffer(29777) := X"00021182";
        ram_buffer(29778) := X"24420038";
        ram_buffer(29779) := X"10000032";
        ram_buffer(29780) := X"00000000";
        ram_buffer(29781) := X"8FC20014";
        ram_buffer(29782) := X"00000000";
        ram_buffer(29783) := X"00021242";
        ram_buffer(29784) := X"2C420015";
        ram_buffer(29785) := X"10400007";
        ram_buffer(29786) := X"00000000";
        ram_buffer(29787) := X"8FC20014";
        ram_buffer(29788) := X"00000000";
        ram_buffer(29789) := X"00021242";
        ram_buffer(29790) := X"2442005B";
        ram_buffer(29791) := X"10000026";
        ram_buffer(29792) := X"00000000";
        ram_buffer(29793) := X"8FC20014";
        ram_buffer(29794) := X"00000000";
        ram_buffer(29795) := X"00021242";
        ram_buffer(29796) := X"2C420055";
        ram_buffer(29797) := X"10400007";
        ram_buffer(29798) := X"00000000";
        ram_buffer(29799) := X"8FC20014";
        ram_buffer(29800) := X"00000000";
        ram_buffer(29801) := X"00021302";
        ram_buffer(29802) := X"2442006E";
        ram_buffer(29803) := X"1000001A";
        ram_buffer(29804) := X"00000000";
        ram_buffer(29805) := X"8FC20014";
        ram_buffer(29806) := X"00000000";
        ram_buffer(29807) := X"00021242";
        ram_buffer(29808) := X"2C420155";
        ram_buffer(29809) := X"10400007";
        ram_buffer(29810) := X"00000000";
        ram_buffer(29811) := X"8FC20014";
        ram_buffer(29812) := X"00000000";
        ram_buffer(29813) := X"000213C2";
        ram_buffer(29814) := X"24420077";
        ram_buffer(29815) := X"1000000E";
        ram_buffer(29816) := X"00000000";
        ram_buffer(29817) := X"8FC20014";
        ram_buffer(29818) := X"00000000";
        ram_buffer(29819) := X"00021242";
        ram_buffer(29820) := X"2C420555";
        ram_buffer(29821) := X"10400007";
        ram_buffer(29822) := X"00000000";
        ram_buffer(29823) := X"8FC20014";
        ram_buffer(29824) := X"00000000";
        ram_buffer(29825) := X"00021482";
        ram_buffer(29826) := X"2442007C";
        ram_buffer(29827) := X"10000002";
        ram_buffer(29828) := X"00000000";
        ram_buffer(29829) := X"2402007E";
        ram_buffer(29830) := X"AFC20034";
        ram_buffer(29831) := X"8FC20034";
        ram_buffer(29832) := X"00000000";
        ram_buffer(29833) := X"24420001";
        ram_buffer(29834) := X"00021040";
        ram_buffer(29835) := X"00021880";
        ram_buffer(29836) := X"3C02100D";
        ram_buffer(29837) := X"2442CBE0";
        ram_buffer(29838) := X"00621021";
        ram_buffer(29839) := X"2442FFF8";
        ram_buffer(29840) := X"AFC20018";
        ram_buffer(29841) := X"8FC20018";
        ram_buffer(29842) := X"00000000";
        ram_buffer(29843) := X"8C420008";
        ram_buffer(29844) := X"00000000";
        ram_buffer(29845) := X"AFC2001C";
        ram_buffer(29846) := X"8FC3001C";
        ram_buffer(29847) := X"8FC20018";
        ram_buffer(29848) := X"00000000";
        ram_buffer(29849) := X"14620018";
        ram_buffer(29850) := X"00000000";
        ram_buffer(29851) := X"3C02100D";
        ram_buffer(29852) := X"2443CBE0";
        ram_buffer(29853) := X"3C02100D";
        ram_buffer(29854) := X"2442CBE0";
        ram_buffer(29855) := X"8C440004";
        ram_buffer(29856) := X"8FC20034";
        ram_buffer(29857) := X"00000000";
        ram_buffer(29858) := X"04410002";
        ram_buffer(29859) := X"00000000";
        ram_buffer(29860) := X"24420003";
        ram_buffer(29861) := X"00021083";
        ram_buffer(29862) := X"00402821";
        ram_buffer(29863) := X"24020001";
        ram_buffer(29864) := X"00A21004";
        ram_buffer(29865) := X"00821025";
        ram_buffer(29866) := X"AC620004";
        ram_buffer(29867) := X"1000001A";
        ram_buffer(29868) := X"00000000";
        ram_buffer(29869) := X"8FC2001C";
        ram_buffer(29870) := X"00000000";
        ram_buffer(29871) := X"8C420008";
        ram_buffer(29872) := X"00000000";
        ram_buffer(29873) := X"AFC2001C";
        ram_buffer(29874) := X"8FC3001C";
        ram_buffer(29875) := X"8FC20018";
        ram_buffer(29876) := X"00000000";
        ram_buffer(29877) := X"1062000B";
        ram_buffer(29878) := X"00000000";
        ram_buffer(29879) := X"8FC2001C";
        ram_buffer(29880) := X"00000000";
        ram_buffer(29881) := X"8C430004";
        ram_buffer(29882) := X"2402FFFC";
        ram_buffer(29883) := X"00621824";
        ram_buffer(29884) := X"8FC20014";
        ram_buffer(29885) := X"00000000";
        ram_buffer(29886) := X"0043102B";
        ram_buffer(29887) := X"1440FFED";
        ram_buffer(29888) := X"00000000";
        ram_buffer(29889) := X"8FC2001C";
        ram_buffer(29890) := X"00000000";
        ram_buffer(29891) := X"8C42000C";
        ram_buffer(29892) := X"00000000";
        ram_buffer(29893) := X"AFC20018";
        ram_buffer(29894) := X"8FC20010";
        ram_buffer(29895) := X"8FC30018";
        ram_buffer(29896) := X"00000000";
        ram_buffer(29897) := X"AC43000C";
        ram_buffer(29898) := X"8FC20010";
        ram_buffer(29899) := X"8FC3001C";
        ram_buffer(29900) := X"00000000";
        ram_buffer(29901) := X"AC430008";
        ram_buffer(29902) := X"8FC20018";
        ram_buffer(29903) := X"8FC30010";
        ram_buffer(29904) := X"00000000";
        ram_buffer(29905) := X"AC430008";
        ram_buffer(29906) := X"8FC20018";
        ram_buffer(29907) := X"00000000";
        ram_buffer(29908) := X"8C430008";
        ram_buffer(29909) := X"8FC2001C";
        ram_buffer(29910) := X"00000000";
        ram_buffer(29911) := X"AC43000C";
        ram_buffer(29912) := X"8FC40040";
        ram_buffer(29913) := X"0C0280CD";
        ram_buffer(29914) := X"00000000";
        ram_buffer(29915) := X"10000002";
        ram_buffer(29916) := X"00000000";
        ram_buffer(29917) := X"00000000";
        ram_buffer(29918) := X"03C0E821";
        ram_buffer(29919) := X"8FBF003C";
        ram_buffer(29920) := X"8FBE0038";
        ram_buffer(29921) := X"27BD0040";
        ram_buffer(29922) := X"03E00008";
        ram_buffer(29923) := X"00000000";
        ram_buffer(29924) := X"27BDFFD0";
        ram_buffer(29925) := X"AFBF002C";
        ram_buffer(29926) := X"AFBE0028";
        ram_buffer(29927) := X"03A0F021";
        ram_buffer(29928) := X"AFC40030";
        ram_buffer(29929) := X"AFC50034";
        ram_buffer(29930) := X"24021000";
        ram_buffer(29931) := X"AFC20010";
        ram_buffer(29932) := X"8FC40030";
        ram_buffer(29933) := X"0C0280C3";
        ram_buffer(29934) := X"00000000";
        ram_buffer(29935) := X"3C02100D";
        ram_buffer(29936) := X"2442CBE0";
        ram_buffer(29937) := X"8C420008";
        ram_buffer(29938) := X"00000000";
        ram_buffer(29939) := X"8C420004";
        ram_buffer(29940) := X"00000000";
        ram_buffer(29941) := X"00401821";
        ram_buffer(29942) := X"2402FFFC";
        ram_buffer(29943) := X"00621024";
        ram_buffer(29944) := X"AFC20014";
        ram_buffer(29945) := X"8FC30014";
        ram_buffer(29946) := X"8FC20034";
        ram_buffer(29947) := X"00000000";
        ram_buffer(29948) := X"00621823";
        ram_buffer(29949) := X"8FC20010";
        ram_buffer(29950) := X"00000000";
        ram_buffer(29951) := X"00621021";
        ram_buffer(29952) := X"2443FFEF";
        ram_buffer(29953) := X"8FC20010";
        ram_buffer(29954) := X"00000000";
        ram_buffer(29955) := X"14400002";
        ram_buffer(29956) := X"0062001B";
        ram_buffer(29957) := X"0007000D";
        ram_buffer(29958) := X"00001010";
        ram_buffer(29959) := X"00001012";
        ram_buffer(29960) := X"2443FFFF";
        ram_buffer(29961) := X"8FC20010";
        ram_buffer(29962) := X"00000000";
        ram_buffer(29963) := X"00620018";
        ram_buffer(29964) := X"00001012";
        ram_buffer(29965) := X"AFC20018";
        ram_buffer(29966) := X"8FC20010";
        ram_buffer(29967) := X"8FC30018";
        ram_buffer(29968) := X"00000000";
        ram_buffer(29969) := X"0062102A";
        ram_buffer(29970) := X"10400007";
        ram_buffer(29971) := X"00000000";
        ram_buffer(29972) := X"8FC40030";
        ram_buffer(29973) := X"0C0280CD";
        ram_buffer(29974) := X"00000000";
        ram_buffer(29975) := X"00001021";
        ram_buffer(29976) := X"1000005A";
        ram_buffer(29977) := X"00000000";
        ram_buffer(29978) := X"00002821";
        ram_buffer(29979) := X"8FC40030";
        ram_buffer(29980) := X"0C028390";
        ram_buffer(29981) := X"00000000";
        ram_buffer(29982) := X"AFC2001C";
        ram_buffer(29983) := X"3C02100D";
        ram_buffer(29984) := X"2442CBE0";
        ram_buffer(29985) := X"8C430008";
        ram_buffer(29986) := X"8FC20014";
        ram_buffer(29987) := X"00000000";
        ram_buffer(29988) := X"00621821";
        ram_buffer(29989) := X"8FC2001C";
        ram_buffer(29990) := X"00000000";
        ram_buffer(29991) := X"10620007";
        ram_buffer(29992) := X"00000000";
        ram_buffer(29993) := X"8FC40030";
        ram_buffer(29994) := X"0C0280CD";
        ram_buffer(29995) := X"00000000";
        ram_buffer(29996) := X"00001021";
        ram_buffer(29997) := X"10000045";
        ram_buffer(29998) := X"00000000";
        ram_buffer(29999) := X"8FC20018";
        ram_buffer(30000) := X"00000000";
        ram_buffer(30001) := X"00021023";
        ram_buffer(30002) := X"00402821";
        ram_buffer(30003) := X"8FC40030";
        ram_buffer(30004) := X"0C028390";
        ram_buffer(30005) := X"00000000";
        ram_buffer(30006) := X"AFC20020";
        ram_buffer(30007) := X"8FC30020";
        ram_buffer(30008) := X"2402FFFF";
        ram_buffer(30009) := X"14620025";
        ram_buffer(30010) := X"00000000";
        ram_buffer(30011) := X"00002821";
        ram_buffer(30012) := X"8FC40030";
        ram_buffer(30013) := X"0C028390";
        ram_buffer(30014) := X"00000000";
        ram_buffer(30015) := X"AFC2001C";
        ram_buffer(30016) := X"8FC2001C";
        ram_buffer(30017) := X"3C03100D";
        ram_buffer(30018) := X"2463CBE0";
        ram_buffer(30019) := X"8C630008";
        ram_buffer(30020) := X"00000000";
        ram_buffer(30021) := X"00431023";
        ram_buffer(30022) := X"AFC20014";
        ram_buffer(30023) := X"8FC20014";
        ram_buffer(30024) := X"00000000";
        ram_buffer(30025) := X"28420010";
        ram_buffer(30026) := X"1440000E";
        ram_buffer(30027) := X"00000000";
        ram_buffer(30028) := X"8FC2001C";
        ram_buffer(30029) := X"8F8380A4";
        ram_buffer(30030) := X"00000000";
        ram_buffer(30031) := X"00431823";
        ram_buffer(30032) := X"3C02100D";
        ram_buffer(30033) := X"AC43D260";
        ram_buffer(30034) := X"3C02100D";
        ram_buffer(30035) := X"2442CBE0";
        ram_buffer(30036) := X"8C420008";
        ram_buffer(30037) := X"8FC30014";
        ram_buffer(30038) := X"00000000";
        ram_buffer(30039) := X"34630001";
        ram_buffer(30040) := X"AC430004";
        ram_buffer(30041) := X"8FC40030";
        ram_buffer(30042) := X"0C0280CD";
        ram_buffer(30043) := X"00000000";
        ram_buffer(30044) := X"00001021";
        ram_buffer(30045) := X"10000015";
        ram_buffer(30046) := X"00000000";
        ram_buffer(30047) := X"3C02100D";
        ram_buffer(30048) := X"2442CBE0";
        ram_buffer(30049) := X"8C420008";
        ram_buffer(30050) := X"8FC40014";
        ram_buffer(30051) := X"8FC30018";
        ram_buffer(30052) := X"00000000";
        ram_buffer(30053) := X"00831823";
        ram_buffer(30054) := X"34630001";
        ram_buffer(30055) := X"AC430004";
        ram_buffer(30056) := X"3C02100D";
        ram_buffer(30057) := X"8C43D260";
        ram_buffer(30058) := X"8FC20018";
        ram_buffer(30059) := X"00000000";
        ram_buffer(30060) := X"00621823";
        ram_buffer(30061) := X"3C02100D";
        ram_buffer(30062) := X"AC43D260";
        ram_buffer(30063) := X"8FC40030";
        ram_buffer(30064) := X"0C0280CD";
        ram_buffer(30065) := X"00000000";
        ram_buffer(30066) := X"24020001";
        ram_buffer(30067) := X"03C0E821";
        ram_buffer(30068) := X"8FBF002C";
        ram_buffer(30069) := X"8FBE0028";
        ram_buffer(30070) := X"27BD0030";
        ram_buffer(30071) := X"03E00008";
        ram_buffer(30072) := X"00000000";
        ram_buffer(30073) := X"27BDFFE8";
        ram_buffer(30074) := X"AFBF0014";
        ram_buffer(30075) := X"AFBE0010";
        ram_buffer(30076) := X"03A0F021";
        ram_buffer(30077) := X"AFC40018";
        ram_buffer(30078) := X"00A01021";
        ram_buffer(30079) := X"AFC60020";
        ram_buffer(30080) := X"AFC70024";
        ram_buffer(30081) := X"8FC70024";
        ram_buffer(30082) := X"8FC60020";
        ram_buffer(30083) := X"00402821";
        ram_buffer(30084) := X"8FC40018";
        ram_buffer(30085) := X"0C0275A1";
        ram_buffer(30086) := X"00000000";
        ram_buffer(30087) := X"03C0E821";
        ram_buffer(30088) := X"8FBF0014";
        ram_buffer(30089) := X"8FBE0010";
        ram_buffer(30090) := X"27BD0018";
        ram_buffer(30091) := X"03E00008";
        ram_buffer(30092) := X"00000000";
        ram_buffer(30093) := X"27BDFFE8";
        ram_buffer(30094) := X"AFBF0014";
        ram_buffer(30095) := X"AFBE0010";
        ram_buffer(30096) := X"03A0F021";
        ram_buffer(30097) := X"00801821";
        ram_buffer(30098) := X"AFC5001C";
        ram_buffer(30099) := X"AFC60020";
        ram_buffer(30100) := X"8F828098";
        ram_buffer(30101) := X"8FC70020";
        ram_buffer(30102) := X"8FC6001C";
        ram_buffer(30103) := X"00602821";
        ram_buffer(30104) := X"00402021";
        ram_buffer(30105) := X"0C027579";
        ram_buffer(30106) := X"00000000";
        ram_buffer(30107) := X"03C0E821";
        ram_buffer(30108) := X"8FBF0014";
        ram_buffer(30109) := X"8FBE0010";
        ram_buffer(30110) := X"27BD0018";
        ram_buffer(30111) := X"03E00008";
        ram_buffer(30112) := X"00000000";
        ram_buffer(30113) := X"27BDFF88";
        ram_buffer(30114) := X"AFBF0074";
        ram_buffer(30115) := X"AFBE0070";
        ram_buffer(30116) := X"AFB0006C";
        ram_buffer(30117) := X"03A0F021";
        ram_buffer(30118) := X"AFC40078";
        ram_buffer(30119) := X"00A08021";
        ram_buffer(30120) := X"AFC60080";
        ram_buffer(30121) := X"AFC70084";
        ram_buffer(30122) := X"AFC00014";
        ram_buffer(30123) := X"8FC20078";
        ram_buffer(30124) := X"00000000";
        ram_buffer(30125) := X"AFC20020";
        ram_buffer(30126) := X"8FC20020";
        ram_buffer(30127) := X"00000000";
        ram_buffer(30128) := X"1040000A";
        ram_buffer(30129) := X"00000000";
        ram_buffer(30130) := X"8FC20020";
        ram_buffer(30131) := X"00000000";
        ram_buffer(30132) := X"8C420038";
        ram_buffer(30133) := X"00000000";
        ram_buffer(30134) := X"14400004";
        ram_buffer(30135) := X"00000000";
        ram_buffer(30136) := X"8FC40020";
        ram_buffer(30137) := X"0C027069";
        ram_buffer(30138) := X"00000000";
        ram_buffer(30139) := X"8602000C";
        ram_buffer(30140) := X"00000000";
        ram_buffer(30141) := X"3042FFFF";
        ram_buffer(30142) := X"30420100";
        ram_buffer(30143) := X"1040000B";
        ram_buffer(30144) := X"00000000";
        ram_buffer(30145) := X"8602000C";
        ram_buffer(30146) := X"00000000";
        ram_buffer(30147) := X"3042FFFF";
        ram_buffer(30148) := X"30420008";
        ram_buffer(30149) := X"10400005";
        ram_buffer(30150) := X"00000000";
        ram_buffer(30151) := X"02002821";
        ram_buffer(30152) := X"8FC40078";
        ram_buffer(30153) := X"0C026EE1";
        ram_buffer(30154) := X"00000000";
        ram_buffer(30155) := X"8E020028";
        ram_buffer(30156) := X"00000000";
        ram_buffer(30157) := X"AFC20024";
        ram_buffer(30158) := X"8FC20024";
        ram_buffer(30159) := X"00000000";
        ram_buffer(30160) := X"14400007";
        ram_buffer(30161) := X"00000000";
        ram_buffer(30162) := X"8FC20078";
        ram_buffer(30163) := X"2403001D";
        ram_buffer(30164) := X"AC430000";
        ram_buffer(30165) := X"2402FFFF";
        ram_buffer(30166) := X"100001F1";
        ram_buffer(30167) := X"00000000";
        ram_buffer(30168) := X"8FC20084";
        ram_buffer(30169) := X"24030001";
        ram_buffer(30170) := X"10430008";
        ram_buffer(30171) := X"00000000";
        ram_buffer(30172) := X"24030002";
        ram_buffer(30173) := X"10430058";
        ram_buffer(30174) := X"00000000";
        ram_buffer(30175) := X"10400056";
        ram_buffer(30176) := X"00000000";
        ram_buffer(30177) := X"10000057";
        ram_buffer(30178) := X"00000000";
        ram_buffer(30179) := X"02002821";
        ram_buffer(30180) := X"8FC40078";
        ram_buffer(30181) := X"0C026EE1";
        ram_buffer(30182) := X"00000000";
        ram_buffer(30183) := X"8602000C";
        ram_buffer(30184) := X"00000000";
        ram_buffer(30185) := X"3042FFFF";
        ram_buffer(30186) := X"30421000";
        ram_buffer(30187) := X"10400006";
        ram_buffer(30188) := X"00000000";
        ram_buffer(30189) := X"8E020050";
        ram_buffer(30190) := X"00000000";
        ram_buffer(30191) := X"AFC20014";
        ram_buffer(30192) := X"10000011";
        ram_buffer(30193) := X"00000000";
        ram_buffer(30194) := X"8E03001C";
        ram_buffer(30195) := X"8FC20024";
        ram_buffer(30196) := X"24070001";
        ram_buffer(30197) := X"00003021";
        ram_buffer(30198) := X"00602821";
        ram_buffer(30199) := X"8FC40078";
        ram_buffer(30200) := X"0040F809";
        ram_buffer(30201) := X"00000000";
        ram_buffer(30202) := X"AFC20014";
        ram_buffer(30203) := X"8FC30014";
        ram_buffer(30204) := X"2402FFFF";
        ram_buffer(30205) := X"14620004";
        ram_buffer(30206) := X"00000000";
        ram_buffer(30207) := X"2402FFFF";
        ram_buffer(30208) := X"100001C7";
        ram_buffer(30209) := X"00000000";
        ram_buffer(30210) := X"8602000C";
        ram_buffer(30211) := X"00000000";
        ram_buffer(30212) := X"3042FFFF";
        ram_buffer(30213) := X"30420004";
        ram_buffer(30214) := X"10400011";
        ram_buffer(30215) := X"00000000";
        ram_buffer(30216) := X"8E020004";
        ram_buffer(30217) := X"8FC30014";
        ram_buffer(30218) := X"00000000";
        ram_buffer(30219) := X"00621023";
        ram_buffer(30220) := X"AFC20014";
        ram_buffer(30221) := X"8E020030";
        ram_buffer(30222) := X"00000000";
        ram_buffer(30223) := X"1040001C";
        ram_buffer(30224) := X"00000000";
        ram_buffer(30225) := X"8E02003C";
        ram_buffer(30226) := X"8FC30014";
        ram_buffer(30227) := X"00000000";
        ram_buffer(30228) := X"00621023";
        ram_buffer(30229) := X"AFC20014";
        ram_buffer(30230) := X"10000015";
        ram_buffer(30231) := X"00000000";
        ram_buffer(30232) := X"8602000C";
        ram_buffer(30233) := X"00000000";
        ram_buffer(30234) := X"3042FFFF";
        ram_buffer(30235) := X"30420008";
        ram_buffer(30236) := X"1040000F";
        ram_buffer(30237) := X"00000000";
        ram_buffer(30238) := X"8E020000";
        ram_buffer(30239) := X"00000000";
        ram_buffer(30240) := X"1040000B";
        ram_buffer(30241) := X"00000000";
        ram_buffer(30242) := X"8E020000";
        ram_buffer(30243) := X"00000000";
        ram_buffer(30244) := X"00401821";
        ram_buffer(30245) := X"8E020010";
        ram_buffer(30246) := X"00000000";
        ram_buffer(30247) := X"00621023";
        ram_buffer(30248) := X"8FC30014";
        ram_buffer(30249) := X"00000000";
        ram_buffer(30250) := X"00621021";
        ram_buffer(30251) := X"AFC20014";
        ram_buffer(30252) := X"8FC30080";
        ram_buffer(30253) := X"8FC20014";
        ram_buffer(30254) := X"00000000";
        ram_buffer(30255) := X"00621021";
        ram_buffer(30256) := X"AFC20080";
        ram_buffer(30257) := X"AFC00084";
        ram_buffer(30258) := X"24020001";
        ram_buffer(30259) := X"AFC2001C";
        ram_buffer(30260) := X"1000000A";
        ram_buffer(30261) := X"00000000";
        ram_buffer(30262) := X"AFC0001C";
        ram_buffer(30263) := X"10000007";
        ram_buffer(30264) := X"00000000";
        ram_buffer(30265) := X"8FC20078";
        ram_buffer(30266) := X"24030016";
        ram_buffer(30267) := X"AC430000";
        ram_buffer(30268) := X"2402FFFF";
        ram_buffer(30269) := X"1000018A";
        ram_buffer(30270) := X"00000000";
        ram_buffer(30271) := X"8E020010";
        ram_buffer(30272) := X"00000000";
        ram_buffer(30273) := X"14400005";
        ram_buffer(30274) := X"00000000";
        ram_buffer(30275) := X"02002821";
        ram_buffer(30276) := X"8FC40078";
        ram_buffer(30277) := X"0C027999";
        ram_buffer(30278) := X"00000000";
        ram_buffer(30279) := X"8602000C";
        ram_buffer(30280) := X"00000000";
        ram_buffer(30281) := X"3042FFFF";
        ram_buffer(30282) := X"3042081A";
        ram_buffer(30283) := X"14400137";
        ram_buffer(30284) := X"00000000";
        ram_buffer(30285) := X"8602000C";
        ram_buffer(30286) := X"00000000";
        ram_buffer(30287) := X"3042FFFF";
        ram_buffer(30288) := X"30420400";
        ram_buffer(30289) := X"1440002B";
        ram_buffer(30290) := X"00000000";
        ram_buffer(30291) := X"8FC30024";
        ram_buffer(30292) := X"3C02100A";
        ram_buffer(30293) := X"24421360";
        ram_buffer(30294) := X"14620016";
        ram_buffer(30295) := X"00000000";
        ram_buffer(30296) := X"8602000E";
        ram_buffer(30297) := X"00000000";
        ram_buffer(30298) := X"04400012";
        ram_buffer(30299) := X"00000000";
        ram_buffer(30300) := X"8602000E";
        ram_buffer(30301) := X"00000000";
        ram_buffer(30302) := X"00401821";
        ram_buffer(30303) := X"27C20028";
        ram_buffer(30304) := X"00403021";
        ram_buffer(30305) := X"00602821";
        ram_buffer(30306) := X"8FC40078";
        ram_buffer(30307) := X"0C0277E3";
        ram_buffer(30308) := X"00000000";
        ram_buffer(30309) := X"14400007";
        ram_buffer(30310) := X"00000000";
        ram_buffer(30311) := X"8FC2002C";
        ram_buffer(30312) := X"00000000";
        ram_buffer(30313) := X"3043F000";
        ram_buffer(30314) := X"34028000";
        ram_buffer(30315) := X"10620009";
        ram_buffer(30316) := X"00000000";
        ram_buffer(30317) := X"8602000C";
        ram_buffer(30318) := X"00000000";
        ram_buffer(30319) := X"34420800";
        ram_buffer(30320) := X"00021400";
        ram_buffer(30321) := X"00021403";
        ram_buffer(30322) := X"A602000C";
        ram_buffer(30323) := X"10000119";
        ram_buffer(30324) := X"00000000";
        ram_buffer(30325) := X"24020400";
        ram_buffer(30326) := X"AE02004C";
        ram_buffer(30327) := X"8602000C";
        ram_buffer(30328) := X"00000000";
        ram_buffer(30329) := X"34420400";
        ram_buffer(30330) := X"00021400";
        ram_buffer(30331) := X"00021403";
        ram_buffer(30332) := X"A602000C";
        ram_buffer(30333) := X"8FC20084";
        ram_buffer(30334) := X"00000000";
        ram_buffer(30335) := X"14400006";
        ram_buffer(30336) := X"00000000";
        ram_buffer(30337) := X"8FC20080";
        ram_buffer(30338) := X"00000000";
        ram_buffer(30339) := X"AFC20010";
        ram_buffer(30340) := X"10000011";
        ram_buffer(30341) := X"00000000";
        ram_buffer(30342) := X"8602000E";
        ram_buffer(30343) := X"00000000";
        ram_buffer(30344) := X"00401821";
        ram_buffer(30345) := X"27C20028";
        ram_buffer(30346) := X"00403021";
        ram_buffer(30347) := X"00602821";
        ram_buffer(30348) := X"8FC40078";
        ram_buffer(30349) := X"0C0277E3";
        ram_buffer(30350) := X"00000000";
        ram_buffer(30351) := X"144000F6";
        ram_buffer(30352) := X"00000000";
        ram_buffer(30353) := X"8FC30038";
        ram_buffer(30354) := X"8FC20080";
        ram_buffer(30355) := X"00000000";
        ram_buffer(30356) := X"00621021";
        ram_buffer(30357) := X"AFC20010";
        ram_buffer(30358) := X"8FC2001C";
        ram_buffer(30359) := X"00000000";
        ram_buffer(30360) := X"14400027";
        ram_buffer(30361) := X"00000000";
        ram_buffer(30362) := X"8602000C";
        ram_buffer(30363) := X"00000000";
        ram_buffer(30364) := X"3042FFFF";
        ram_buffer(30365) := X"30421000";
        ram_buffer(30366) := X"10400006";
        ram_buffer(30367) := X"00000000";
        ram_buffer(30368) := X"8E020050";
        ram_buffer(30369) := X"00000000";
        ram_buffer(30370) := X"AFC20014";
        ram_buffer(30371) := X"1000000E";
        ram_buffer(30372) := X"00000000";
        ram_buffer(30373) := X"8E03001C";
        ram_buffer(30374) := X"8FC20024";
        ram_buffer(30375) := X"24070001";
        ram_buffer(30376) := X"00003021";
        ram_buffer(30377) := X"00602821";
        ram_buffer(30378) := X"8FC40078";
        ram_buffer(30379) := X"0040F809";
        ram_buffer(30380) := X"00000000";
        ram_buffer(30381) := X"AFC20014";
        ram_buffer(30382) := X"8FC30014";
        ram_buffer(30383) := X"2402FFFF";
        ram_buffer(30384) := X"106200D8";
        ram_buffer(30385) := X"00000000";
        ram_buffer(30386) := X"8E020004";
        ram_buffer(30387) := X"8FC30014";
        ram_buffer(30388) := X"00000000";
        ram_buffer(30389) := X"00621023";
        ram_buffer(30390) := X"AFC20014";
        ram_buffer(30391) := X"8E020030";
        ram_buffer(30392) := X"00000000";
        ram_buffer(30393) := X"10400006";
        ram_buffer(30394) := X"00000000";
        ram_buffer(30395) := X"8E02003C";
        ram_buffer(30396) := X"8FC30014";
        ram_buffer(30397) := X"00000000";
        ram_buffer(30398) := X"00621023";
        ram_buffer(30399) := X"AFC20014";
        ram_buffer(30400) := X"8E020030";
        ram_buffer(30401) := X"00000000";
        ram_buffer(30402) := X"1040001B";
        ram_buffer(30403) := X"00000000";
        ram_buffer(30404) := X"8E020004";
        ram_buffer(30405) := X"8FC30014";
        ram_buffer(30406) := X"00000000";
        ram_buffer(30407) := X"00621021";
        ram_buffer(30408) := X"AFC20014";
        ram_buffer(30409) := X"8E020038";
        ram_buffer(30410) := X"00000000";
        ram_buffer(30411) := X"00401821";
        ram_buffer(30412) := X"8E020010";
        ram_buffer(30413) := X"00000000";
        ram_buffer(30414) := X"00621023";
        ram_buffer(30415) := X"AFC20018";
        ram_buffer(30416) := X"8FC30014";
        ram_buffer(30417) := X"8FC20018";
        ram_buffer(30418) := X"00000000";
        ram_buffer(30419) := X"00621023";
        ram_buffer(30420) := X"AFC20014";
        ram_buffer(30421) := X"8E02003C";
        ram_buffer(30422) := X"00000000";
        ram_buffer(30423) := X"00401821";
        ram_buffer(30424) := X"8FC20018";
        ram_buffer(30425) := X"00000000";
        ram_buffer(30426) := X"00431021";
        ram_buffer(30427) := X"AFC20018";
        ram_buffer(30428) := X"10000014";
        ram_buffer(30429) := X"00000000";
        ram_buffer(30430) := X"8E020000";
        ram_buffer(30431) := X"00000000";
        ram_buffer(30432) := X"00401821";
        ram_buffer(30433) := X"8E020010";
        ram_buffer(30434) := X"00000000";
        ram_buffer(30435) := X"00621023";
        ram_buffer(30436) := X"AFC20018";
        ram_buffer(30437) := X"8FC30014";
        ram_buffer(30438) := X"8FC20018";
        ram_buffer(30439) := X"00000000";
        ram_buffer(30440) := X"00621023";
        ram_buffer(30441) := X"AFC20014";
        ram_buffer(30442) := X"8E020004";
        ram_buffer(30443) := X"00000000";
        ram_buffer(30444) := X"00401821";
        ram_buffer(30445) := X"8FC20018";
        ram_buffer(30446) := X"00000000";
        ram_buffer(30447) := X"00431021";
        ram_buffer(30448) := X"AFC20018";
        ram_buffer(30449) := X"8FC30010";
        ram_buffer(30450) := X"8FC20014";
        ram_buffer(30451) := X"00000000";
        ram_buffer(30452) := X"0062102A";
        ram_buffer(30453) := X"14400035";
        ram_buffer(30454) := X"00000000";
        ram_buffer(30455) := X"8FC30014";
        ram_buffer(30456) := X"8FC20018";
        ram_buffer(30457) := X"00000000";
        ram_buffer(30458) := X"00621821";
        ram_buffer(30459) := X"8FC20010";
        ram_buffer(30460) := X"00000000";
        ram_buffer(30461) := X"0043102B";
        ram_buffer(30462) := X"1040002C";
        ram_buffer(30463) := X"00000000";
        ram_buffer(30464) := X"8FC30010";
        ram_buffer(30465) := X"8FC20014";
        ram_buffer(30466) := X"00000000";
        ram_buffer(30467) := X"0062F823";
        ram_buffer(30468) := X"8E020010";
        ram_buffer(30469) := X"03E01821";
        ram_buffer(30470) := X"00431021";
        ram_buffer(30471) := X"AE020000";
        ram_buffer(30472) := X"03E01821";
        ram_buffer(30473) := X"8FC20018";
        ram_buffer(30474) := X"00000000";
        ram_buffer(30475) := X"00431023";
        ram_buffer(30476) := X"AE020004";
        ram_buffer(30477) := X"8E020030";
        ram_buffer(30478) := X"00000000";
        ram_buffer(30479) := X"1040000C";
        ram_buffer(30480) := X"00000000";
        ram_buffer(30481) := X"8E030030";
        ram_buffer(30482) := X"26020040";
        ram_buffer(30483) := X"10620007";
        ram_buffer(30484) := X"00000000";
        ram_buffer(30485) := X"8E020030";
        ram_buffer(30486) := X"00000000";
        ram_buffer(30487) := X"00402821";
        ram_buffer(30488) := X"8FC40078";
        ram_buffer(30489) := X"0C027301";
        ram_buffer(30490) := X"00000000";
        ram_buffer(30491) := X"AE000030";
        ram_buffer(30492) := X"8603000C";
        ram_buffer(30493) := X"2402FFDF";
        ram_buffer(30494) := X"00621024";
        ram_buffer(30495) := X"00021400";
        ram_buffer(30496) := X"00021403";
        ram_buffer(30497) := X"A602000C";
        ram_buffer(30498) := X"2602005C";
        ram_buffer(30499) := X"24060008";
        ram_buffer(30500) := X"00002821";
        ram_buffer(30501) := X"00402021";
        ram_buffer(30502) := X"0C02801D";
        ram_buffer(30503) := X"00000000";
        ram_buffer(30504) := X"00001021";
        ram_buffer(30505) := X"1000009E";
        ram_buffer(30506) := X"00000000";
        ram_buffer(30507) := X"8E02004C";
        ram_buffer(30508) := X"00000000";
        ram_buffer(30509) := X"00021823";
        ram_buffer(30510) := X"8FC20010";
        ram_buffer(30511) := X"00000000";
        ram_buffer(30512) := X"00621024";
        ram_buffer(30513) := X"AFC20014";
        ram_buffer(30514) := X"8E03001C";
        ram_buffer(30515) := X"8FC20024";
        ram_buffer(30516) := X"00003821";
        ram_buffer(30517) := X"8FC60014";
        ram_buffer(30518) := X"00602821";
        ram_buffer(30519) := X"8FC40078";
        ram_buffer(30520) := X"0040F809";
        ram_buffer(30521) := X"00000000";
        ram_buffer(30522) := X"00401821";
        ram_buffer(30523) := X"2402FFFF";
        ram_buffer(30524) := X"1062004F";
        ram_buffer(30525) := X"00000000";
        ram_buffer(30526) := X"AE000004";
        ram_buffer(30527) := X"8E020010";
        ram_buffer(30528) := X"00000000";
        ram_buffer(30529) := X"AE020000";
        ram_buffer(30530) := X"8E020030";
        ram_buffer(30531) := X"00000000";
        ram_buffer(30532) := X"1040000C";
        ram_buffer(30533) := X"00000000";
        ram_buffer(30534) := X"8E030030";
        ram_buffer(30535) := X"26020040";
        ram_buffer(30536) := X"10620007";
        ram_buffer(30537) := X"00000000";
        ram_buffer(30538) := X"8E020030";
        ram_buffer(30539) := X"00000000";
        ram_buffer(30540) := X"00402821";
        ram_buffer(30541) := X"8FC40078";
        ram_buffer(30542) := X"0C027301";
        ram_buffer(30543) := X"00000000";
        ram_buffer(30544) := X"AE000030";
        ram_buffer(30545) := X"8603000C";
        ram_buffer(30546) := X"2402FFDF";
        ram_buffer(30547) := X"00621024";
        ram_buffer(30548) := X"00021400";
        ram_buffer(30549) := X"00021403";
        ram_buffer(30550) := X"A602000C";
        ram_buffer(30551) := X"8FC30010";
        ram_buffer(30552) := X"8FC20014";
        ram_buffer(30553) := X"00000000";
        ram_buffer(30554) := X"00621023";
        ram_buffer(30555) := X"AFC20018";
        ram_buffer(30556) := X"8FC20018";
        ram_buffer(30557) := X"00000000";
        ram_buffer(30558) := X"1040001B";
        ram_buffer(30559) := X"00000000";
        ram_buffer(30560) := X"02002821";
        ram_buffer(30561) := X"8FC40078";
        ram_buffer(30562) := X"0C028274";
        ram_buffer(30563) := X"00000000";
        ram_buffer(30564) := X"14400028";
        ram_buffer(30565) := X"00000000";
        ram_buffer(30566) := X"8E020004";
        ram_buffer(30567) := X"00000000";
        ram_buffer(30568) := X"00401821";
        ram_buffer(30569) := X"8FC20018";
        ram_buffer(30570) := X"00000000";
        ram_buffer(30571) := X"0062102B";
        ram_buffer(30572) := X"14400020";
        ram_buffer(30573) := X"00000000";
        ram_buffer(30574) := X"8E030000";
        ram_buffer(30575) := X"8FC20018";
        ram_buffer(30576) := X"00000000";
        ram_buffer(30577) := X"00621021";
        ram_buffer(30578) := X"AE020000";
        ram_buffer(30579) := X"8E020004";
        ram_buffer(30580) := X"00000000";
        ram_buffer(30581) := X"00401821";
        ram_buffer(30582) := X"8FC20018";
        ram_buffer(30583) := X"00000000";
        ram_buffer(30584) := X"00621023";
        ram_buffer(30585) := X"AE020004";
        ram_buffer(30586) := X"2602005C";
        ram_buffer(30587) := X"24060008";
        ram_buffer(30588) := X"00002821";
        ram_buffer(30589) := X"00402021";
        ram_buffer(30590) := X"0C02801D";
        ram_buffer(30591) := X"00000000";
        ram_buffer(30592) := X"00001021";
        ram_buffer(30593) := X"10000046";
        ram_buffer(30594) := X"00000000";
        ram_buffer(30595) := X"00000000";
        ram_buffer(30596) := X"10000008";
        ram_buffer(30597) := X"00000000";
        ram_buffer(30598) := X"00000000";
        ram_buffer(30599) := X"10000005";
        ram_buffer(30600) := X"00000000";
        ram_buffer(30601) := X"00000000";
        ram_buffer(30602) := X"10000002";
        ram_buffer(30603) := X"00000000";
        ram_buffer(30604) := X"00000000";
        ram_buffer(30605) := X"02002821";
        ram_buffer(30606) := X"8FC40078";
        ram_buffer(30607) := X"0C026EE1";
        ram_buffer(30608) := X"00000000";
        ram_buffer(30609) := X"1440000D";
        ram_buffer(30610) := X"00000000";
        ram_buffer(30611) := X"8E03001C";
        ram_buffer(30612) := X"8FC20024";
        ram_buffer(30613) := X"8FC70084";
        ram_buffer(30614) := X"8FC60080";
        ram_buffer(30615) := X"00602821";
        ram_buffer(30616) := X"8FC40078";
        ram_buffer(30617) := X"0040F809";
        ram_buffer(30618) := X"00000000";
        ram_buffer(30619) := X"00401821";
        ram_buffer(30620) := X"2402FFFF";
        ram_buffer(30621) := X"14620004";
        ram_buffer(30622) := X"00000000";
        ram_buffer(30623) := X"2402FFFF";
        ram_buffer(30624) := X"10000027";
        ram_buffer(30625) := X"00000000";
        ram_buffer(30626) := X"8E020030";
        ram_buffer(30627) := X"00000000";
        ram_buffer(30628) := X"1040000C";
        ram_buffer(30629) := X"00000000";
        ram_buffer(30630) := X"8E030030";
        ram_buffer(30631) := X"26020040";
        ram_buffer(30632) := X"10620007";
        ram_buffer(30633) := X"00000000";
        ram_buffer(30634) := X"8E020030";
        ram_buffer(30635) := X"00000000";
        ram_buffer(30636) := X"00402821";
        ram_buffer(30637) := X"8FC40078";
        ram_buffer(30638) := X"0C027301";
        ram_buffer(30639) := X"00000000";
        ram_buffer(30640) := X"AE000030";
        ram_buffer(30641) := X"8E020010";
        ram_buffer(30642) := X"00000000";
        ram_buffer(30643) := X"AE020000";
        ram_buffer(30644) := X"AE000004";
        ram_buffer(30645) := X"8603000C";
        ram_buffer(30646) := X"2402FFDF";
        ram_buffer(30647) := X"00621024";
        ram_buffer(30648) := X"00021400";
        ram_buffer(30649) := X"00021403";
        ram_buffer(30650) := X"A602000C";
        ram_buffer(30651) := X"8603000C";
        ram_buffer(30652) := X"2402F7FF";
        ram_buffer(30653) := X"00621024";
        ram_buffer(30654) := X"00021400";
        ram_buffer(30655) := X"00021403";
        ram_buffer(30656) := X"A602000C";
        ram_buffer(30657) := X"2602005C";
        ram_buffer(30658) := X"24060008";
        ram_buffer(30659) := X"00002821";
        ram_buffer(30660) := X"00402021";
        ram_buffer(30661) := X"0C02801D";
        ram_buffer(30662) := X"00000000";
        ram_buffer(30663) := X"00001021";
        ram_buffer(30664) := X"03C0E821";
        ram_buffer(30665) := X"8FBF0074";
        ram_buffer(30666) := X"8FBE0070";
        ram_buffer(30667) := X"8FB0006C";
        ram_buffer(30668) := X"27BD0078";
        ram_buffer(30669) := X"03E00008";
        ram_buffer(30670) := X"00000000";
        ram_buffer(30671) := X"27BDFFE8";
        ram_buffer(30672) := X"AFBF0014";
        ram_buffer(30673) := X"AFBE0010";
        ram_buffer(30674) := X"03A0F021";
        ram_buffer(30675) := X"00801821";
        ram_buffer(30676) := X"AFC5001C";
        ram_buffer(30677) := X"AFC60020";
        ram_buffer(30678) := X"8F828098";
        ram_buffer(30679) := X"8FC70020";
        ram_buffer(30680) := X"8FC6001C";
        ram_buffer(30681) := X"00602821";
        ram_buffer(30682) := X"00402021";
        ram_buffer(30683) := X"0C0275A1";
        ram_buffer(30684) := X"00000000";
        ram_buffer(30685) := X"03C0E821";
        ram_buffer(30686) := X"8FBF0014";
        ram_buffer(30687) := X"8FBE0010";
        ram_buffer(30688) := X"27BD0018";
        ram_buffer(30689) := X"03E00008";
        ram_buffer(30690) := X"00000000";
        ram_buffer(30691) := X"27BDFFE0";
        ram_buffer(30692) := X"AFBF001C";
        ram_buffer(30693) := X"AFBE0018";
        ram_buffer(30694) := X"03A0F021";
        ram_buffer(30695) := X"AFC40020";
        ram_buffer(30696) := X"AFC50024";
        ram_buffer(30697) := X"AFC60028";
        ram_buffer(30698) := X"AF8081EC";
        ram_buffer(30699) := X"8FC50028";
        ram_buffer(30700) := X"8FC40024";
        ram_buffer(30701) := X"0C02FB83";
        ram_buffer(30702) := X"00000000";
        ram_buffer(30703) := X"AFC20010";
        ram_buffer(30704) := X"8FC30010";
        ram_buffer(30705) := X"2402FFFF";
        ram_buffer(30706) := X"14620009";
        ram_buffer(30707) := X"00000000";
        ram_buffer(30708) := X"8F8281EC";
        ram_buffer(30709) := X"00000000";
        ram_buffer(30710) := X"10400005";
        ram_buffer(30711) := X"00000000";
        ram_buffer(30712) := X"8F8381EC";
        ram_buffer(30713) := X"8FC20020";
        ram_buffer(30714) := X"00000000";
        ram_buffer(30715) := X"AC430000";
        ram_buffer(30716) := X"8FC20010";
        ram_buffer(30717) := X"03C0E821";
        ram_buffer(30718) := X"8FBF001C";
        ram_buffer(30719) := X"8FBE0018";
        ram_buffer(30720) := X"27BD0020";
        ram_buffer(30721) := X"03E00008";
        ram_buffer(30722) := X"00000000";
        ram_buffer(30723) := X"27BDFFD0";
        ram_buffer(30724) := X"AFBF002C";
        ram_buffer(30725) := X"AFBE0028";
        ram_buffer(30726) := X"AFB40024";
        ram_buffer(30727) := X"AFB30020";
        ram_buffer(30728) := X"AFB2001C";
        ram_buffer(30729) := X"AFB10018";
        ram_buffer(30730) := X"AFB00014";
        ram_buffer(30731) := X"03A0F021";
        ram_buffer(30732) := X"AFC40030";
        ram_buffer(30733) := X"00A0A021";
        ram_buffer(30734) := X"00009821";
        ram_buffer(30735) := X"8FC20030";
        ram_buffer(30736) := X"00000000";
        ram_buffer(30737) := X"245102E0";
        ram_buffer(30738) := X"1000001B";
        ram_buffer(30739) := X"00000000";
        ram_buffer(30740) := X"8E300008";
        ram_buffer(30741) := X"8E320004";
        ram_buffer(30742) := X"10000012";
        ram_buffer(30743) := X"00000000";
        ram_buffer(30744) := X"8602000C";
        ram_buffer(30745) := X"00000000";
        ram_buffer(30746) := X"1040000D";
        ram_buffer(30747) := X"00000000";
        ram_buffer(30748) := X"8603000C";
        ram_buffer(30749) := X"24020001";
        ram_buffer(30750) := X"10620009";
        ram_buffer(30751) := X"00000000";
        ram_buffer(30752) := X"8603000E";
        ram_buffer(30753) := X"2402FFFF";
        ram_buffer(30754) := X"10620005";
        ram_buffer(30755) := X"00000000";
        ram_buffer(30756) := X"02002021";
        ram_buffer(30757) := X"0280F809";
        ram_buffer(30758) := X"00000000";
        ram_buffer(30759) := X"02629825";
        ram_buffer(30760) := X"26100068";
        ram_buffer(30761) := X"2652FFFF";
        ram_buffer(30762) := X"0641FFED";
        ram_buffer(30763) := X"00000000";
        ram_buffer(30764) := X"8E310000";
        ram_buffer(30765) := X"00000000";
        ram_buffer(30766) := X"1620FFE5";
        ram_buffer(30767) := X"00000000";
        ram_buffer(30768) := X"02601021";
        ram_buffer(30769) := X"03C0E821";
        ram_buffer(30770) := X"8FBF002C";
        ram_buffer(30771) := X"8FBE0028";
        ram_buffer(30772) := X"8FB40024";
        ram_buffer(30773) := X"8FB30020";
        ram_buffer(30774) := X"8FB2001C";
        ram_buffer(30775) := X"8FB10018";
        ram_buffer(30776) := X"8FB00014";
        ram_buffer(30777) := X"27BD0030";
        ram_buffer(30778) := X"03E00008";
        ram_buffer(30779) := X"00000000";
        ram_buffer(30780) := X"27BDFFD0";
        ram_buffer(30781) := X"AFBF002C";
        ram_buffer(30782) := X"AFBE0028";
        ram_buffer(30783) := X"AFB40024";
        ram_buffer(30784) := X"AFB30020";
        ram_buffer(30785) := X"AFB2001C";
        ram_buffer(30786) := X"AFB10018";
        ram_buffer(30787) := X"AFB00014";
        ram_buffer(30788) := X"03A0F021";
        ram_buffer(30789) := X"AFC40030";
        ram_buffer(30790) := X"00A0A021";
        ram_buffer(30791) := X"00009821";
        ram_buffer(30792) := X"8FC20030";
        ram_buffer(30793) := X"00000000";
        ram_buffer(30794) := X"245102E0";
        ram_buffer(30795) := X"1000001C";
        ram_buffer(30796) := X"00000000";
        ram_buffer(30797) := X"8E300008";
        ram_buffer(30798) := X"8E320004";
        ram_buffer(30799) := X"10000013";
        ram_buffer(30800) := X"00000000";
        ram_buffer(30801) := X"8602000C";
        ram_buffer(30802) := X"00000000";
        ram_buffer(30803) := X"1040000E";
        ram_buffer(30804) := X"00000000";
        ram_buffer(30805) := X"8603000C";
        ram_buffer(30806) := X"24020001";
        ram_buffer(30807) := X"1062000A";
        ram_buffer(30808) := X"00000000";
        ram_buffer(30809) := X"8603000E";
        ram_buffer(30810) := X"2402FFFF";
        ram_buffer(30811) := X"10620006";
        ram_buffer(30812) := X"00000000";
        ram_buffer(30813) := X"02002821";
        ram_buffer(30814) := X"8FC40030";
        ram_buffer(30815) := X"0280F809";
        ram_buffer(30816) := X"00000000";
        ram_buffer(30817) := X"02629825";
        ram_buffer(30818) := X"26100068";
        ram_buffer(30819) := X"2652FFFF";
        ram_buffer(30820) := X"0641FFEC";
        ram_buffer(30821) := X"00000000";
        ram_buffer(30822) := X"8E310000";
        ram_buffer(30823) := X"00000000";
        ram_buffer(30824) := X"1620FFE4";
        ram_buffer(30825) := X"00000000";
        ram_buffer(30826) := X"02601021";
        ram_buffer(30827) := X"03C0E821";
        ram_buffer(30828) := X"8FBF002C";
        ram_buffer(30829) := X"8FBE0028";
        ram_buffer(30830) := X"8FB40024";
        ram_buffer(30831) := X"8FB30020";
        ram_buffer(30832) := X"8FB2001C";
        ram_buffer(30833) := X"8FB10018";
        ram_buffer(30834) := X"8FB00014";
        ram_buffer(30835) := X"27BD0030";
        ram_buffer(30836) := X"03E00008";
        ram_buffer(30837) := X"00000000";
        ram_buffer(30838) := X"27BDFFC8";
        ram_buffer(30839) := X"AFBF0034";
        ram_buffer(30840) := X"AFBE0030";
        ram_buffer(30841) := X"03A0F021";
        ram_buffer(30842) := X"AFC40038";
        ram_buffer(30843) := X"AFC5003C";
        ram_buffer(30844) := X"AFC60040";
        ram_buffer(30845) := X"AFC70044";
        ram_buffer(30846) := X"8FC2003C";
        ram_buffer(30847) := X"00000000";
        ram_buffer(30848) := X"AFC20024";
        ram_buffer(30849) := X"8FC30044";
        ram_buffer(30850) := X"8FC20040";
        ram_buffer(30851) := X"00000000";
        ram_buffer(30852) := X"00620018";
        ram_buffer(30853) := X"00001012";
        ram_buffer(30854) := X"AFC20010";
        ram_buffer(30855) := X"8FC20010";
        ram_buffer(30856) := X"00000000";
        ram_buffer(30857) := X"AFC20028";
        ram_buffer(30858) := X"8FC20028";
        ram_buffer(30859) := X"00000000";
        ram_buffer(30860) := X"AFC20020";
        ram_buffer(30861) := X"27C20024";
        ram_buffer(30862) := X"AFC20018";
        ram_buffer(30863) := X"24020001";
        ram_buffer(30864) := X"AFC2001C";
        ram_buffer(30865) := X"8FC20038";
        ram_buffer(30866) := X"00000000";
        ram_buffer(30867) := X"AFC20014";
        ram_buffer(30868) := X"8FC20014";
        ram_buffer(30869) := X"00000000";
        ram_buffer(30870) := X"1040000A";
        ram_buffer(30871) := X"00000000";
        ram_buffer(30872) := X"8FC20014";
        ram_buffer(30873) := X"00000000";
        ram_buffer(30874) := X"8C420038";
        ram_buffer(30875) := X"00000000";
        ram_buffer(30876) := X"14400004";
        ram_buffer(30877) := X"00000000";
        ram_buffer(30878) := X"8FC40014";
        ram_buffer(30879) := X"0C027069";
        ram_buffer(30880) := X"00000000";
        ram_buffer(30881) := X"8FC20048";
        ram_buffer(30882) := X"00000000";
        ram_buffer(30883) := X"8442000C";
        ram_buffer(30884) := X"00000000";
        ram_buffer(30885) := X"3042FFFF";
        ram_buffer(30886) := X"30422000";
        ram_buffer(30887) := X"14400013";
        ram_buffer(30888) := X"00000000";
        ram_buffer(30889) := X"8FC20048";
        ram_buffer(30890) := X"00000000";
        ram_buffer(30891) := X"8442000C";
        ram_buffer(30892) := X"00000000";
        ram_buffer(30893) := X"34422000";
        ram_buffer(30894) := X"00021C00";
        ram_buffer(30895) := X"00031C03";
        ram_buffer(30896) := X"8FC20048";
        ram_buffer(30897) := X"00000000";
        ram_buffer(30898) := X"A443000C";
        ram_buffer(30899) := X"8FC20048";
        ram_buffer(30900) := X"00000000";
        ram_buffer(30901) := X"8C430064";
        ram_buffer(30902) := X"2402DFFF";
        ram_buffer(30903) := X"00621824";
        ram_buffer(30904) := X"8FC20048";
        ram_buffer(30905) := X"00000000";
        ram_buffer(30906) := X"AC430064";
        ram_buffer(30907) := X"27C20018";
        ram_buffer(30908) := X"00403021";
        ram_buffer(30909) := X"8FC50048";
        ram_buffer(30910) := X"8FC40038";
        ram_buffer(30911) := X"0C02B89A";
        ram_buffer(30912) := X"00000000";
        ram_buffer(30913) := X"14400004";
        ram_buffer(30914) := X"00000000";
        ram_buffer(30915) := X"8FC20044";
        ram_buffer(30916) := X"1000000C";
        ram_buffer(30917) := X"00000000";
        ram_buffer(30918) := X"8FC20020";
        ram_buffer(30919) := X"8FC30010";
        ram_buffer(30920) := X"00000000";
        ram_buffer(30921) := X"00621823";
        ram_buffer(30922) := X"8FC20040";
        ram_buffer(30923) := X"00000000";
        ram_buffer(30924) := X"14400002";
        ram_buffer(30925) := X"0062001B";
        ram_buffer(30926) := X"0007000D";
        ram_buffer(30927) := X"00001010";
        ram_buffer(30928) := X"00001012";
        ram_buffer(30929) := X"03C0E821";
        ram_buffer(30930) := X"8FBF0034";
        ram_buffer(30931) := X"8FBE0030";
        ram_buffer(30932) := X"27BD0038";
        ram_buffer(30933) := X"03E00008";
        ram_buffer(30934) := X"00000000";
        ram_buffer(30935) := X"27BDFFE0";
        ram_buffer(30936) := X"AFBF001C";
        ram_buffer(30937) := X"AFBE0018";
        ram_buffer(30938) := X"03A0F021";
        ram_buffer(30939) := X"AFC40020";
        ram_buffer(30940) := X"AFC50024";
        ram_buffer(30941) := X"AFC60028";
        ram_buffer(30942) := X"AFC7002C";
        ram_buffer(30943) := X"8F838098";
        ram_buffer(30944) := X"8FC2002C";
        ram_buffer(30945) := X"00000000";
        ram_buffer(30946) := X"AFA20010";
        ram_buffer(30947) := X"8FC70028";
        ram_buffer(30948) := X"8FC60024";
        ram_buffer(30949) := X"8FC50020";
        ram_buffer(30950) := X"00602021";
        ram_buffer(30951) := X"0C027876";
        ram_buffer(30952) := X"00000000";
        ram_buffer(30953) := X"03C0E821";
        ram_buffer(30954) := X"8FBF001C";
        ram_buffer(30955) := X"8FBE0018";
        ram_buffer(30956) := X"27BD0020";
        ram_buffer(30957) := X"03E00008";
        ram_buffer(30958) := X"00000000";
        ram_buffer(30959) := X"27BDFFE8";
        ram_buffer(30960) := X"AFBF0014";
        ram_buffer(30961) := X"AFBE0010";
        ram_buffer(30962) := X"03A0F021";
        ram_buffer(30963) := X"00801821";
        ram_buffer(30964) := X"AFC5001C";
        ram_buffer(30965) := X"8F828098";
        ram_buffer(30966) := X"8FC6001C";
        ram_buffer(30967) := X"00602821";
        ram_buffer(30968) := X"00402021";
        ram_buffer(30969) := X"0C027913";
        ram_buffer(30970) := X"00000000";
        ram_buffer(30971) := X"03C0E821";
        ram_buffer(30972) := X"8FBF0014";
        ram_buffer(30973) := X"8FBE0010";
        ram_buffer(30974) := X"27BD0018";
        ram_buffer(30975) := X"03E00008";
        ram_buffer(30976) := X"00000000";
        ram_buffer(30977) := X"27BDFFE0";
        ram_buffer(30978) := X"AFBF001C";
        ram_buffer(30979) := X"AFBE0018";
        ram_buffer(30980) := X"03A0F021";
        ram_buffer(30981) := X"AFC40020";
        ram_buffer(30982) := X"8F828098";
        ram_buffer(30983) := X"27C30010";
        ram_buffer(30984) := X"00603021";
        ram_buffer(30985) := X"8FC50020";
        ram_buffer(30986) := X"00402021";
        ram_buffer(30987) := X"0C027913";
        ram_buffer(30988) := X"00000000";
        ram_buffer(30989) := X"03C0E821";
        ram_buffer(30990) := X"8FBF001C";
        ram_buffer(30991) := X"8FBE0018";
        ram_buffer(30992) := X"27BD0020";
        ram_buffer(30993) := X"03E00008";
        ram_buffer(30994) := X"00000000";
        ram_buffer(30995) := X"27BDFFD0";
        ram_buffer(30996) := X"AFBF002C";
        ram_buffer(30997) := X"AFBE0028";
        ram_buffer(30998) := X"AFB20024";
        ram_buffer(30999) := X"AFB10020";
        ram_buffer(31000) := X"AFB0001C";
        ram_buffer(31001) := X"03A0F021";
        ram_buffer(31002) := X"AFC40030";
        ram_buffer(31003) := X"00A08821";
        ram_buffer(31004) := X"AFC60038";
        ram_buffer(31005) := X"8FC40030";
        ram_buffer(31006) := X"0C02B832";
        ram_buffer(31007) := X"00000000";
        ram_buffer(31008) := X"8F828094";
        ram_buffer(31009) := X"00000000";
        ram_buffer(31010) := X"8C420000";
        ram_buffer(31011) := X"00000000";
        ram_buffer(31012) := X"14400007";
        ram_buffer(31013) := X"00000000";
        ram_buffer(31014) := X"8FC40030";
        ram_buffer(31015) := X"0C02B83C";
        ram_buffer(31016) := X"00000000";
        ram_buffer(31017) := X"00001021";
        ram_buffer(31018) := X"10000053";
        ram_buffer(31019) := X"00000000";
        ram_buffer(31020) := X"AFD10010";
        ram_buffer(31021) := X"10000005";
        ram_buffer(31022) := X"00000000";
        ram_buffer(31023) := X"8FC20010";
        ram_buffer(31024) := X"00000000";
        ram_buffer(31025) := X"24420001";
        ram_buffer(31026) := X"AFC20010";
        ram_buffer(31027) := X"8FC20010";
        ram_buffer(31028) := X"00000000";
        ram_buffer(31029) := X"80420000";
        ram_buffer(31030) := X"00000000";
        ram_buffer(31031) := X"10400007";
        ram_buffer(31032) := X"00000000";
        ram_buffer(31033) := X"8FC20010";
        ram_buffer(31034) := X"00000000";
        ram_buffer(31035) := X"80430000";
        ram_buffer(31036) := X"2402003D";
        ram_buffer(31037) := X"1462FFF1";
        ram_buffer(31038) := X"00000000";
        ram_buffer(31039) := X"8FC20010";
        ram_buffer(31040) := X"00000000";
        ram_buffer(31041) := X"80430000";
        ram_buffer(31042) := X"2402003D";
        ram_buffer(31043) := X"10620036";
        ram_buffer(31044) := X"00000000";
        ram_buffer(31045) := X"8FC20010";
        ram_buffer(31046) := X"02201821";
        ram_buffer(31047) := X"00439023";
        ram_buffer(31048) := X"8F828094";
        ram_buffer(31049) := X"00000000";
        ram_buffer(31050) := X"8C500000";
        ram_buffer(31051) := X"1000002A";
        ram_buffer(31052) := X"00000000";
        ram_buffer(31053) := X"8E020000";
        ram_buffer(31054) := X"02401821";
        ram_buffer(31055) := X"00603021";
        ram_buffer(31056) := X"02202821";
        ram_buffer(31057) := X"00402021";
        ram_buffer(31058) := X"0C028525";
        ram_buffer(31059) := X"00000000";
        ram_buffer(31060) := X"14400020";
        ram_buffer(31061) := X"00000000";
        ram_buffer(31062) := X"8E020000";
        ram_buffer(31063) := X"02401821";
        ram_buffer(31064) := X"00431021";
        ram_buffer(31065) := X"AFC20010";
        ram_buffer(31066) := X"8FC20010";
        ram_buffer(31067) := X"00000000";
        ram_buffer(31068) := X"80430000";
        ram_buffer(31069) := X"2402003D";
        ram_buffer(31070) := X"14620016";
        ram_buffer(31071) := X"00000000";
        ram_buffer(31072) := X"02001821";
        ram_buffer(31073) := X"8F828094";
        ram_buffer(31074) := X"00000000";
        ram_buffer(31075) := X"8C420000";
        ram_buffer(31076) := X"00000000";
        ram_buffer(31077) := X"00621023";
        ram_buffer(31078) := X"00021083";
        ram_buffer(31079) := X"00401821";
        ram_buffer(31080) := X"8FC20038";
        ram_buffer(31081) := X"00000000";
        ram_buffer(31082) := X"AC430000";
        ram_buffer(31083) := X"8FC40030";
        ram_buffer(31084) := X"0C02B83C";
        ram_buffer(31085) := X"00000000";
        ram_buffer(31086) := X"8FC20010";
        ram_buffer(31087) := X"00000000";
        ram_buffer(31088) := X"24420001";
        ram_buffer(31089) := X"AFC20010";
        ram_buffer(31090) := X"8FC20010";
        ram_buffer(31091) := X"1000000A";
        ram_buffer(31092) := X"00000000";
        ram_buffer(31093) := X"26100004";
        ram_buffer(31094) := X"8E020000";
        ram_buffer(31095) := X"00000000";
        ram_buffer(31096) := X"1440FFD4";
        ram_buffer(31097) := X"00000000";
        ram_buffer(31098) := X"8FC40030";
        ram_buffer(31099) := X"0C02B83C";
        ram_buffer(31100) := X"00000000";
        ram_buffer(31101) := X"00001021";
        ram_buffer(31102) := X"03C0E821";
        ram_buffer(31103) := X"8FBF002C";
        ram_buffer(31104) := X"8FBE0028";
        ram_buffer(31105) := X"8FB20024";
        ram_buffer(31106) := X"8FB10020";
        ram_buffer(31107) := X"8FB0001C";
        ram_buffer(31108) := X"27BD0030";
        ram_buffer(31109) := X"03E00008";
        ram_buffer(31110) := X"00000000";
        ram_buffer(31111) := X"27BDFFE0";
        ram_buffer(31112) := X"AFBF001C";
        ram_buffer(31113) := X"AFBE0018";
        ram_buffer(31114) := X"03A0F021";
        ram_buffer(31115) := X"AFC40020";
        ram_buffer(31116) := X"AFC50024";
        ram_buffer(31117) := X"27C20010";
        ram_buffer(31118) := X"00403021";
        ram_buffer(31119) := X"8FC50024";
        ram_buffer(31120) := X"8FC40020";
        ram_buffer(31121) := X"0C027913";
        ram_buffer(31122) := X"00000000";
        ram_buffer(31123) := X"03C0E821";
        ram_buffer(31124) := X"8FBF001C";
        ram_buffer(31125) := X"8FBE0018";
        ram_buffer(31126) := X"27BD0020";
        ram_buffer(31127) := X"03E00008";
        ram_buffer(31128) := X"00000000";
        ram_buffer(31129) := X"27BDFF98";
        ram_buffer(31130) := X"AFBF0064";
        ram_buffer(31131) := X"AFBE0060";
        ram_buffer(31132) := X"AFB3005C";
        ram_buffer(31133) := X"AFB20058";
        ram_buffer(31134) := X"AFB10054";
        ram_buffer(31135) := X"AFB00050";
        ram_buffer(31136) := X"03A0F021";
        ram_buffer(31137) := X"AFC40068";
        ram_buffer(31138) := X"00A08021";
        ram_buffer(31139) := X"8602000C";
        ram_buffer(31140) := X"00000000";
        ram_buffer(31141) := X"3042FFFF";
        ram_buffer(31142) := X"30420002";
        ram_buffer(31143) := X"1040000A";
        ram_buffer(31144) := X"00000000";
        ram_buffer(31145) := X"26020043";
        ram_buffer(31146) := X"AE020000";
        ram_buffer(31147) := X"8E020000";
        ram_buffer(31148) := X"00000000";
        ram_buffer(31149) := X"AE020010";
        ram_buffer(31150) := X"24020001";
        ram_buffer(31151) := X"AE020014";
        ram_buffer(31152) := X"10000082";
        ram_buffer(31153) := X"00000000";
        ram_buffer(31154) := X"8602000E";
        ram_buffer(31155) := X"00000000";
        ram_buffer(31156) := X"0440000C";
        ram_buffer(31157) := X"00000000";
        ram_buffer(31158) := X"8602000E";
        ram_buffer(31159) := X"00000000";
        ram_buffer(31160) := X"00401821";
        ram_buffer(31161) := X"27C20010";
        ram_buffer(31162) := X"00403021";
        ram_buffer(31163) := X"00602821";
        ram_buffer(31164) := X"8FC40068";
        ram_buffer(31165) := X"0C0277E3";
        ram_buffer(31166) := X"00000000";
        ram_buffer(31167) := X"04410014";
        ram_buffer(31168) := X"00000000";
        ram_buffer(31169) := X"00009821";
        ram_buffer(31170) := X"8602000C";
        ram_buffer(31171) := X"00000000";
        ram_buffer(31172) := X"3042FFFF";
        ram_buffer(31173) := X"30420080";
        ram_buffer(31174) := X"10400004";
        ram_buffer(31175) := X"00000000";
        ram_buffer(31176) := X"24110040";
        ram_buffer(31177) := X"10000002";
        ram_buffer(31178) := X"00000000";
        ram_buffer(31179) := X"24110400";
        ram_buffer(31180) := X"8602000C";
        ram_buffer(31181) := X"00000000";
        ram_buffer(31182) := X"34420800";
        ram_buffer(31183) := X"00021400";
        ram_buffer(31184) := X"00021403";
        ram_buffer(31185) := X"A602000C";
        ram_buffer(31186) := X"10000024";
        ram_buffer(31187) := X"00000000";
        ram_buffer(31188) := X"8FC20014";
        ram_buffer(31189) := X"00000000";
        ram_buffer(31190) := X"3042F000";
        ram_buffer(31191) := X"38422000";
        ram_buffer(31192) := X"2C420001";
        ram_buffer(31193) := X"304200FF";
        ram_buffer(31194) := X"00409821";
        ram_buffer(31195) := X"24110400";
        ram_buffer(31196) := X"8FC20014";
        ram_buffer(31197) := X"00000000";
        ram_buffer(31198) := X"3043F000";
        ram_buffer(31199) := X"34028000";
        ram_buffer(31200) := X"14620010";
        ram_buffer(31201) := X"00000000";
        ram_buffer(31202) := X"8E030028";
        ram_buffer(31203) := X"3C02100A";
        ram_buffer(31204) := X"24421360";
        ram_buffer(31205) := X"1462000B";
        ram_buffer(31206) := X"00000000";
        ram_buffer(31207) := X"8602000C";
        ram_buffer(31208) := X"00000000";
        ram_buffer(31209) := X"34420400";
        ram_buffer(31210) := X"00021400";
        ram_buffer(31211) := X"00021403";
        ram_buffer(31212) := X"A602000C";
        ram_buffer(31213) := X"24020400";
        ram_buffer(31214) := X"AE02004C";
        ram_buffer(31215) := X"10000007";
        ram_buffer(31216) := X"00000000";
        ram_buffer(31217) := X"8602000C";
        ram_buffer(31218) := X"00000000";
        ram_buffer(31219) := X"34420800";
        ram_buffer(31220) := X"00021400";
        ram_buffer(31221) := X"00021403";
        ram_buffer(31222) := X"A602000C";
        ram_buffer(31223) := X"02202821";
        ram_buffer(31224) := X"8FC40068";
        ram_buffer(31225) := X"0C027B8F";
        ram_buffer(31226) := X"00000000";
        ram_buffer(31227) := X"00409021";
        ram_buffer(31228) := X"16400016";
        ram_buffer(31229) := X"00000000";
        ram_buffer(31230) := X"8602000C";
        ram_buffer(31231) := X"00000000";
        ram_buffer(31232) := X"3042FFFF";
        ram_buffer(31233) := X"30420200";
        ram_buffer(31234) := X"14400030";
        ram_buffer(31235) := X"00000000";
        ram_buffer(31236) := X"8602000C";
        ram_buffer(31237) := X"00000000";
        ram_buffer(31238) := X"34420002";
        ram_buffer(31239) := X"00021400";
        ram_buffer(31240) := X"00021403";
        ram_buffer(31241) := X"A602000C";
        ram_buffer(31242) := X"26020043";
        ram_buffer(31243) := X"AE020000";
        ram_buffer(31244) := X"8E020000";
        ram_buffer(31245) := X"00000000";
        ram_buffer(31246) := X"AE020010";
        ram_buffer(31247) := X"24020001";
        ram_buffer(31248) := X"AE020014";
        ram_buffer(31249) := X"10000021";
        ram_buffer(31250) := X"00000000";
        ram_buffer(31251) := X"8FC20068";
        ram_buffer(31252) := X"3C03100A";
        ram_buffer(31253) := X"2463C118";
        ram_buffer(31254) := X"AC43003C";
        ram_buffer(31255) := X"8602000C";
        ram_buffer(31256) := X"00000000";
        ram_buffer(31257) := X"34420080";
        ram_buffer(31258) := X"00021400";
        ram_buffer(31259) := X"00021403";
        ram_buffer(31260) := X"A602000C";
        ram_buffer(31261) := X"AE120000";
        ram_buffer(31262) := X"8E020000";
        ram_buffer(31263) := X"00000000";
        ram_buffer(31264) := X"AE020010";
        ram_buffer(31265) := X"02201021";
        ram_buffer(31266) := X"AE020014";
        ram_buffer(31267) := X"1260000F";
        ram_buffer(31268) := X"00000000";
        ram_buffer(31269) := X"8602000E";
        ram_buffer(31270) := X"00000000";
        ram_buffer(31271) := X"00402821";
        ram_buffer(31272) := X"8FC40068";
        ram_buffer(31273) := X"0C02BA9C";
        ram_buffer(31274) := X"00000000";
        ram_buffer(31275) := X"10400007";
        ram_buffer(31276) := X"00000000";
        ram_buffer(31277) := X"8602000C";
        ram_buffer(31278) := X"00000000";
        ram_buffer(31279) := X"34420001";
        ram_buffer(31280) := X"00021400";
        ram_buffer(31281) := X"00021403";
        ram_buffer(31282) := X"A602000C";
        ram_buffer(31283) := X"03C0E821";
        ram_buffer(31284) := X"8FBF0064";
        ram_buffer(31285) := X"8FBE0060";
        ram_buffer(31286) := X"8FB3005C";
        ram_buffer(31287) := X"8FB20058";
        ram_buffer(31288) := X"8FB10054";
        ram_buffer(31289) := X"8FB00050";
        ram_buffer(31290) := X"27BD0068";
        ram_buffer(31291) := X"03E00008";
        ram_buffer(31292) := X"00000000";
        ram_buffer(31293) := X"27BDFFE8";
        ram_buffer(31294) := X"AFBF0014";
        ram_buffer(31295) := X"AFBE0010";
        ram_buffer(31296) := X"03A0F021";
        ram_buffer(31297) := X"AFC40018";
        ram_buffer(31298) := X"8F828098";
        ram_buffer(31299) := X"8FC50018";
        ram_buffer(31300) := X"00402021";
        ram_buffer(31301) := X"0C027B8F";
        ram_buffer(31302) := X"00000000";
        ram_buffer(31303) := X"03C0E821";
        ram_buffer(31304) := X"8FBF0014";
        ram_buffer(31305) := X"8FBE0010";
        ram_buffer(31306) := X"27BD0018";
        ram_buffer(31307) := X"03E00008";
        ram_buffer(31308) := X"00000000";
        ram_buffer(31309) := X"27BDFFE8";
        ram_buffer(31310) := X"AFBF0014";
        ram_buffer(31311) := X"AFBE0010";
        ram_buffer(31312) := X"03A0F021";
        ram_buffer(31313) := X"AFC40018";
        ram_buffer(31314) := X"8F828098";
        ram_buffer(31315) := X"8FC50018";
        ram_buffer(31316) := X"00402021";
        ram_buffer(31317) := X"0C027301";
        ram_buffer(31318) := X"00000000";
        ram_buffer(31319) := X"00000000";
        ram_buffer(31320) := X"03C0E821";
        ram_buffer(31321) := X"8FBF0014";
        ram_buffer(31322) := X"8FBE0010";
        ram_buffer(31323) := X"27BD0018";
        ram_buffer(31324) := X"03E00008";
        ram_buffer(31325) := X"00000000";
        ram_buffer(31326) := X"27BDFFB8";
        ram_buffer(31327) := X"AFBF0044";
        ram_buffer(31328) := X"AFBE0040";
        ram_buffer(31329) := X"03A0F021";
        ram_buffer(31330) := X"AFC40048";
        ram_buffer(31331) := X"AFC5004C";
        ram_buffer(31332) := X"AFC00020";
        ram_buffer(31333) := X"3C02100D";
        ram_buffer(31334) := X"2442CBE0";
        ram_buffer(31335) := X"8C420008";
        ram_buffer(31336) := X"00000000";
        ram_buffer(31337) := X"AFC20024";
        ram_buffer(31338) := X"8FC20024";
        ram_buffer(31339) := X"00000000";
        ram_buffer(31340) := X"8C430004";
        ram_buffer(31341) := X"2402FFFC";
        ram_buffer(31342) := X"00621024";
        ram_buffer(31343) := X"AFC20028";
        ram_buffer(31344) := X"8FC30024";
        ram_buffer(31345) := X"8FC20028";
        ram_buffer(31346) := X"00000000";
        ram_buffer(31347) := X"00621021";
        ram_buffer(31348) := X"AFC2002C";
        ram_buffer(31349) := X"8F8381B4";
        ram_buffer(31350) := X"8FC2004C";
        ram_buffer(31351) := X"00000000";
        ram_buffer(31352) := X"00621021";
        ram_buffer(31353) := X"24420010";
        ram_buffer(31354) := X"AFC2001C";
        ram_buffer(31355) := X"24021000";
        ram_buffer(31356) := X"AFC20030";
        ram_buffer(31357) := X"8F8380A4";
        ram_buffer(31358) := X"2402FFFF";
        ram_buffer(31359) := X"1062000B";
        ram_buffer(31360) := X"00000000";
        ram_buffer(31361) := X"8FC30030";
        ram_buffer(31362) := X"8FC2001C";
        ram_buffer(31363) := X"00000000";
        ram_buffer(31364) := X"00621021";
        ram_buffer(31365) := X"2443FFFF";
        ram_buffer(31366) := X"8FC20030";
        ram_buffer(31367) := X"00000000";
        ram_buffer(31368) := X"00021023";
        ram_buffer(31369) := X"00621024";
        ram_buffer(31370) := X"AFC2001C";
        ram_buffer(31371) := X"8FC2001C";
        ram_buffer(31372) := X"00000000";
        ram_buffer(31373) := X"00402821";
        ram_buffer(31374) := X"8FC40048";
        ram_buffer(31375) := X"0C028390";
        ram_buffer(31376) := X"00000000";
        ram_buffer(31377) := X"AFC20010";
        ram_buffer(31378) := X"8FC30010";
        ram_buffer(31379) := X"2402FFFF";
        ram_buffer(31380) := X"106200F3";
        ram_buffer(31381) := X"00000000";
        ram_buffer(31382) := X"8FC30010";
        ram_buffer(31383) := X"8FC2002C";
        ram_buffer(31384) := X"00000000";
        ram_buffer(31385) := X"0062102B";
        ram_buffer(31386) := X"10400007";
        ram_buffer(31387) := X"00000000";
        ram_buffer(31388) := X"3C02100D";
        ram_buffer(31389) := X"2442CBE0";
        ram_buffer(31390) := X"8FC30024";
        ram_buffer(31391) := X"00000000";
        ram_buffer(31392) := X"146200E7";
        ram_buffer(31393) := X"00000000";
        ram_buffer(31394) := X"3C02100D";
        ram_buffer(31395) := X"8C42D260";
        ram_buffer(31396) := X"00000000";
        ram_buffer(31397) := X"00401821";
        ram_buffer(31398) := X"8FC2001C";
        ram_buffer(31399) := X"00000000";
        ram_buffer(31400) := X"00621021";
        ram_buffer(31401) := X"00401821";
        ram_buffer(31402) := X"3C02100D";
        ram_buffer(31403) := X"AC43D260";
        ram_buffer(31404) := X"8FC30010";
        ram_buffer(31405) := X"8FC2002C";
        ram_buffer(31406) := X"00000000";
        ram_buffer(31407) := X"14620017";
        ram_buffer(31408) := X"00000000";
        ram_buffer(31409) := X"8FC20030";
        ram_buffer(31410) := X"00000000";
        ram_buffer(31411) := X"2443FFFF";
        ram_buffer(31412) := X"8FC2002C";
        ram_buffer(31413) := X"00000000";
        ram_buffer(31414) := X"00621024";
        ram_buffer(31415) := X"1440000F";
        ram_buffer(31416) := X"00000000";
        ram_buffer(31417) := X"8FC3001C";
        ram_buffer(31418) := X"8FC20028";
        ram_buffer(31419) := X"00000000";
        ram_buffer(31420) := X"00621021";
        ram_buffer(31421) := X"AFC20034";
        ram_buffer(31422) := X"3C02100D";
        ram_buffer(31423) := X"2442CBE0";
        ram_buffer(31424) := X"8C420008";
        ram_buffer(31425) := X"8FC30034";
        ram_buffer(31426) := X"00000000";
        ram_buffer(31427) := X"34630001";
        ram_buffer(31428) := X"AC430004";
        ram_buffer(31429) := X"100000A6";
        ram_buffer(31430) := X"00000000";
        ram_buffer(31431) := X"8F8380A4";
        ram_buffer(31432) := X"2402FFFF";
        ram_buffer(31433) := X"14620006";
        ram_buffer(31434) := X"00000000";
        ram_buffer(31435) := X"8FC20010";
        ram_buffer(31436) := X"00000000";
        ram_buffer(31437) := X"AF8280A4";
        ram_buffer(31438) := X"1000000A";
        ram_buffer(31439) := X"00000000";
        ram_buffer(31440) := X"3C02100D";
        ram_buffer(31441) := X"8C43D260";
        ram_buffer(31442) := X"8FC40010";
        ram_buffer(31443) := X"8FC2002C";
        ram_buffer(31444) := X"00000000";
        ram_buffer(31445) := X"00821023";
        ram_buffer(31446) := X"00621821";
        ram_buffer(31447) := X"3C02100D";
        ram_buffer(31448) := X"AC43D260";
        ram_buffer(31449) := X"8FC20010";
        ram_buffer(31450) := X"00000000";
        ram_buffer(31451) := X"24420008";
        ram_buffer(31452) := X"30420007";
        ram_buffer(31453) := X"AFC20038";
        ram_buffer(31454) := X"8FC20038";
        ram_buffer(31455) := X"00000000";
        ram_buffer(31456) := X"1040000D";
        ram_buffer(31457) := X"00000000";
        ram_buffer(31458) := X"24030008";
        ram_buffer(31459) := X"8FC20038";
        ram_buffer(31460) := X"00000000";
        ram_buffer(31461) := X"00621023";
        ram_buffer(31462) := X"AFC20014";
        ram_buffer(31463) := X"8FC30010";
        ram_buffer(31464) := X"8FC20014";
        ram_buffer(31465) := X"00000000";
        ram_buffer(31466) := X"00621021";
        ram_buffer(31467) := X"AFC20010";
        ram_buffer(31468) := X"10000002";
        ram_buffer(31469) := X"00000000";
        ram_buffer(31470) := X"AFC00014";
        ram_buffer(31471) := X"8FC30010";
        ram_buffer(31472) := X"8FC2001C";
        ram_buffer(31473) := X"00000000";
        ram_buffer(31474) := X"00621021";
        ram_buffer(31475) := X"00401821";
        ram_buffer(31476) := X"8FC20030";
        ram_buffer(31477) := X"00000000";
        ram_buffer(31478) := X"2442FFFF";
        ram_buffer(31479) := X"00621024";
        ram_buffer(31480) := X"8FC30030";
        ram_buffer(31481) := X"00000000";
        ram_buffer(31482) := X"00621023";
        ram_buffer(31483) := X"8FC30014";
        ram_buffer(31484) := X"00000000";
        ram_buffer(31485) := X"00621021";
        ram_buffer(31486) := X"AFC20014";
        ram_buffer(31487) := X"8FC20014";
        ram_buffer(31488) := X"00000000";
        ram_buffer(31489) := X"00402821";
        ram_buffer(31490) := X"8FC40048";
        ram_buffer(31491) := X"0C028390";
        ram_buffer(31492) := X"00000000";
        ram_buffer(31493) := X"AFC20018";
        ram_buffer(31494) := X"8FC30018";
        ram_buffer(31495) := X"2402FFFF";
        ram_buffer(31496) := X"14620007";
        ram_buffer(31497) := X"00000000";
        ram_buffer(31498) := X"AFC00014";
        ram_buffer(31499) := X"24020001";
        ram_buffer(31500) := X"AFC20020";
        ram_buffer(31501) := X"8FC20010";
        ram_buffer(31502) := X"00000000";
        ram_buffer(31503) := X"AFC20018";
        ram_buffer(31504) := X"3C02100D";
        ram_buffer(31505) := X"8C42D260";
        ram_buffer(31506) := X"00000000";
        ram_buffer(31507) := X"00401821";
        ram_buffer(31508) := X"8FC20014";
        ram_buffer(31509) := X"00000000";
        ram_buffer(31510) := X"00621021";
        ram_buffer(31511) := X"00401821";
        ram_buffer(31512) := X"3C02100D";
        ram_buffer(31513) := X"AC43D260";
        ram_buffer(31514) := X"3C02100D";
        ram_buffer(31515) := X"2442CBE0";
        ram_buffer(31516) := X"8FC30010";
        ram_buffer(31517) := X"00000000";
        ram_buffer(31518) := X"AC430008";
        ram_buffer(31519) := X"8FC30018";
        ram_buffer(31520) := X"8FC20010";
        ram_buffer(31521) := X"00000000";
        ram_buffer(31522) := X"00621023";
        ram_buffer(31523) := X"00401821";
        ram_buffer(31524) := X"8FC20014";
        ram_buffer(31525) := X"00000000";
        ram_buffer(31526) := X"00621021";
        ram_buffer(31527) := X"AFC20034";
        ram_buffer(31528) := X"3C02100D";
        ram_buffer(31529) := X"2442CBE0";
        ram_buffer(31530) := X"8C420008";
        ram_buffer(31531) := X"8FC30034";
        ram_buffer(31532) := X"00000000";
        ram_buffer(31533) := X"34630001";
        ram_buffer(31534) := X"AC430004";
        ram_buffer(31535) := X"3C02100D";
        ram_buffer(31536) := X"2442CBE0";
        ram_buffer(31537) := X"8FC30024";
        ram_buffer(31538) := X"00000000";
        ram_buffer(31539) := X"10620038";
        ram_buffer(31540) := X"00000000";
        ram_buffer(31541) := X"8FC20028";
        ram_buffer(31542) := X"00000000";
        ram_buffer(31543) := X"2C420010";
        ram_buffer(31544) := X"10400008";
        ram_buffer(31545) := X"00000000";
        ram_buffer(31546) := X"3C02100D";
        ram_buffer(31547) := X"2442CBE0";
        ram_buffer(31548) := X"8C420008";
        ram_buffer(31549) := X"24030001";
        ram_buffer(31550) := X"AC430004";
        ram_buffer(31551) := X"10000049";
        ram_buffer(31552) := X"00000000";
        ram_buffer(31553) := X"8FC20028";
        ram_buffer(31554) := X"00000000";
        ram_buffer(31555) := X"2443FFF4";
        ram_buffer(31556) := X"2402FFF8";
        ram_buffer(31557) := X"00621024";
        ram_buffer(31558) := X"AFC20028";
        ram_buffer(31559) := X"8FC20024";
        ram_buffer(31560) := X"00000000";
        ram_buffer(31561) := X"8C420004";
        ram_buffer(31562) := X"00000000";
        ram_buffer(31563) := X"30430001";
        ram_buffer(31564) := X"8FC20028";
        ram_buffer(31565) := X"00000000";
        ram_buffer(31566) := X"00621825";
        ram_buffer(31567) := X"8FC20024";
        ram_buffer(31568) := X"00000000";
        ram_buffer(31569) := X"AC430004";
        ram_buffer(31570) := X"8FC30024";
        ram_buffer(31571) := X"8FC20028";
        ram_buffer(31572) := X"00000000";
        ram_buffer(31573) := X"00621021";
        ram_buffer(31574) := X"24030005";
        ram_buffer(31575) := X"AC430004";
        ram_buffer(31576) := X"8FC20028";
        ram_buffer(31577) := X"00000000";
        ram_buffer(31578) := X"24420004";
        ram_buffer(31579) := X"8FC30024";
        ram_buffer(31580) := X"00000000";
        ram_buffer(31581) := X"00621021";
        ram_buffer(31582) := X"24030005";
        ram_buffer(31583) := X"AC430004";
        ram_buffer(31584) := X"8FC20028";
        ram_buffer(31585) := X"00000000";
        ram_buffer(31586) := X"2C420010";
        ram_buffer(31587) := X"14400008";
        ram_buffer(31588) := X"00000000";
        ram_buffer(31589) := X"8FC20024";
        ram_buffer(31590) := X"00000000";
        ram_buffer(31591) := X"24420008";
        ram_buffer(31592) := X"00402821";
        ram_buffer(31593) := X"8FC40048";
        ram_buffer(31594) := X"0C027301";
        ram_buffer(31595) := X"00000000";
        ram_buffer(31596) := X"3C02100D";
        ram_buffer(31597) := X"8C42D260";
        ram_buffer(31598) := X"00000000";
        ram_buffer(31599) := X"00401821";
        ram_buffer(31600) := X"8F8281B8";
        ram_buffer(31601) := X"00000000";
        ram_buffer(31602) := X"0043102B";
        ram_buffer(31603) := X"10400005";
        ram_buffer(31604) := X"00000000";
        ram_buffer(31605) := X"3C02100D";
        ram_buffer(31606) := X"8C42D260";
        ram_buffer(31607) := X"00000000";
        ram_buffer(31608) := X"AF8281B8";
        ram_buffer(31609) := X"3C02100D";
        ram_buffer(31610) := X"8C42D260";
        ram_buffer(31611) := X"00000000";
        ram_buffer(31612) := X"00401821";
        ram_buffer(31613) := X"8F8281BC";
        ram_buffer(31614) := X"00000000";
        ram_buffer(31615) := X"0043102B";
        ram_buffer(31616) := X"10400008";
        ram_buffer(31617) := X"00000000";
        ram_buffer(31618) := X"3C02100D";
        ram_buffer(31619) := X"8C42D260";
        ram_buffer(31620) := X"00000000";
        ram_buffer(31621) := X"AF8281BC";
        ram_buffer(31622) := X"10000002";
        ram_buffer(31623) := X"00000000";
        ram_buffer(31624) := X"00000000";
        ram_buffer(31625) := X"03C0E821";
        ram_buffer(31626) := X"8FBF0044";
        ram_buffer(31627) := X"8FBE0040";
        ram_buffer(31628) := X"27BD0048";
        ram_buffer(31629) := X"03E00008";
        ram_buffer(31630) := X"00000000";
        ram_buffer(31631) := X"27BDFFB0";
        ram_buffer(31632) := X"AFBF004C";
        ram_buffer(31633) := X"AFBE0048";
        ram_buffer(31634) := X"03A0F021";
        ram_buffer(31635) := X"AFC40050";
        ram_buffer(31636) := X"AFC50054";
        ram_buffer(31637) := X"8FC20054";
        ram_buffer(31638) := X"00000000";
        ram_buffer(31639) := X"2442000B";
        ram_buffer(31640) := X"2C420017";
        ram_buffer(31641) := X"14400008";
        ram_buffer(31642) := X"00000000";
        ram_buffer(31643) := X"8FC20054";
        ram_buffer(31644) := X"00000000";
        ram_buffer(31645) := X"2443000B";
        ram_buffer(31646) := X"2402FFF8";
        ram_buffer(31647) := X"00621024";
        ram_buffer(31648) := X"10000002";
        ram_buffer(31649) := X"00000000";
        ram_buffer(31650) := X"24020010";
        ram_buffer(31651) := X"AFC20034";
        ram_buffer(31652) := X"8FC20034";
        ram_buffer(31653) := X"00000000";
        ram_buffer(31654) := X"04400007";
        ram_buffer(31655) := X"00000000";
        ram_buffer(31656) := X"8FC30034";
        ram_buffer(31657) := X"8FC20054";
        ram_buffer(31658) := X"00000000";
        ram_buffer(31659) := X"0062102B";
        ram_buffer(31660) := X"10400007";
        ram_buffer(31661) := X"00000000";
        ram_buffer(31662) := X"8FC20050";
        ram_buffer(31663) := X"2403000C";
        ram_buffer(31664) := X"AC430000";
        ram_buffer(31665) := X"00001021";
        ram_buffer(31666) := X"100003DA";
        ram_buffer(31667) := X"00000000";
        ram_buffer(31668) := X"8FC40050";
        ram_buffer(31669) := X"0C0280C3";
        ram_buffer(31670) := X"00000000";
        ram_buffer(31671) := X"8FC20034";
        ram_buffer(31672) := X"00000000";
        ram_buffer(31673) := X"2C4201F8";
        ram_buffer(31674) := X"10400059";
        ram_buffer(31675) := X"00000000";
        ram_buffer(31676) := X"8FC20034";
        ram_buffer(31677) := X"00000000";
        ram_buffer(31678) := X"000210C2";
        ram_buffer(31679) := X"AFC20014";
        ram_buffer(31680) := X"8FC20014";
        ram_buffer(31681) := X"00000000";
        ram_buffer(31682) := X"24420001";
        ram_buffer(31683) := X"00021040";
        ram_buffer(31684) := X"00021880";
        ram_buffer(31685) := X"3C02100D";
        ram_buffer(31686) := X"2442CBE0";
        ram_buffer(31687) := X"00621021";
        ram_buffer(31688) := X"2442FFF8";
        ram_buffer(31689) := X"AFC20030";
        ram_buffer(31690) := X"8FC20030";
        ram_buffer(31691) := X"00000000";
        ram_buffer(31692) := X"8C42000C";
        ram_buffer(31693) := X"00000000";
        ram_buffer(31694) := X"AFC20010";
        ram_buffer(31695) := X"8FC30010";
        ram_buffer(31696) := X"8FC20030";
        ram_buffer(31697) := X"00000000";
        ram_buffer(31698) := X"1462000A";
        ram_buffer(31699) := X"00000000";
        ram_buffer(31700) := X"8FC20030";
        ram_buffer(31701) := X"00000000";
        ram_buffer(31702) := X"24420008";
        ram_buffer(31703) := X"AFC20030";
        ram_buffer(31704) := X"8FC20030";
        ram_buffer(31705) := X"00000000";
        ram_buffer(31706) := X"8C42000C";
        ram_buffer(31707) := X"00000000";
        ram_buffer(31708) := X"AFC20010";
        ram_buffer(31709) := X"8FC30010";
        ram_buffer(31710) := X"8FC20030";
        ram_buffer(31711) := X"00000000";
        ram_buffer(31712) := X"1062002D";
        ram_buffer(31713) := X"00000000";
        ram_buffer(31714) := X"8FC20010";
        ram_buffer(31715) := X"00000000";
        ram_buffer(31716) := X"8C430004";
        ram_buffer(31717) := X"2402FFFC";
        ram_buffer(31718) := X"00621024";
        ram_buffer(31719) := X"AFC20038";
        ram_buffer(31720) := X"8FC20010";
        ram_buffer(31721) := X"00000000";
        ram_buffer(31722) := X"8C42000C";
        ram_buffer(31723) := X"00000000";
        ram_buffer(31724) := X"AFC2002C";
        ram_buffer(31725) := X"8FC20010";
        ram_buffer(31726) := X"00000000";
        ram_buffer(31727) := X"8C420008";
        ram_buffer(31728) := X"00000000";
        ram_buffer(31729) := X"AFC20028";
        ram_buffer(31730) := X"8FC20028";
        ram_buffer(31731) := X"8FC3002C";
        ram_buffer(31732) := X"00000000";
        ram_buffer(31733) := X"AC43000C";
        ram_buffer(31734) := X"8FC2002C";
        ram_buffer(31735) := X"8FC30028";
        ram_buffer(31736) := X"00000000";
        ram_buffer(31737) := X"AC430008";
        ram_buffer(31738) := X"8FC30010";
        ram_buffer(31739) := X"8FC20038";
        ram_buffer(31740) := X"00000000";
        ram_buffer(31741) := X"00621021";
        ram_buffer(31742) := X"8FC40010";
        ram_buffer(31743) := X"8FC30038";
        ram_buffer(31744) := X"00000000";
        ram_buffer(31745) := X"00831821";
        ram_buffer(31746) := X"8C630004";
        ram_buffer(31747) := X"00000000";
        ram_buffer(31748) := X"34630001";
        ram_buffer(31749) := X"AC430004";
        ram_buffer(31750) := X"8FC40050";
        ram_buffer(31751) := X"0C0280CD";
        ram_buffer(31752) := X"00000000";
        ram_buffer(31753) := X"8FC20010";
        ram_buffer(31754) := X"00000000";
        ram_buffer(31755) := X"24420008";
        ram_buffer(31756) := X"10000380";
        ram_buffer(31757) := X"00000000";
        ram_buffer(31758) := X"8FC20014";
        ram_buffer(31759) := X"00000000";
        ram_buffer(31760) := X"24420002";
        ram_buffer(31761) := X"AFC20014";
        ram_buffer(31762) := X"100000A8";
        ram_buffer(31763) := X"00000000";
        ram_buffer(31764) := X"8FC20034";
        ram_buffer(31765) := X"00000000";
        ram_buffer(31766) := X"00021242";
        ram_buffer(31767) := X"14400006";
        ram_buffer(31768) := X"00000000";
        ram_buffer(31769) := X"8FC20034";
        ram_buffer(31770) := X"00000000";
        ram_buffer(31771) := X"000210C2";
        ram_buffer(31772) := X"1000003E";
        ram_buffer(31773) := X"00000000";
        ram_buffer(31774) := X"8FC20034";
        ram_buffer(31775) := X"00000000";
        ram_buffer(31776) := X"00021242";
        ram_buffer(31777) := X"2C420005";
        ram_buffer(31778) := X"10400007";
        ram_buffer(31779) := X"00000000";
        ram_buffer(31780) := X"8FC20034";
        ram_buffer(31781) := X"00000000";
        ram_buffer(31782) := X"00021182";
        ram_buffer(31783) := X"24420038";
        ram_buffer(31784) := X"10000032";
        ram_buffer(31785) := X"00000000";
        ram_buffer(31786) := X"8FC20034";
        ram_buffer(31787) := X"00000000";
        ram_buffer(31788) := X"00021242";
        ram_buffer(31789) := X"2C420015";
        ram_buffer(31790) := X"10400007";
        ram_buffer(31791) := X"00000000";
        ram_buffer(31792) := X"8FC20034";
        ram_buffer(31793) := X"00000000";
        ram_buffer(31794) := X"00021242";
        ram_buffer(31795) := X"2442005B";
        ram_buffer(31796) := X"10000026";
        ram_buffer(31797) := X"00000000";
        ram_buffer(31798) := X"8FC20034";
        ram_buffer(31799) := X"00000000";
        ram_buffer(31800) := X"00021242";
        ram_buffer(31801) := X"2C420055";
        ram_buffer(31802) := X"10400007";
        ram_buffer(31803) := X"00000000";
        ram_buffer(31804) := X"8FC20034";
        ram_buffer(31805) := X"00000000";
        ram_buffer(31806) := X"00021302";
        ram_buffer(31807) := X"2442006E";
        ram_buffer(31808) := X"1000001A";
        ram_buffer(31809) := X"00000000";
        ram_buffer(31810) := X"8FC20034";
        ram_buffer(31811) := X"00000000";
        ram_buffer(31812) := X"00021242";
        ram_buffer(31813) := X"2C420155";
        ram_buffer(31814) := X"10400007";
        ram_buffer(31815) := X"00000000";
        ram_buffer(31816) := X"8FC20034";
        ram_buffer(31817) := X"00000000";
        ram_buffer(31818) := X"000213C2";
        ram_buffer(31819) := X"24420077";
        ram_buffer(31820) := X"1000000E";
        ram_buffer(31821) := X"00000000";
        ram_buffer(31822) := X"8FC20034";
        ram_buffer(31823) := X"00000000";
        ram_buffer(31824) := X"00021242";
        ram_buffer(31825) := X"2C420555";
        ram_buffer(31826) := X"10400007";
        ram_buffer(31827) := X"00000000";
        ram_buffer(31828) := X"8FC20034";
        ram_buffer(31829) := X"00000000";
        ram_buffer(31830) := X"00021482";
        ram_buffer(31831) := X"2442007C";
        ram_buffer(31832) := X"10000002";
        ram_buffer(31833) := X"00000000";
        ram_buffer(31834) := X"2402007E";
        ram_buffer(31835) := X"AFC20014";
        ram_buffer(31836) := X"8FC20014";
        ram_buffer(31837) := X"00000000";
        ram_buffer(31838) := X"24420001";
        ram_buffer(31839) := X"00021040";
        ram_buffer(31840) := X"00021880";
        ram_buffer(31841) := X"3C02100D";
        ram_buffer(31842) := X"2442CBE0";
        ram_buffer(31843) := X"00621021";
        ram_buffer(31844) := X"2442FFF8";
        ram_buffer(31845) := X"AFC20018";
        ram_buffer(31846) := X"8FC20018";
        ram_buffer(31847) := X"00000000";
        ram_buffer(31848) := X"8C42000C";
        ram_buffer(31849) := X"00000000";
        ram_buffer(31850) := X"AFC20010";
        ram_buffer(31851) := X"10000046";
        ram_buffer(31852) := X"00000000";
        ram_buffer(31853) := X"8FC20010";
        ram_buffer(31854) := X"00000000";
        ram_buffer(31855) := X"8C430004";
        ram_buffer(31856) := X"2402FFFC";
        ram_buffer(31857) := X"00621024";
        ram_buffer(31858) := X"AFC20038";
        ram_buffer(31859) := X"8FC30038";
        ram_buffer(31860) := X"8FC20034";
        ram_buffer(31861) := X"00000000";
        ram_buffer(31862) := X"00621023";
        ram_buffer(31863) := X"AFC2001C";
        ram_buffer(31864) := X"8FC2001C";
        ram_buffer(31865) := X"00000000";
        ram_buffer(31866) := X"28420010";
        ram_buffer(31867) := X"14400007";
        ram_buffer(31868) := X"00000000";
        ram_buffer(31869) := X"8FC20014";
        ram_buffer(31870) := X"00000000";
        ram_buffer(31871) := X"2442FFFF";
        ram_buffer(31872) := X"AFC20014";
        ram_buffer(31873) := X"10000035";
        ram_buffer(31874) := X"00000000";
        ram_buffer(31875) := X"8FC2001C";
        ram_buffer(31876) := X"00000000";
        ram_buffer(31877) := X"04400027";
        ram_buffer(31878) := X"00000000";
        ram_buffer(31879) := X"8FC20010";
        ram_buffer(31880) := X"00000000";
        ram_buffer(31881) := X"8C42000C";
        ram_buffer(31882) := X"00000000";
        ram_buffer(31883) := X"AFC2002C";
        ram_buffer(31884) := X"8FC20010";
        ram_buffer(31885) := X"00000000";
        ram_buffer(31886) := X"8C420008";
        ram_buffer(31887) := X"00000000";
        ram_buffer(31888) := X"AFC20028";
        ram_buffer(31889) := X"8FC20028";
        ram_buffer(31890) := X"8FC3002C";
        ram_buffer(31891) := X"00000000";
        ram_buffer(31892) := X"AC43000C";
        ram_buffer(31893) := X"8FC2002C";
        ram_buffer(31894) := X"8FC30028";
        ram_buffer(31895) := X"00000000";
        ram_buffer(31896) := X"AC430008";
        ram_buffer(31897) := X"8FC30010";
        ram_buffer(31898) := X"8FC20038";
        ram_buffer(31899) := X"00000000";
        ram_buffer(31900) := X"00621021";
        ram_buffer(31901) := X"8FC40010";
        ram_buffer(31902) := X"8FC30038";
        ram_buffer(31903) := X"00000000";
        ram_buffer(31904) := X"00831821";
        ram_buffer(31905) := X"8C630004";
        ram_buffer(31906) := X"00000000";
        ram_buffer(31907) := X"34630001";
        ram_buffer(31908) := X"AC430004";
        ram_buffer(31909) := X"8FC40050";
        ram_buffer(31910) := X"0C0280CD";
        ram_buffer(31911) := X"00000000";
        ram_buffer(31912) := X"8FC20010";
        ram_buffer(31913) := X"00000000";
        ram_buffer(31914) := X"24420008";
        ram_buffer(31915) := X"100002E1";
        ram_buffer(31916) := X"00000000";
        ram_buffer(31917) := X"8FC20010";
        ram_buffer(31918) := X"00000000";
        ram_buffer(31919) := X"8C42000C";
        ram_buffer(31920) := X"00000000";
        ram_buffer(31921) := X"AFC20010";
        ram_buffer(31922) := X"8FC30010";
        ram_buffer(31923) := X"8FC20018";
        ram_buffer(31924) := X"00000000";
        ram_buffer(31925) := X"1462FFB7";
        ram_buffer(31926) := X"00000000";
        ram_buffer(31927) := X"8FC20014";
        ram_buffer(31928) := X"00000000";
        ram_buffer(31929) := X"24420001";
        ram_buffer(31930) := X"AFC20014";
        ram_buffer(31931) := X"3C02100D";
        ram_buffer(31932) := X"2442CBE8";
        ram_buffer(31933) := X"8C420008";
        ram_buffer(31934) := X"00000000";
        ram_buffer(31935) := X"AFC20010";
        ram_buffer(31936) := X"3C02100D";
        ram_buffer(31937) := X"2442CBE8";
        ram_buffer(31938) := X"8FC30010";
        ram_buffer(31939) := X"00000000";
        ram_buffer(31940) := X"1062013E";
        ram_buffer(31941) := X"00000000";
        ram_buffer(31942) := X"8FC20010";
        ram_buffer(31943) := X"00000000";
        ram_buffer(31944) := X"8C430004";
        ram_buffer(31945) := X"2402FFFC";
        ram_buffer(31946) := X"00621024";
        ram_buffer(31947) := X"AFC20038";
        ram_buffer(31948) := X"8FC30038";
        ram_buffer(31949) := X"8FC20034";
        ram_buffer(31950) := X"00000000";
        ram_buffer(31951) := X"00621023";
        ram_buffer(31952) := X"AFC2001C";
        ram_buffer(31953) := X"8FC2001C";
        ram_buffer(31954) := X"00000000";
        ram_buffer(31955) := X"28420010";
        ram_buffer(31956) := X"14400037";
        ram_buffer(31957) := X"00000000";
        ram_buffer(31958) := X"8FC30010";
        ram_buffer(31959) := X"8FC20034";
        ram_buffer(31960) := X"00000000";
        ram_buffer(31961) := X"00621021";
        ram_buffer(31962) := X"AFC2003C";
        ram_buffer(31963) := X"8FC20034";
        ram_buffer(31964) := X"00000000";
        ram_buffer(31965) := X"34430001";
        ram_buffer(31966) := X"8FC20010";
        ram_buffer(31967) := X"00000000";
        ram_buffer(31968) := X"AC430004";
        ram_buffer(31969) := X"3C02100D";
        ram_buffer(31970) := X"2443CBE8";
        ram_buffer(31971) := X"3C02100D";
        ram_buffer(31972) := X"2442CBE8";
        ram_buffer(31973) := X"8FC4003C";
        ram_buffer(31974) := X"00000000";
        ram_buffer(31975) := X"AC44000C";
        ram_buffer(31976) := X"8C42000C";
        ram_buffer(31977) := X"00000000";
        ram_buffer(31978) := X"AC620008";
        ram_buffer(31979) := X"3C02100D";
        ram_buffer(31980) := X"2443CBE8";
        ram_buffer(31981) := X"8FC2003C";
        ram_buffer(31982) := X"00000000";
        ram_buffer(31983) := X"AC43000C";
        ram_buffer(31984) := X"8FC2003C";
        ram_buffer(31985) := X"00000000";
        ram_buffer(31986) := X"8C43000C";
        ram_buffer(31987) := X"8FC2003C";
        ram_buffer(31988) := X"00000000";
        ram_buffer(31989) := X"AC430008";
        ram_buffer(31990) := X"8FC2001C";
        ram_buffer(31991) := X"00000000";
        ram_buffer(31992) := X"34420001";
        ram_buffer(31993) := X"00401821";
        ram_buffer(31994) := X"8FC2003C";
        ram_buffer(31995) := X"00000000";
        ram_buffer(31996) := X"AC430004";
        ram_buffer(31997) := X"8FC2001C";
        ram_buffer(31998) := X"8FC3003C";
        ram_buffer(31999) := X"00000000";
        ram_buffer(32000) := X"00621021";
        ram_buffer(32001) := X"8FC3001C";
        ram_buffer(32002) := X"00000000";
        ram_buffer(32003) := X"AC430000";
        ram_buffer(32004) := X"8FC40050";
        ram_buffer(32005) := X"0C0280CD";
        ram_buffer(32006) := X"00000000";
        ram_buffer(32007) := X"8FC20010";
        ram_buffer(32008) := X"00000000";
        ram_buffer(32009) := X"24420008";
        ram_buffer(32010) := X"10000282";
        ram_buffer(32011) := X"00000000";
        ram_buffer(32012) := X"3C02100D";
        ram_buffer(32013) := X"2443CBE8";
        ram_buffer(32014) := X"3C02100D";
        ram_buffer(32015) := X"2442CBE8";
        ram_buffer(32016) := X"3C04100D";
        ram_buffer(32017) := X"2484CBE8";
        ram_buffer(32018) := X"AC44000C";
        ram_buffer(32019) := X"8C42000C";
        ram_buffer(32020) := X"00000000";
        ram_buffer(32021) := X"AC620008";
        ram_buffer(32022) := X"8FC2001C";
        ram_buffer(32023) := X"00000000";
        ram_buffer(32024) := X"04400015";
        ram_buffer(32025) := X"00000000";
        ram_buffer(32026) := X"8FC30010";
        ram_buffer(32027) := X"8FC20038";
        ram_buffer(32028) := X"00000000";
        ram_buffer(32029) := X"00621021";
        ram_buffer(32030) := X"8FC40010";
        ram_buffer(32031) := X"8FC30038";
        ram_buffer(32032) := X"00000000";
        ram_buffer(32033) := X"00831821";
        ram_buffer(32034) := X"8C630004";
        ram_buffer(32035) := X"00000000";
        ram_buffer(32036) := X"34630001";
        ram_buffer(32037) := X"AC430004";
        ram_buffer(32038) := X"8FC40050";
        ram_buffer(32039) := X"0C0280CD";
        ram_buffer(32040) := X"00000000";
        ram_buffer(32041) := X"8FC20010";
        ram_buffer(32042) := X"00000000";
        ram_buffer(32043) := X"24420008";
        ram_buffer(32044) := X"10000260";
        ram_buffer(32045) := X"00000000";
        ram_buffer(32046) := X"8FC20038";
        ram_buffer(32047) := X"00000000";
        ram_buffer(32048) := X"2C420200";
        ram_buffer(32049) := X"10400038";
        ram_buffer(32050) := X"00000000";
        ram_buffer(32051) := X"8FC20038";
        ram_buffer(32052) := X"00000000";
        ram_buffer(32053) := X"000210C2";
        ram_buffer(32054) := X"AFC20040";
        ram_buffer(32055) := X"3C02100D";
        ram_buffer(32056) := X"2443CBE0";
        ram_buffer(32057) := X"3C02100D";
        ram_buffer(32058) := X"2442CBE0";
        ram_buffer(32059) := X"8C440004";
        ram_buffer(32060) := X"8FC20040";
        ram_buffer(32061) := X"00000000";
        ram_buffer(32062) := X"04410002";
        ram_buffer(32063) := X"00000000";
        ram_buffer(32064) := X"24420003";
        ram_buffer(32065) := X"00021083";
        ram_buffer(32066) := X"00402821";
        ram_buffer(32067) := X"24020001";
        ram_buffer(32068) := X"00A21004";
        ram_buffer(32069) := X"00821025";
        ram_buffer(32070) := X"AC620004";
        ram_buffer(32071) := X"8FC20040";
        ram_buffer(32072) := X"00000000";
        ram_buffer(32073) := X"24420001";
        ram_buffer(32074) := X"00021040";
        ram_buffer(32075) := X"00021880";
        ram_buffer(32076) := X"3C02100D";
        ram_buffer(32077) := X"2442CBE0";
        ram_buffer(32078) := X"00621021";
        ram_buffer(32079) := X"2442FFF8";
        ram_buffer(32080) := X"AFC2002C";
        ram_buffer(32081) := X"8FC2002C";
        ram_buffer(32082) := X"00000000";
        ram_buffer(32083) := X"8C420008";
        ram_buffer(32084) := X"00000000";
        ram_buffer(32085) := X"AFC20028";
        ram_buffer(32086) := X"8FC20010";
        ram_buffer(32087) := X"8FC3002C";
        ram_buffer(32088) := X"00000000";
        ram_buffer(32089) := X"AC43000C";
        ram_buffer(32090) := X"8FC20010";
        ram_buffer(32091) := X"8FC30028";
        ram_buffer(32092) := X"00000000";
        ram_buffer(32093) := X"AC430008";
        ram_buffer(32094) := X"8FC2002C";
        ram_buffer(32095) := X"8FC30010";
        ram_buffer(32096) := X"00000000";
        ram_buffer(32097) := X"AC430008";
        ram_buffer(32098) := X"8FC2002C";
        ram_buffer(32099) := X"00000000";
        ram_buffer(32100) := X"8C430008";
        ram_buffer(32101) := X"8FC20028";
        ram_buffer(32102) := X"00000000";
        ram_buffer(32103) := X"AC43000C";
        ram_buffer(32104) := X"1000009A";
        ram_buffer(32105) := X"00000000";
        ram_buffer(32106) := X"8FC20038";
        ram_buffer(32107) := X"00000000";
        ram_buffer(32108) := X"00021242";
        ram_buffer(32109) := X"14400006";
        ram_buffer(32110) := X"00000000";
        ram_buffer(32111) := X"8FC20038";
        ram_buffer(32112) := X"00000000";
        ram_buffer(32113) := X"000210C2";
        ram_buffer(32114) := X"1000003E";
        ram_buffer(32115) := X"00000000";
        ram_buffer(32116) := X"8FC20038";
        ram_buffer(32117) := X"00000000";
        ram_buffer(32118) := X"00021242";
        ram_buffer(32119) := X"2C420005";
        ram_buffer(32120) := X"10400007";
        ram_buffer(32121) := X"00000000";
        ram_buffer(32122) := X"8FC20038";
        ram_buffer(32123) := X"00000000";
        ram_buffer(32124) := X"00021182";
        ram_buffer(32125) := X"24420038";
        ram_buffer(32126) := X"10000032";
        ram_buffer(32127) := X"00000000";
        ram_buffer(32128) := X"8FC20038";
        ram_buffer(32129) := X"00000000";
        ram_buffer(32130) := X"00021242";
        ram_buffer(32131) := X"2C420015";
        ram_buffer(32132) := X"10400007";
        ram_buffer(32133) := X"00000000";
        ram_buffer(32134) := X"8FC20038";
        ram_buffer(32135) := X"00000000";
        ram_buffer(32136) := X"00021242";
        ram_buffer(32137) := X"2442005B";
        ram_buffer(32138) := X"10000026";
        ram_buffer(32139) := X"00000000";
        ram_buffer(32140) := X"8FC20038";
        ram_buffer(32141) := X"00000000";
        ram_buffer(32142) := X"00021242";
        ram_buffer(32143) := X"2C420055";
        ram_buffer(32144) := X"10400007";
        ram_buffer(32145) := X"00000000";
        ram_buffer(32146) := X"8FC20038";
        ram_buffer(32147) := X"00000000";
        ram_buffer(32148) := X"00021302";
        ram_buffer(32149) := X"2442006E";
        ram_buffer(32150) := X"1000001A";
        ram_buffer(32151) := X"00000000";
        ram_buffer(32152) := X"8FC20038";
        ram_buffer(32153) := X"00000000";
        ram_buffer(32154) := X"00021242";
        ram_buffer(32155) := X"2C420155";
        ram_buffer(32156) := X"10400007";
        ram_buffer(32157) := X"00000000";
        ram_buffer(32158) := X"8FC20038";
        ram_buffer(32159) := X"00000000";
        ram_buffer(32160) := X"000213C2";
        ram_buffer(32161) := X"24420077";
        ram_buffer(32162) := X"1000000E";
        ram_buffer(32163) := X"00000000";
        ram_buffer(32164) := X"8FC20038";
        ram_buffer(32165) := X"00000000";
        ram_buffer(32166) := X"00021242";
        ram_buffer(32167) := X"2C420555";
        ram_buffer(32168) := X"10400007";
        ram_buffer(32169) := X"00000000";
        ram_buffer(32170) := X"8FC20038";
        ram_buffer(32171) := X"00000000";
        ram_buffer(32172) := X"00021482";
        ram_buffer(32173) := X"2442007C";
        ram_buffer(32174) := X"10000002";
        ram_buffer(32175) := X"00000000";
        ram_buffer(32176) := X"2402007E";
        ram_buffer(32177) := X"AFC20040";
        ram_buffer(32178) := X"8FC20040";
        ram_buffer(32179) := X"00000000";
        ram_buffer(32180) := X"24420001";
        ram_buffer(32181) := X"00021040";
        ram_buffer(32182) := X"00021880";
        ram_buffer(32183) := X"3C02100D";
        ram_buffer(32184) := X"2442CBE0";
        ram_buffer(32185) := X"00621021";
        ram_buffer(32186) := X"2442FFF8";
        ram_buffer(32187) := X"AFC2002C";
        ram_buffer(32188) := X"8FC2002C";
        ram_buffer(32189) := X"00000000";
        ram_buffer(32190) := X"8C420008";
        ram_buffer(32191) := X"00000000";
        ram_buffer(32192) := X"AFC20028";
        ram_buffer(32193) := X"8FC30028";
        ram_buffer(32194) := X"8FC2002C";
        ram_buffer(32195) := X"00000000";
        ram_buffer(32196) := X"14620018";
        ram_buffer(32197) := X"00000000";
        ram_buffer(32198) := X"3C02100D";
        ram_buffer(32199) := X"2443CBE0";
        ram_buffer(32200) := X"3C02100D";
        ram_buffer(32201) := X"2442CBE0";
        ram_buffer(32202) := X"8C440004";
        ram_buffer(32203) := X"8FC20040";
        ram_buffer(32204) := X"00000000";
        ram_buffer(32205) := X"04410002";
        ram_buffer(32206) := X"00000000";
        ram_buffer(32207) := X"24420003";
        ram_buffer(32208) := X"00021083";
        ram_buffer(32209) := X"00402821";
        ram_buffer(32210) := X"24020001";
        ram_buffer(32211) := X"00A21004";
        ram_buffer(32212) := X"00821025";
        ram_buffer(32213) := X"AC620004";
        ram_buffer(32214) := X"1000001A";
        ram_buffer(32215) := X"00000000";
        ram_buffer(32216) := X"8FC20028";
        ram_buffer(32217) := X"00000000";
        ram_buffer(32218) := X"8C420008";
        ram_buffer(32219) := X"00000000";
        ram_buffer(32220) := X"AFC20028";
        ram_buffer(32221) := X"8FC30028";
        ram_buffer(32222) := X"8FC2002C";
        ram_buffer(32223) := X"00000000";
        ram_buffer(32224) := X"1062000B";
        ram_buffer(32225) := X"00000000";
        ram_buffer(32226) := X"8FC20028";
        ram_buffer(32227) := X"00000000";
        ram_buffer(32228) := X"8C430004";
        ram_buffer(32229) := X"2402FFFC";
        ram_buffer(32230) := X"00621824";
        ram_buffer(32231) := X"8FC20038";
        ram_buffer(32232) := X"00000000";
        ram_buffer(32233) := X"0043102B";
        ram_buffer(32234) := X"1440FFED";
        ram_buffer(32235) := X"00000000";
        ram_buffer(32236) := X"8FC20028";
        ram_buffer(32237) := X"00000000";
        ram_buffer(32238) := X"8C42000C";
        ram_buffer(32239) := X"00000000";
        ram_buffer(32240) := X"AFC2002C";
        ram_buffer(32241) := X"8FC20010";
        ram_buffer(32242) := X"8FC3002C";
        ram_buffer(32243) := X"00000000";
        ram_buffer(32244) := X"AC43000C";
        ram_buffer(32245) := X"8FC20010";
        ram_buffer(32246) := X"8FC30028";
        ram_buffer(32247) := X"00000000";
        ram_buffer(32248) := X"AC430008";
        ram_buffer(32249) := X"8FC2002C";
        ram_buffer(32250) := X"8FC30010";
        ram_buffer(32251) := X"00000000";
        ram_buffer(32252) := X"AC430008";
        ram_buffer(32253) := X"8FC2002C";
        ram_buffer(32254) := X"00000000";
        ram_buffer(32255) := X"8C430008";
        ram_buffer(32256) := X"8FC20028";
        ram_buffer(32257) := X"00000000";
        ram_buffer(32258) := X"AC43000C";
        ram_buffer(32259) := X"8FC20014";
        ram_buffer(32260) := X"00000000";
        ram_buffer(32261) := X"04410002";
        ram_buffer(32262) := X"00000000";
        ram_buffer(32263) := X"24420003";
        ram_buffer(32264) := X"00021083";
        ram_buffer(32265) := X"00401821";
        ram_buffer(32266) := X"24020001";
        ram_buffer(32267) := X"00621004";
        ram_buffer(32268) := X"AFC20020";
        ram_buffer(32269) := X"3C02100D";
        ram_buffer(32270) := X"2442CBE0";
        ram_buffer(32271) := X"8C420004";
        ram_buffer(32272) := X"8FC30020";
        ram_buffer(32273) := X"00000000";
        ram_buffer(32274) := X"0043102B";
        ram_buffer(32275) := X"14400118";
        ram_buffer(32276) := X"00000000";
        ram_buffer(32277) := X"3C02100D";
        ram_buffer(32278) := X"2442CBE0";
        ram_buffer(32279) := X"8C430004";
        ram_buffer(32280) := X"8FC20020";
        ram_buffer(32281) := X"00000000";
        ram_buffer(32282) := X"00621024";
        ram_buffer(32283) := X"1440001C";
        ram_buffer(32284) := X"00000000";
        ram_buffer(32285) := X"8FC30014";
        ram_buffer(32286) := X"2402FFFC";
        ram_buffer(32287) := X"00621024";
        ram_buffer(32288) := X"24420004";
        ram_buffer(32289) := X"AFC20014";
        ram_buffer(32290) := X"8FC20020";
        ram_buffer(32291) := X"00000000";
        ram_buffer(32292) := X"00021040";
        ram_buffer(32293) := X"AFC20020";
        ram_buffer(32294) := X"10000009";
        ram_buffer(32295) := X"00000000";
        ram_buffer(32296) := X"8FC20014";
        ram_buffer(32297) := X"00000000";
        ram_buffer(32298) := X"24420004";
        ram_buffer(32299) := X"AFC20014";
        ram_buffer(32300) := X"8FC20020";
        ram_buffer(32301) := X"00000000";
        ram_buffer(32302) := X"00021040";
        ram_buffer(32303) := X"AFC20020";
        ram_buffer(32304) := X"3C02100D";
        ram_buffer(32305) := X"2442CBE0";
        ram_buffer(32306) := X"8C430004";
        ram_buffer(32307) := X"8FC20020";
        ram_buffer(32308) := X"00000000";
        ram_buffer(32309) := X"00621024";
        ram_buffer(32310) := X"1040FFF1";
        ram_buffer(32311) := X"00000000";
        ram_buffer(32312) := X"8FC20014";
        ram_buffer(32313) := X"00000000";
        ram_buffer(32314) := X"AFC20024";
        ram_buffer(32315) := X"8FC20014";
        ram_buffer(32316) := X"00000000";
        ram_buffer(32317) := X"24420001";
        ram_buffer(32318) := X"00021040";
        ram_buffer(32319) := X"00021880";
        ram_buffer(32320) := X"3C02100D";
        ram_buffer(32321) := X"2442CBE0";
        ram_buffer(32322) := X"00621021";
        ram_buffer(32323) := X"2442FFF8";
        ram_buffer(32324) := X"AFC20018";
        ram_buffer(32325) := X"8FC20018";
        ram_buffer(32326) := X"00000000";
        ram_buffer(32327) := X"AFC20030";
        ram_buffer(32328) := X"8FC20018";
        ram_buffer(32329) := X"00000000";
        ram_buffer(32330) := X"8C42000C";
        ram_buffer(32331) := X"00000000";
        ram_buffer(32332) := X"AFC20010";
        ram_buffer(32333) := X"10000088";
        ram_buffer(32334) := X"00000000";
        ram_buffer(32335) := X"8FC20010";
        ram_buffer(32336) := X"00000000";
        ram_buffer(32337) := X"8C430004";
        ram_buffer(32338) := X"2402FFFC";
        ram_buffer(32339) := X"00621024";
        ram_buffer(32340) := X"AFC20038";
        ram_buffer(32341) := X"8FC30038";
        ram_buffer(32342) := X"8FC20034";
        ram_buffer(32343) := X"00000000";
        ram_buffer(32344) := X"00621023";
        ram_buffer(32345) := X"AFC2001C";
        ram_buffer(32346) := X"8FC2001C";
        ram_buffer(32347) := X"00000000";
        ram_buffer(32348) := X"28420010";
        ram_buffer(32349) := X"14400049";
        ram_buffer(32350) := X"00000000";
        ram_buffer(32351) := X"8FC30010";
        ram_buffer(32352) := X"8FC20034";
        ram_buffer(32353) := X"00000000";
        ram_buffer(32354) := X"00621021";
        ram_buffer(32355) := X"AFC2003C";
        ram_buffer(32356) := X"8FC20034";
        ram_buffer(32357) := X"00000000";
        ram_buffer(32358) := X"34430001";
        ram_buffer(32359) := X"8FC20010";
        ram_buffer(32360) := X"00000000";
        ram_buffer(32361) := X"AC430004";
        ram_buffer(32362) := X"8FC20010";
        ram_buffer(32363) := X"00000000";
        ram_buffer(32364) := X"8C42000C";
        ram_buffer(32365) := X"00000000";
        ram_buffer(32366) := X"AFC2002C";
        ram_buffer(32367) := X"8FC20010";
        ram_buffer(32368) := X"00000000";
        ram_buffer(32369) := X"8C420008";
        ram_buffer(32370) := X"00000000";
        ram_buffer(32371) := X"AFC20028";
        ram_buffer(32372) := X"8FC20028";
        ram_buffer(32373) := X"8FC3002C";
        ram_buffer(32374) := X"00000000";
        ram_buffer(32375) := X"AC43000C";
        ram_buffer(32376) := X"8FC2002C";
        ram_buffer(32377) := X"8FC30028";
        ram_buffer(32378) := X"00000000";
        ram_buffer(32379) := X"AC430008";
        ram_buffer(32380) := X"3C02100D";
        ram_buffer(32381) := X"2443CBE8";
        ram_buffer(32382) := X"3C02100D";
        ram_buffer(32383) := X"2442CBE8";
        ram_buffer(32384) := X"8FC4003C";
        ram_buffer(32385) := X"00000000";
        ram_buffer(32386) := X"AC44000C";
        ram_buffer(32387) := X"8C42000C";
        ram_buffer(32388) := X"00000000";
        ram_buffer(32389) := X"AC620008";
        ram_buffer(32390) := X"3C02100D";
        ram_buffer(32391) := X"2443CBE8";
        ram_buffer(32392) := X"8FC2003C";
        ram_buffer(32393) := X"00000000";
        ram_buffer(32394) := X"AC43000C";
        ram_buffer(32395) := X"8FC2003C";
        ram_buffer(32396) := X"00000000";
        ram_buffer(32397) := X"8C43000C";
        ram_buffer(32398) := X"8FC2003C";
        ram_buffer(32399) := X"00000000";
        ram_buffer(32400) := X"AC430008";
        ram_buffer(32401) := X"8FC2001C";
        ram_buffer(32402) := X"00000000";
        ram_buffer(32403) := X"34420001";
        ram_buffer(32404) := X"00401821";
        ram_buffer(32405) := X"8FC2003C";
        ram_buffer(32406) := X"00000000";
        ram_buffer(32407) := X"AC430004";
        ram_buffer(32408) := X"8FC2001C";
        ram_buffer(32409) := X"8FC3003C";
        ram_buffer(32410) := X"00000000";
        ram_buffer(32411) := X"00621021";
        ram_buffer(32412) := X"8FC3001C";
        ram_buffer(32413) := X"00000000";
        ram_buffer(32414) := X"AC430000";
        ram_buffer(32415) := X"8FC40050";
        ram_buffer(32416) := X"0C0280CD";
        ram_buffer(32417) := X"00000000";
        ram_buffer(32418) := X"8FC20010";
        ram_buffer(32419) := X"00000000";
        ram_buffer(32420) := X"24420008";
        ram_buffer(32421) := X"100000E7";
        ram_buffer(32422) := X"00000000";
        ram_buffer(32423) := X"8FC2001C";
        ram_buffer(32424) := X"00000000";
        ram_buffer(32425) := X"04400027";
        ram_buffer(32426) := X"00000000";
        ram_buffer(32427) := X"8FC30010";
        ram_buffer(32428) := X"8FC20038";
        ram_buffer(32429) := X"00000000";
        ram_buffer(32430) := X"00621021";
        ram_buffer(32431) := X"8FC40010";
        ram_buffer(32432) := X"8FC30038";
        ram_buffer(32433) := X"00000000";
        ram_buffer(32434) := X"00831821";
        ram_buffer(32435) := X"8C630004";
        ram_buffer(32436) := X"00000000";
        ram_buffer(32437) := X"34630001";
        ram_buffer(32438) := X"AC430004";
        ram_buffer(32439) := X"8FC20010";
        ram_buffer(32440) := X"00000000";
        ram_buffer(32441) := X"8C42000C";
        ram_buffer(32442) := X"00000000";
        ram_buffer(32443) := X"AFC2002C";
        ram_buffer(32444) := X"8FC20010";
        ram_buffer(32445) := X"00000000";
        ram_buffer(32446) := X"8C420008";
        ram_buffer(32447) := X"00000000";
        ram_buffer(32448) := X"AFC20028";
        ram_buffer(32449) := X"8FC20028";
        ram_buffer(32450) := X"8FC3002C";
        ram_buffer(32451) := X"00000000";
        ram_buffer(32452) := X"AC43000C";
        ram_buffer(32453) := X"8FC2002C";
        ram_buffer(32454) := X"8FC30028";
        ram_buffer(32455) := X"00000000";
        ram_buffer(32456) := X"AC430008";
        ram_buffer(32457) := X"8FC40050";
        ram_buffer(32458) := X"0C0280CD";
        ram_buffer(32459) := X"00000000";
        ram_buffer(32460) := X"8FC20010";
        ram_buffer(32461) := X"00000000";
        ram_buffer(32462) := X"24420008";
        ram_buffer(32463) := X"100000BD";
        ram_buffer(32464) := X"00000000";
        ram_buffer(32465) := X"8FC20010";
        ram_buffer(32466) := X"00000000";
        ram_buffer(32467) := X"8C42000C";
        ram_buffer(32468) := X"00000000";
        ram_buffer(32469) := X"AFC20010";
        ram_buffer(32470) := X"8FC30010";
        ram_buffer(32471) := X"8FC20018";
        ram_buffer(32472) := X"00000000";
        ram_buffer(32473) := X"1462FF75";
        ram_buffer(32474) := X"00000000";
        ram_buffer(32475) := X"8FC20018";
        ram_buffer(32476) := X"00000000";
        ram_buffer(32477) := X"24420008";
        ram_buffer(32478) := X"AFC20018";
        ram_buffer(32479) := X"8FC20014";
        ram_buffer(32480) := X"00000000";
        ram_buffer(32481) := X"24420001";
        ram_buffer(32482) := X"AFC20014";
        ram_buffer(32483) := X"8FC20014";
        ram_buffer(32484) := X"00000000";
        ram_buffer(32485) := X"30420003";
        ram_buffer(32486) := X"1440FF61";
        ram_buffer(32487) := X"00000000";
        ram_buffer(32488) := X"8FC20024";
        ram_buffer(32489) := X"00000000";
        ram_buffer(32490) := X"30420003";
        ram_buffer(32491) := X"1440000D";
        ram_buffer(32492) := X"00000000";
        ram_buffer(32493) := X"3C02100D";
        ram_buffer(32494) := X"2442CBE0";
        ram_buffer(32495) := X"3C03100D";
        ram_buffer(32496) := X"2463CBE0";
        ram_buffer(32497) := X"8C640004";
        ram_buffer(32498) := X"8FC30020";
        ram_buffer(32499) := X"00000000";
        ram_buffer(32500) := X"00031827";
        ram_buffer(32501) := X"00831824";
        ram_buffer(32502) := X"AC430004";
        ram_buffer(32503) := X"10000010";
        ram_buffer(32504) := X"00000000";
        ram_buffer(32505) := X"8FC20024";
        ram_buffer(32506) := X"00000000";
        ram_buffer(32507) := X"2442FFFF";
        ram_buffer(32508) := X"AFC20024";
        ram_buffer(32509) := X"8FC20030";
        ram_buffer(32510) := X"00000000";
        ram_buffer(32511) := X"2442FFF8";
        ram_buffer(32512) := X"AFC20030";
        ram_buffer(32513) := X"8FC20030";
        ram_buffer(32514) := X"00000000";
        ram_buffer(32515) := X"8C430008";
        ram_buffer(32516) := X"8FC20030";
        ram_buffer(32517) := X"00000000";
        ram_buffer(32518) := X"1062FFE1";
        ram_buffer(32519) := X"00000000";
        ram_buffer(32520) := X"8FC20020";
        ram_buffer(32521) := X"00000000";
        ram_buffer(32522) := X"00021040";
        ram_buffer(32523) := X"AFC20020";
        ram_buffer(32524) := X"3C02100D";
        ram_buffer(32525) := X"2442CBE0";
        ram_buffer(32526) := X"8C420004";
        ram_buffer(32527) := X"8FC30020";
        ram_buffer(32528) := X"00000000";
        ram_buffer(32529) := X"0043102B";
        ram_buffer(32530) := X"14400019";
        ram_buffer(32531) := X"00000000";
        ram_buffer(32532) := X"8FC20020";
        ram_buffer(32533) := X"00000000";
        ram_buffer(32534) := X"10400015";
        ram_buffer(32535) := X"00000000";
        ram_buffer(32536) := X"10000009";
        ram_buffer(32537) := X"00000000";
        ram_buffer(32538) := X"8FC20014";
        ram_buffer(32539) := X"00000000";
        ram_buffer(32540) := X"24420004";
        ram_buffer(32541) := X"AFC20014";
        ram_buffer(32542) := X"8FC20020";
        ram_buffer(32543) := X"00000000";
        ram_buffer(32544) := X"00021040";
        ram_buffer(32545) := X"AFC20020";
        ram_buffer(32546) := X"3C02100D";
        ram_buffer(32547) := X"2442CBE0";
        ram_buffer(32548) := X"8C430004";
        ram_buffer(32549) := X"8FC20020";
        ram_buffer(32550) := X"00000000";
        ram_buffer(32551) := X"00621024";
        ram_buffer(32552) := X"1040FFF1";
        ram_buffer(32553) := X"00000000";
        ram_buffer(32554) := X"1000FF0D";
        ram_buffer(32555) := X"00000000";
        ram_buffer(32556) := X"3C02100D";
        ram_buffer(32557) := X"2442CBE0";
        ram_buffer(32558) := X"8C420008";
        ram_buffer(32559) := X"00000000";
        ram_buffer(32560) := X"8C430004";
        ram_buffer(32561) := X"2402FFFC";
        ram_buffer(32562) := X"00621824";
        ram_buffer(32563) := X"8FC20034";
        ram_buffer(32564) := X"00000000";
        ram_buffer(32565) := X"00621023";
        ram_buffer(32566) := X"AFC2001C";
        ram_buffer(32567) := X"3C02100D";
        ram_buffer(32568) := X"2442CBE0";
        ram_buffer(32569) := X"8C420008";
        ram_buffer(32570) := X"00000000";
        ram_buffer(32571) := X"8C430004";
        ram_buffer(32572) := X"2402FFFC";
        ram_buffer(32573) := X"00621824";
        ram_buffer(32574) := X"8FC20034";
        ram_buffer(32575) := X"00000000";
        ram_buffer(32576) := X"0062102B";
        ram_buffer(32577) := X"14400006";
        ram_buffer(32578) := X"00000000";
        ram_buffer(32579) := X"8FC2001C";
        ram_buffer(32580) := X"00000000";
        ram_buffer(32581) := X"28420010";
        ram_buffer(32582) := X"10400027";
        ram_buffer(32583) := X"00000000";
        ram_buffer(32584) := X"8FC50034";
        ram_buffer(32585) := X"8FC40050";
        ram_buffer(32586) := X"0C027A5E";
        ram_buffer(32587) := X"00000000";
        ram_buffer(32588) := X"3C02100D";
        ram_buffer(32589) := X"2442CBE0";
        ram_buffer(32590) := X"8C420008";
        ram_buffer(32591) := X"00000000";
        ram_buffer(32592) := X"8C430004";
        ram_buffer(32593) := X"2402FFFC";
        ram_buffer(32594) := X"00621824";
        ram_buffer(32595) := X"8FC20034";
        ram_buffer(32596) := X"00000000";
        ram_buffer(32597) := X"00621023";
        ram_buffer(32598) := X"AFC2001C";
        ram_buffer(32599) := X"3C02100D";
        ram_buffer(32600) := X"2442CBE0";
        ram_buffer(32601) := X"8C420008";
        ram_buffer(32602) := X"00000000";
        ram_buffer(32603) := X"8C430004";
        ram_buffer(32604) := X"2402FFFC";
        ram_buffer(32605) := X"00621824";
        ram_buffer(32606) := X"8FC20034";
        ram_buffer(32607) := X"00000000";
        ram_buffer(32608) := X"0062102B";
        ram_buffer(32609) := X"14400006";
        ram_buffer(32610) := X"00000000";
        ram_buffer(32611) := X"8FC2001C";
        ram_buffer(32612) := X"00000000";
        ram_buffer(32613) := X"28420010";
        ram_buffer(32614) := X"10400007";
        ram_buffer(32615) := X"00000000";
        ram_buffer(32616) := X"8FC40050";
        ram_buffer(32617) := X"0C0280CD";
        ram_buffer(32618) := X"00000000";
        ram_buffer(32619) := X"00001021";
        ram_buffer(32620) := X"10000020";
        ram_buffer(32621) := X"00000000";
        ram_buffer(32622) := X"3C02100D";
        ram_buffer(32623) := X"2442CBE0";
        ram_buffer(32624) := X"8C420008";
        ram_buffer(32625) := X"00000000";
        ram_buffer(32626) := X"AFC20010";
        ram_buffer(32627) := X"8FC20034";
        ram_buffer(32628) := X"00000000";
        ram_buffer(32629) := X"34430001";
        ram_buffer(32630) := X"8FC20010";
        ram_buffer(32631) := X"00000000";
        ram_buffer(32632) := X"AC430004";
        ram_buffer(32633) := X"3C02100D";
        ram_buffer(32634) := X"2442CBE0";
        ram_buffer(32635) := X"8FC40010";
        ram_buffer(32636) := X"8FC30034";
        ram_buffer(32637) := X"00000000";
        ram_buffer(32638) := X"00831821";
        ram_buffer(32639) := X"AC430008";
        ram_buffer(32640) := X"3C02100D";
        ram_buffer(32641) := X"2442CBE0";
        ram_buffer(32642) := X"8C420008";
        ram_buffer(32643) := X"8FC3001C";
        ram_buffer(32644) := X"00000000";
        ram_buffer(32645) := X"34630001";
        ram_buffer(32646) := X"AC430004";
        ram_buffer(32647) := X"8FC40050";
        ram_buffer(32648) := X"0C0280CD";
        ram_buffer(32649) := X"00000000";
        ram_buffer(32650) := X"8FC20010";
        ram_buffer(32651) := X"00000000";
        ram_buffer(32652) := X"24420008";
        ram_buffer(32653) := X"03C0E821";
        ram_buffer(32654) := X"8FBF004C";
        ram_buffer(32655) := X"8FBE0048";
        ram_buffer(32656) := X"27BD0050";
        ram_buffer(32657) := X"03E00008";
        ram_buffer(32658) := X"00000000";
        ram_buffer(32659) := X"27BDFFE8";
        ram_buffer(32660) := X"AFBE0014";
        ram_buffer(32661) := X"03A0F021";
        ram_buffer(32662) := X"AFC40018";
        ram_buffer(32663) := X"AFC5001C";
        ram_buffer(32664) := X"AFC60020";
        ram_buffer(32665) := X"8FC20018";
        ram_buffer(32666) := X"00000000";
        ram_buffer(32667) := X"AFC20000";
        ram_buffer(32668) := X"8FC2001C";
        ram_buffer(32669) := X"00000000";
        ram_buffer(32670) := X"AFC20004";
        ram_buffer(32671) := X"8FC20020";
        ram_buffer(32672) := X"00000000";
        ram_buffer(32673) := X"2C420010";
        ram_buffer(32674) := X"1440006E";
        ram_buffer(32675) := X"00000000";
        ram_buffer(32676) := X"8FC30004";
        ram_buffer(32677) := X"8FC20000";
        ram_buffer(32678) := X"00000000";
        ram_buffer(32679) := X"00621025";
        ram_buffer(32680) := X"30420003";
        ram_buffer(32681) := X"14400067";
        ram_buffer(32682) := X"00000000";
        ram_buffer(32683) := X"8FC20000";
        ram_buffer(32684) := X"00000000";
        ram_buffer(32685) := X"AFC20008";
        ram_buffer(32686) := X"8FC20004";
        ram_buffer(32687) := X"00000000";
        ram_buffer(32688) := X"AFC2000C";
        ram_buffer(32689) := X"10000031";
        ram_buffer(32690) := X"00000000";
        ram_buffer(32691) := X"8FC20008";
        ram_buffer(32692) := X"00000000";
        ram_buffer(32693) := X"24430004";
        ram_buffer(32694) := X"AFC30008";
        ram_buffer(32695) := X"8FC3000C";
        ram_buffer(32696) := X"00000000";
        ram_buffer(32697) := X"24640004";
        ram_buffer(32698) := X"AFC4000C";
        ram_buffer(32699) := X"8C630000";
        ram_buffer(32700) := X"00000000";
        ram_buffer(32701) := X"AC430000";
        ram_buffer(32702) := X"8FC20008";
        ram_buffer(32703) := X"00000000";
        ram_buffer(32704) := X"24430004";
        ram_buffer(32705) := X"AFC30008";
        ram_buffer(32706) := X"8FC3000C";
        ram_buffer(32707) := X"00000000";
        ram_buffer(32708) := X"24640004";
        ram_buffer(32709) := X"AFC4000C";
        ram_buffer(32710) := X"8C630000";
        ram_buffer(32711) := X"00000000";
        ram_buffer(32712) := X"AC430000";
        ram_buffer(32713) := X"8FC20008";
        ram_buffer(32714) := X"00000000";
        ram_buffer(32715) := X"24430004";
        ram_buffer(32716) := X"AFC30008";
        ram_buffer(32717) := X"8FC3000C";
        ram_buffer(32718) := X"00000000";
        ram_buffer(32719) := X"24640004";
        ram_buffer(32720) := X"AFC4000C";
        ram_buffer(32721) := X"8C630000";
        ram_buffer(32722) := X"00000000";
        ram_buffer(32723) := X"AC430000";
        ram_buffer(32724) := X"8FC20008";
        ram_buffer(32725) := X"00000000";
        ram_buffer(32726) := X"24430004";
        ram_buffer(32727) := X"AFC30008";
        ram_buffer(32728) := X"8FC3000C";
        ram_buffer(32729) := X"00000000";
        ram_buffer(32730) := X"24640004";
        ram_buffer(32731) := X"AFC4000C";
        ram_buffer(32732) := X"8C630000";
        ram_buffer(32733) := X"00000000";
        ram_buffer(32734) := X"AC430000";
        ram_buffer(32735) := X"8FC20020";
        ram_buffer(32736) := X"00000000";
        ram_buffer(32737) := X"2442FFF0";
        ram_buffer(32738) := X"AFC20020";
        ram_buffer(32739) := X"8FC20020";
        ram_buffer(32740) := X"00000000";
        ram_buffer(32741) := X"2C420010";
        ram_buffer(32742) := X"1040FFCC";
        ram_buffer(32743) := X"00000000";
        ram_buffer(32744) := X"10000010";
        ram_buffer(32745) := X"00000000";
        ram_buffer(32746) := X"8FC20008";
        ram_buffer(32747) := X"00000000";
        ram_buffer(32748) := X"24430004";
        ram_buffer(32749) := X"AFC30008";
        ram_buffer(32750) := X"8FC3000C";
        ram_buffer(32751) := X"00000000";
        ram_buffer(32752) := X"24640004";
        ram_buffer(32753) := X"AFC4000C";
        ram_buffer(32754) := X"8C630000";
        ram_buffer(32755) := X"00000000";
        ram_buffer(32756) := X"AC430000";
        ram_buffer(32757) := X"8FC20020";
        ram_buffer(32758) := X"00000000";
        ram_buffer(32759) := X"2442FFFC";
        ram_buffer(32760) := X"AFC20020";
        ram_buffer(32761) := X"8FC20020";
        ram_buffer(32762) := X"00000000";
        ram_buffer(32763) := X"2C420004";
        ram_buffer(32764) := X"1040FFED";
        ram_buffer(32765) := X"00000000";
        ram_buffer(32766) := X"8FC20008";
        ram_buffer(32767) := X"00000000";
        ram_buffer(32768) := X"AFC20000";
        ram_buffer(32769) := X"8FC2000C";
        ram_buffer(32770) := X"00000000";
        ram_buffer(32771) := X"AFC20004";
        ram_buffer(32772) := X"1000000C";
        ram_buffer(32773) := X"00000000";
        ram_buffer(32774) := X"8FC20000";
        ram_buffer(32775) := X"00000000";
        ram_buffer(32776) := X"24430001";
        ram_buffer(32777) := X"AFC30000";
        ram_buffer(32778) := X"8FC30004";
        ram_buffer(32779) := X"00000000";
        ram_buffer(32780) := X"24640001";
        ram_buffer(32781) := X"AFC40004";
        ram_buffer(32782) := X"80630000";
        ram_buffer(32783) := X"00000000";
        ram_buffer(32784) := X"A0430000";
        ram_buffer(32785) := X"8FC20020";
        ram_buffer(32786) := X"00000000";
        ram_buffer(32787) := X"2443FFFF";
        ram_buffer(32788) := X"AFC30020";
        ram_buffer(32789) := X"1440FFF0";
        ram_buffer(32790) := X"00000000";
        ram_buffer(32791) := X"8FC20018";
        ram_buffer(32792) := X"03C0E821";
        ram_buffer(32793) := X"8FBE0014";
        ram_buffer(32794) := X"27BD0018";
        ram_buffer(32795) := X"03E00008";
        ram_buffer(32796) := X"00000000";
        ram_buffer(32797) := X"27BDFFE0";
        ram_buffer(32798) := X"AFBE001C";
        ram_buffer(32799) := X"03A0F021";
        ram_buffer(32800) := X"AFC40020";
        ram_buffer(32801) := X"AFC50024";
        ram_buffer(32802) := X"AFC60028";
        ram_buffer(32803) := X"8FC20020";
        ram_buffer(32804) := X"00000000";
        ram_buffer(32805) := X"AFC20000";
        ram_buffer(32806) := X"8FC20024";
        ram_buffer(32807) := X"00000000";
        ram_buffer(32808) := X"304200FF";
        ram_buffer(32809) := X"AFC20010";
        ram_buffer(32810) := X"10000015";
        ram_buffer(32811) := X"00000000";
        ram_buffer(32812) := X"8FC20028";
        ram_buffer(32813) := X"00000000";
        ram_buffer(32814) := X"2443FFFF";
        ram_buffer(32815) := X"AFC30028";
        ram_buffer(32816) := X"1040000C";
        ram_buffer(32817) := X"00000000";
        ram_buffer(32818) := X"8FC20000";
        ram_buffer(32819) := X"00000000";
        ram_buffer(32820) := X"24430001";
        ram_buffer(32821) := X"AFC30000";
        ram_buffer(32822) := X"8FC30024";
        ram_buffer(32823) := X"00000000";
        ram_buffer(32824) := X"00031E00";
        ram_buffer(32825) := X"00031E03";
        ram_buffer(32826) := X"A0430000";
        ram_buffer(32827) := X"10000004";
        ram_buffer(32828) := X"00000000";
        ram_buffer(32829) := X"8FC20020";
        ram_buffer(32830) := X"1000007F";
        ram_buffer(32831) := X"00000000";
        ram_buffer(32832) := X"8FC20000";
        ram_buffer(32833) := X"00000000";
        ram_buffer(32834) := X"30420003";
        ram_buffer(32835) := X"1440FFE8";
        ram_buffer(32836) := X"00000000";
        ram_buffer(32837) := X"8FC20028";
        ram_buffer(32838) := X"00000000";
        ram_buffer(32839) := X"2C420004";
        ram_buffer(32840) := X"1440006E";
        ram_buffer(32841) := X"00000000";
        ram_buffer(32842) := X"8FC20000";
        ram_buffer(32843) := X"00000000";
        ram_buffer(32844) := X"AFC2000C";
        ram_buffer(32845) := X"8FC20010";
        ram_buffer(32846) := X"00000000";
        ram_buffer(32847) := X"00021A00";
        ram_buffer(32848) := X"8FC20010";
        ram_buffer(32849) := X"00000000";
        ram_buffer(32850) := X"00621025";
        ram_buffer(32851) := X"AFC20008";
        ram_buffer(32852) := X"8FC20008";
        ram_buffer(32853) := X"00000000";
        ram_buffer(32854) := X"00021400";
        ram_buffer(32855) := X"8FC30008";
        ram_buffer(32856) := X"00000000";
        ram_buffer(32857) := X"00621025";
        ram_buffer(32858) := X"AFC20008";
        ram_buffer(32859) := X"24020020";
        ram_buffer(32860) := X"AFC20004";
        ram_buffer(32861) := X"1000000D";
        ram_buffer(32862) := X"00000000";
        ram_buffer(32863) := X"8FC30008";
        ram_buffer(32864) := X"8FC20004";
        ram_buffer(32865) := X"00000000";
        ram_buffer(32866) := X"00431004";
        ram_buffer(32867) := X"8FC30008";
        ram_buffer(32868) := X"00000000";
        ram_buffer(32869) := X"00621025";
        ram_buffer(32870) := X"AFC20008";
        ram_buffer(32871) := X"8FC20004";
        ram_buffer(32872) := X"00000000";
        ram_buffer(32873) := X"00021040";
        ram_buffer(32874) := X"AFC20004";
        ram_buffer(32875) := X"8FC20004";
        ram_buffer(32876) := X"00000000";
        ram_buffer(32877) := X"2C420020";
        ram_buffer(32878) := X"1440FFF0";
        ram_buffer(32879) := X"00000000";
        ram_buffer(32880) := X"10000021";
        ram_buffer(32881) := X"00000000";
        ram_buffer(32882) := X"8FC2000C";
        ram_buffer(32883) := X"00000000";
        ram_buffer(32884) := X"24430004";
        ram_buffer(32885) := X"AFC3000C";
        ram_buffer(32886) := X"8FC30008";
        ram_buffer(32887) := X"00000000";
        ram_buffer(32888) := X"AC430000";
        ram_buffer(32889) := X"8FC2000C";
        ram_buffer(32890) := X"00000000";
        ram_buffer(32891) := X"24430004";
        ram_buffer(32892) := X"AFC3000C";
        ram_buffer(32893) := X"8FC30008";
        ram_buffer(32894) := X"00000000";
        ram_buffer(32895) := X"AC430000";
        ram_buffer(32896) := X"8FC2000C";
        ram_buffer(32897) := X"00000000";
        ram_buffer(32898) := X"24430004";
        ram_buffer(32899) := X"AFC3000C";
        ram_buffer(32900) := X"8FC30008";
        ram_buffer(32901) := X"00000000";
        ram_buffer(32902) := X"AC430000";
        ram_buffer(32903) := X"8FC2000C";
        ram_buffer(32904) := X"00000000";
        ram_buffer(32905) := X"24430004";
        ram_buffer(32906) := X"AFC3000C";
        ram_buffer(32907) := X"8FC30008";
        ram_buffer(32908) := X"00000000";
        ram_buffer(32909) := X"AC430000";
        ram_buffer(32910) := X"8FC20028";
        ram_buffer(32911) := X"00000000";
        ram_buffer(32912) := X"2442FFF0";
        ram_buffer(32913) := X"AFC20028";
        ram_buffer(32914) := X"8FC20028";
        ram_buffer(32915) := X"00000000";
        ram_buffer(32916) := X"2C420010";
        ram_buffer(32917) := X"1040FFDC";
        ram_buffer(32918) := X"00000000";
        ram_buffer(32919) := X"1000000C";
        ram_buffer(32920) := X"00000000";
        ram_buffer(32921) := X"8FC2000C";
        ram_buffer(32922) := X"00000000";
        ram_buffer(32923) := X"24430004";
        ram_buffer(32924) := X"AFC3000C";
        ram_buffer(32925) := X"8FC30008";
        ram_buffer(32926) := X"00000000";
        ram_buffer(32927) := X"AC430000";
        ram_buffer(32928) := X"8FC20028";
        ram_buffer(32929) := X"00000000";
        ram_buffer(32930) := X"2442FFFC";
        ram_buffer(32931) := X"AFC20028";
        ram_buffer(32932) := X"8FC20028";
        ram_buffer(32933) := X"00000000";
        ram_buffer(32934) := X"2C420004";
        ram_buffer(32935) := X"1040FFF1";
        ram_buffer(32936) := X"00000000";
        ram_buffer(32937) := X"8FC2000C";
        ram_buffer(32938) := X"00000000";
        ram_buffer(32939) := X"AFC20000";
        ram_buffer(32940) := X"1000000A";
        ram_buffer(32941) := X"00000000";
        ram_buffer(32942) := X"8FC20000";
        ram_buffer(32943) := X"00000000";
        ram_buffer(32944) := X"24430001";
        ram_buffer(32945) := X"AFC30000";
        ram_buffer(32946) := X"8FC30024";
        ram_buffer(32947) := X"00000000";
        ram_buffer(32948) := X"00031E00";
        ram_buffer(32949) := X"00031E03";
        ram_buffer(32950) := X"A0430000";
        ram_buffer(32951) := X"8FC20028";
        ram_buffer(32952) := X"00000000";
        ram_buffer(32953) := X"2443FFFF";
        ram_buffer(32954) := X"AFC30028";
        ram_buffer(32955) := X"1440FFF2";
        ram_buffer(32956) := X"00000000";
        ram_buffer(32957) := X"8FC20020";
        ram_buffer(32958) := X"03C0E821";
        ram_buffer(32959) := X"8FBE001C";
        ram_buffer(32960) := X"27BD0020";
        ram_buffer(32961) := X"03E00008";
        ram_buffer(32962) := X"00000000";
        ram_buffer(32963) := X"27BDFFF8";
        ram_buffer(32964) := X"AFBE0004";
        ram_buffer(32965) := X"03A0F021";
        ram_buffer(32966) := X"AFC40008";
        ram_buffer(32967) := X"00000000";
        ram_buffer(32968) := X"03C0E821";
        ram_buffer(32969) := X"8FBE0004";
        ram_buffer(32970) := X"27BD0008";
        ram_buffer(32971) := X"03E00008";
        ram_buffer(32972) := X"00000000";
        ram_buffer(32973) := X"27BDFFF8";
        ram_buffer(32974) := X"AFBE0004";
        ram_buffer(32975) := X"03A0F021";
        ram_buffer(32976) := X"AFC40008";
        ram_buffer(32977) := X"00000000";
        ram_buffer(32978) := X"03C0E821";
        ram_buffer(32979) := X"8FBE0004";
        ram_buffer(32980) := X"27BD0008";
        ram_buffer(32981) := X"03E00008";
        ram_buffer(32982) := X"00000000";
        ram_buffer(32983) := X"27BDFFE0";
        ram_buffer(32984) := X"AFBF001C";
        ram_buffer(32985) := X"AFBE0018";
        ram_buffer(32986) := X"03A0F021";
        ram_buffer(32987) := X"AFC40020";
        ram_buffer(32988) := X"AFC50024";
        ram_buffer(32989) := X"AFC60028";
        ram_buffer(32990) := X"AFC7002C";
        ram_buffer(32991) := X"AF8081EC";
        ram_buffer(32992) := X"8FC6002C";
        ram_buffer(32993) := X"8FC50028";
        ram_buffer(32994) := X"8FC40024";
        ram_buffer(32995) := X"0C02FBF6";
        ram_buffer(32996) := X"00000000";
        ram_buffer(32997) := X"AFC20010";
        ram_buffer(32998) := X"8FC30010";
        ram_buffer(32999) := X"2402FFFF";
        ram_buffer(33000) := X"14620009";
        ram_buffer(33001) := X"00000000";
        ram_buffer(33002) := X"8F8281EC";
        ram_buffer(33003) := X"00000000";
        ram_buffer(33004) := X"10400005";
        ram_buffer(33005) := X"00000000";
        ram_buffer(33006) := X"8F8381EC";
        ram_buffer(33007) := X"8FC20020";
        ram_buffer(33008) := X"00000000";
        ram_buffer(33009) := X"AC430000";
        ram_buffer(33010) := X"8FC20010";
        ram_buffer(33011) := X"03C0E821";
        ram_buffer(33012) := X"8FBF001C";
        ram_buffer(33013) := X"8FBE0018";
        ram_buffer(33014) := X"27BD0020";
        ram_buffer(33015) := X"03E00008";
        ram_buffer(33016) := X"00000000";
        ram_buffer(33017) := X"27BDFFE0";
        ram_buffer(33018) := X"AFBF001C";
        ram_buffer(33019) := X"AFBE0018";
        ram_buffer(33020) := X"03A0F021";
        ram_buffer(33021) := X"AFC40020";
        ram_buffer(33022) := X"AFC50024";
        ram_buffer(33023) := X"AFC60028";
        ram_buffer(33024) := X"AFC7002C";
        ram_buffer(33025) := X"27C20028";
        ram_buffer(33026) := X"AFC20014";
        ram_buffer(33027) := X"8FC20020";
        ram_buffer(33028) := X"00000000";
        ram_buffer(33029) := X"8C420008";
        ram_buffer(33030) := X"8FC30014";
        ram_buffer(33031) := X"00000000";
        ram_buffer(33032) := X"00603821";
        ram_buffer(33033) := X"8FC60024";
        ram_buffer(33034) := X"00402821";
        ram_buffer(33035) := X"8FC40020";
        ram_buffer(33036) := X"0C029DFA";
        ram_buffer(33037) := X"00000000";
        ram_buffer(33038) := X"AFC20010";
        ram_buffer(33039) := X"8FC20010";
        ram_buffer(33040) := X"03C0E821";
        ram_buffer(33041) := X"8FBF001C";
        ram_buffer(33042) := X"8FBE0018";
        ram_buffer(33043) := X"27BD0020";
        ram_buffer(33044) := X"03E00008";
        ram_buffer(33045) := X"00000000";
        ram_buffer(33046) := X"27BDFFD8";
        ram_buffer(33047) := X"AFBF0024";
        ram_buffer(33048) := X"AFBE0020";
        ram_buffer(33049) := X"03A0F021";
        ram_buffer(33050) := X"AFC40028";
        ram_buffer(33051) := X"AFC5002C";
        ram_buffer(33052) := X"AFC60030";
        ram_buffer(33053) := X"AFC70034";
        ram_buffer(33054) := X"8F828098";
        ram_buffer(33055) := X"00000000";
        ram_buffer(33056) := X"AFC20010";
        ram_buffer(33057) := X"27C2002C";
        ram_buffer(33058) := X"AFC20018";
        ram_buffer(33059) := X"8FC20010";
        ram_buffer(33060) := X"00000000";
        ram_buffer(33061) := X"8C420008";
        ram_buffer(33062) := X"8FC30018";
        ram_buffer(33063) := X"00000000";
        ram_buffer(33064) := X"00603821";
        ram_buffer(33065) := X"8FC60028";
        ram_buffer(33066) := X"00402821";
        ram_buffer(33067) := X"8FC40010";
        ram_buffer(33068) := X"0C029DFA";
        ram_buffer(33069) := X"00000000";
        ram_buffer(33070) := X"AFC20014";
        ram_buffer(33071) := X"8FC20014";
        ram_buffer(33072) := X"03C0E821";
        ram_buffer(33073) := X"8FBF0024";
        ram_buffer(33074) := X"8FBE0020";
        ram_buffer(33075) := X"27BD0028";
        ram_buffer(33076) := X"03E00008";
        ram_buffer(33077) := X"00000000";
        ram_buffer(33078) := X"27BDFFC0";
        ram_buffer(33079) := X"AFBF003C";
        ram_buffer(33080) := X"AFBE0038";
        ram_buffer(33081) := X"03A0F021";
        ram_buffer(33082) := X"AFC40040";
        ram_buffer(33083) := X"AFC50044";
        ram_buffer(33084) := X"8FC40044";
        ram_buffer(33085) := X"0C02851E";
        ram_buffer(33086) := X"00000000";
        ram_buffer(33087) := X"AFC20010";
        ram_buffer(33088) := X"8FC20044";
        ram_buffer(33089) := X"00000000";
        ram_buffer(33090) := X"AFC20028";
        ram_buffer(33091) := X"8FC20010";
        ram_buffer(33092) := X"00000000";
        ram_buffer(33093) := X"AFC2002C";
        ram_buffer(33094) := X"3C02100D";
        ram_buffer(33095) := X"2442A074";
        ram_buffer(33096) := X"AFC20030";
        ram_buffer(33097) := X"24020001";
        ram_buffer(33098) := X"AFC20034";
        ram_buffer(33099) := X"8FC20010";
        ram_buffer(33100) := X"00000000";
        ram_buffer(33101) := X"24420001";
        ram_buffer(33102) := X"AFC20024";
        ram_buffer(33103) := X"27C20028";
        ram_buffer(33104) := X"AFC2001C";
        ram_buffer(33105) := X"24020002";
        ram_buffer(33106) := X"AFC20020";
        ram_buffer(33107) := X"8FC20040";
        ram_buffer(33108) := X"00000000";
        ram_buffer(33109) := X"8C420008";
        ram_buffer(33110) := X"00000000";
        ram_buffer(33111) := X"AFC20014";
        ram_buffer(33112) := X"8FC20014";
        ram_buffer(33113) := X"00000000";
        ram_buffer(33114) := X"8442000C";
        ram_buffer(33115) := X"00000000";
        ram_buffer(33116) := X"3042FFFF";
        ram_buffer(33117) := X"30422000";
        ram_buffer(33118) := X"14400013";
        ram_buffer(33119) := X"00000000";
        ram_buffer(33120) := X"8FC20014";
        ram_buffer(33121) := X"00000000";
        ram_buffer(33122) := X"8442000C";
        ram_buffer(33123) := X"00000000";
        ram_buffer(33124) := X"34422000";
        ram_buffer(33125) := X"00021C00";
        ram_buffer(33126) := X"00031C03";
        ram_buffer(33127) := X"8FC20014";
        ram_buffer(33128) := X"00000000";
        ram_buffer(33129) := X"A443000C";
        ram_buffer(33130) := X"8FC20014";
        ram_buffer(33131) := X"00000000";
        ram_buffer(33132) := X"8C430064";
        ram_buffer(33133) := X"2402DFFF";
        ram_buffer(33134) := X"00621824";
        ram_buffer(33135) := X"8FC20014";
        ram_buffer(33136) := X"00000000";
        ram_buffer(33137) := X"AC430064";
        ram_buffer(33138) := X"27C2001C";
        ram_buffer(33139) := X"00403021";
        ram_buffer(33140) := X"8FC50014";
        ram_buffer(33141) := X"8FC40040";
        ram_buffer(33142) := X"0C02B89A";
        ram_buffer(33143) := X"00000000";
        ram_buffer(33144) := X"10400004";
        ram_buffer(33145) := X"00000000";
        ram_buffer(33146) := X"2402FFFF";
        ram_buffer(33147) := X"10000002";
        ram_buffer(33148) := X"00000000";
        ram_buffer(33149) := X"2402000A";
        ram_buffer(33150) := X"AFC20018";
        ram_buffer(33151) := X"8FC20018";
        ram_buffer(33152) := X"03C0E821";
        ram_buffer(33153) := X"8FBF003C";
        ram_buffer(33154) := X"8FBE0038";
        ram_buffer(33155) := X"27BD0040";
        ram_buffer(33156) := X"03E00008";
        ram_buffer(33157) := X"00000000";
        ram_buffer(33158) := X"27BDFFE8";
        ram_buffer(33159) := X"AFBF0014";
        ram_buffer(33160) := X"AFBE0010";
        ram_buffer(33161) := X"03A0F021";
        ram_buffer(33162) := X"AFC40018";
        ram_buffer(33163) := X"8F828098";
        ram_buffer(33164) := X"8FC50018";
        ram_buffer(33165) := X"00402021";
        ram_buffer(33166) := X"0C028136";
        ram_buffer(33167) := X"00000000";
        ram_buffer(33168) := X"03C0E821";
        ram_buffer(33169) := X"8FBF0014";
        ram_buffer(33170) := X"8FBE0010";
        ram_buffer(33171) := X"27BD0018";
        ram_buffer(33172) := X"03E00008";
        ram_buffer(33173) := X"00000000";
        ram_buffer(33174) := X"27BDFFE8";
        ram_buffer(33175) := X"AFBF0014";
        ram_buffer(33176) := X"AFBE0010";
        ram_buffer(33177) := X"03A0F021";
        ram_buffer(33178) := X"AFC40018";
        ram_buffer(33179) := X"AFC5001C";
        ram_buffer(33180) := X"8FC2001C";
        ram_buffer(33181) := X"00000000";
        ram_buffer(33182) := X"8C420000";
        ram_buffer(33183) := X"00000000";
        ram_buffer(33184) := X"10400009";
        ram_buffer(33185) := X"00000000";
        ram_buffer(33186) := X"8FC2001C";
        ram_buffer(33187) := X"00000000";
        ram_buffer(33188) := X"8C420000";
        ram_buffer(33189) := X"00000000";
        ram_buffer(33190) := X"00402821";
        ram_buffer(33191) := X"8FC40018";
        ram_buffer(33192) := X"0C028196";
        ram_buffer(33193) := X"00000000";
        ram_buffer(33194) := X"8FC5001C";
        ram_buffer(33195) := X"8FC40018";
        ram_buffer(33196) := X"0C027301";
        ram_buffer(33197) := X"00000000";
        ram_buffer(33198) := X"00000000";
        ram_buffer(33199) := X"03C0E821";
        ram_buffer(33200) := X"8FBF0014";
        ram_buffer(33201) := X"8FBE0010";
        ram_buffer(33202) := X"27BD0018";
        ram_buffer(33203) := X"03E00008";
        ram_buffer(33204) := X"00000000";
        ram_buffer(33205) := X"27BDFFD0";
        ram_buffer(33206) := X"AFBF002C";
        ram_buffer(33207) := X"AFBE0028";
        ram_buffer(33208) := X"03A0F021";
        ram_buffer(33209) := X"AFC40030";
        ram_buffer(33210) := X"8F828098";
        ram_buffer(33211) := X"8FC30030";
        ram_buffer(33212) := X"00000000";
        ram_buffer(33213) := X"10620095";
        ram_buffer(33214) := X"00000000";
        ram_buffer(33215) := X"8FC20030";
        ram_buffer(33216) := X"00000000";
        ram_buffer(33217) := X"8C42004C";
        ram_buffer(33218) := X"00000000";
        ram_buffer(33219) := X"10400031";
        ram_buffer(33220) := X"00000000";
        ram_buffer(33221) := X"AFC00010";
        ram_buffer(33222) := X"10000021";
        ram_buffer(33223) := X"00000000";
        ram_buffer(33224) := X"8FC20030";
        ram_buffer(33225) := X"00000000";
        ram_buffer(33226) := X"8C43004C";
        ram_buffer(33227) := X"8FC20010";
        ram_buffer(33228) := X"00000000";
        ram_buffer(33229) := X"00021080";
        ram_buffer(33230) := X"00621021";
        ram_buffer(33231) := X"8C420000";
        ram_buffer(33232) := X"00000000";
        ram_buffer(33233) := X"AFC20014";
        ram_buffer(33234) := X"1000000D";
        ram_buffer(33235) := X"00000000";
        ram_buffer(33236) := X"8FC20014";
        ram_buffer(33237) := X"00000000";
        ram_buffer(33238) := X"AFC2001C";
        ram_buffer(33239) := X"8FC20014";
        ram_buffer(33240) := X"00000000";
        ram_buffer(33241) := X"8C420000";
        ram_buffer(33242) := X"00000000";
        ram_buffer(33243) := X"AFC20014";
        ram_buffer(33244) := X"8FC5001C";
        ram_buffer(33245) := X"8FC40030";
        ram_buffer(33246) := X"0C027301";
        ram_buffer(33247) := X"00000000";
        ram_buffer(33248) := X"8FC20014";
        ram_buffer(33249) := X"00000000";
        ram_buffer(33250) := X"1440FFF1";
        ram_buffer(33251) := X"00000000";
        ram_buffer(33252) := X"8FC20010";
        ram_buffer(33253) := X"00000000";
        ram_buffer(33254) := X"24420001";
        ram_buffer(33255) := X"AFC20010";
        ram_buffer(33256) := X"8FC20010";
        ram_buffer(33257) := X"00000000";
        ram_buffer(33258) := X"2C420020";
        ram_buffer(33259) := X"1440FFDC";
        ram_buffer(33260) := X"00000000";
        ram_buffer(33261) := X"8FC20030";
        ram_buffer(33262) := X"00000000";
        ram_buffer(33263) := X"8C42004C";
        ram_buffer(33264) := X"00000000";
        ram_buffer(33265) := X"00402821";
        ram_buffer(33266) := X"8FC40030";
        ram_buffer(33267) := X"0C027301";
        ram_buffer(33268) := X"00000000";
        ram_buffer(33269) := X"8FC20030";
        ram_buffer(33270) := X"00000000";
        ram_buffer(33271) := X"8C420040";
        ram_buffer(33272) := X"00000000";
        ram_buffer(33273) := X"10400009";
        ram_buffer(33274) := X"00000000";
        ram_buffer(33275) := X"8FC20030";
        ram_buffer(33276) := X"00000000";
        ram_buffer(33277) := X"8C420040";
        ram_buffer(33278) := X"00000000";
        ram_buffer(33279) := X"00402821";
        ram_buffer(33280) := X"8FC40030";
        ram_buffer(33281) := X"0C027301";
        ram_buffer(33282) := X"00000000";
        ram_buffer(33283) := X"8FC20030";
        ram_buffer(33284) := X"00000000";
        ram_buffer(33285) := X"8C420148";
        ram_buffer(33286) := X"00000000";
        ram_buffer(33287) := X"10400023";
        ram_buffer(33288) := X"00000000";
        ram_buffer(33289) := X"8FC20030";
        ram_buffer(33290) := X"00000000";
        ram_buffer(33291) := X"8C430148";
        ram_buffer(33292) := X"8FC20030";
        ram_buffer(33293) := X"00000000";
        ram_buffer(33294) := X"2442014C";
        ram_buffer(33295) := X"1062001B";
        ram_buffer(33296) := X"00000000";
        ram_buffer(33297) := X"8FC20030";
        ram_buffer(33298) := X"00000000";
        ram_buffer(33299) := X"8C420148";
        ram_buffer(33300) := X"00000000";
        ram_buffer(33301) := X"AFC20018";
        ram_buffer(33302) := X"1000000D";
        ram_buffer(33303) := X"00000000";
        ram_buffer(33304) := X"8FC20018";
        ram_buffer(33305) := X"00000000";
        ram_buffer(33306) := X"AFC20020";
        ram_buffer(33307) := X"8FC20018";
        ram_buffer(33308) := X"00000000";
        ram_buffer(33309) := X"8C420000";
        ram_buffer(33310) := X"00000000";
        ram_buffer(33311) := X"AFC20018";
        ram_buffer(33312) := X"8FC50020";
        ram_buffer(33313) := X"8FC40030";
        ram_buffer(33314) := X"0C027301";
        ram_buffer(33315) := X"00000000";
        ram_buffer(33316) := X"8FC20030";
        ram_buffer(33317) := X"00000000";
        ram_buffer(33318) := X"2443014C";
        ram_buffer(33319) := X"8FC20018";
        ram_buffer(33320) := X"00000000";
        ram_buffer(33321) := X"1462FFEE";
        ram_buffer(33322) := X"00000000";
        ram_buffer(33323) := X"8FC20030";
        ram_buffer(33324) := X"00000000";
        ram_buffer(33325) := X"8C420054";
        ram_buffer(33326) := X"00000000";
        ram_buffer(33327) := X"10400009";
        ram_buffer(33328) := X"00000000";
        ram_buffer(33329) := X"8FC20030";
        ram_buffer(33330) := X"00000000";
        ram_buffer(33331) := X"8C420054";
        ram_buffer(33332) := X"00000000";
        ram_buffer(33333) := X"00402821";
        ram_buffer(33334) := X"8FC40030";
        ram_buffer(33335) := X"0C027301";
        ram_buffer(33336) := X"00000000";
        ram_buffer(33337) := X"8FC20030";
        ram_buffer(33338) := X"00000000";
        ram_buffer(33339) := X"8C420038";
        ram_buffer(33340) := X"00000000";
        ram_buffer(33341) := X"10400015";
        ram_buffer(33342) := X"00000000";
        ram_buffer(33343) := X"8FC20030";
        ram_buffer(33344) := X"00000000";
        ram_buffer(33345) := X"8C42003C";
        ram_buffer(33346) := X"8FC40030";
        ram_buffer(33347) := X"0040F809";
        ram_buffer(33348) := X"00000000";
        ram_buffer(33349) := X"8FC20030";
        ram_buffer(33350) := X"00000000";
        ram_buffer(33351) := X"8C4202E0";
        ram_buffer(33352) := X"00000000";
        ram_buffer(33353) := X"10400009";
        ram_buffer(33354) := X"00000000";
        ram_buffer(33355) := X"8FC20030";
        ram_buffer(33356) := X"00000000";
        ram_buffer(33357) := X"8C4202E0";
        ram_buffer(33358) := X"00000000";
        ram_buffer(33359) := X"00402821";
        ram_buffer(33360) := X"8FC40030";
        ram_buffer(33361) := X"0C028196";
        ram_buffer(33362) := X"00000000";
        ram_buffer(33363) := X"00000000";
        ram_buffer(33364) := X"03C0E821";
        ram_buffer(33365) := X"8FBF002C";
        ram_buffer(33366) := X"8FBE0028";
        ram_buffer(33367) := X"27BD0030";
        ram_buffer(33368) := X"03E00008";
        ram_buffer(33369) := X"00000000";
        ram_buffer(33370) := X"27BDFFE8";
        ram_buffer(33371) := X"AFBF0014";
        ram_buffer(33372) := X"AFBE0010";
        ram_buffer(33373) := X"03A0F021";
        ram_buffer(33374) := X"AFC40018";
        ram_buffer(33375) := X"8FC20018";
        ram_buffer(33376) := X"00000000";
        ram_buffer(33377) := X"8442000C";
        ram_buffer(33378) := X"00000000";
        ram_buffer(33379) := X"3042FFFF";
        ram_buffer(33380) := X"30430009";
        ram_buffer(33381) := X"24020009";
        ram_buffer(33382) := X"14620006";
        ram_buffer(33383) := X"00000000";
        ram_buffer(33384) := X"8FC40018";
        ram_buffer(33385) := X"0C026F0C";
        ram_buffer(33386) := X"00000000";
        ram_buffer(33387) := X"10000002";
        ram_buffer(33388) := X"00000000";
        ram_buffer(33389) := X"00001021";
        ram_buffer(33390) := X"03C0E821";
        ram_buffer(33391) := X"8FBF0014";
        ram_buffer(33392) := X"8FBE0010";
        ram_buffer(33393) := X"27BD0018";
        ram_buffer(33394) := X"03E00008";
        ram_buffer(33395) := X"00000000";
        ram_buffer(33396) := X"27BDFFD8";
        ram_buffer(33397) := X"AFBF0024";
        ram_buffer(33398) := X"AFBE0020";
        ram_buffer(33399) := X"AFB0001C";
        ram_buffer(33400) := X"03A0F021";
        ram_buffer(33401) := X"AFC40028";
        ram_buffer(33402) := X"00A08021";
        ram_buffer(33403) := X"8FC20028";
        ram_buffer(33404) := X"00000000";
        ram_buffer(33405) := X"AFC20010";
        ram_buffer(33406) := X"8FC20010";
        ram_buffer(33407) := X"00000000";
        ram_buffer(33408) := X"1040000A";
        ram_buffer(33409) := X"00000000";
        ram_buffer(33410) := X"8FC20010";
        ram_buffer(33411) := X"00000000";
        ram_buffer(33412) := X"8C420038";
        ram_buffer(33413) := X"00000000";
        ram_buffer(33414) := X"14400004";
        ram_buffer(33415) := X"00000000";
        ram_buffer(33416) := X"8FC40010";
        ram_buffer(33417) := X"0C027069";
        ram_buffer(33418) := X"00000000";
        ram_buffer(33419) := X"8602000C";
        ram_buffer(33420) := X"00000000";
        ram_buffer(33421) := X"3042FFFF";
        ram_buffer(33422) := X"30422000";
        ram_buffer(33423) := X"1440000B";
        ram_buffer(33424) := X"00000000";
        ram_buffer(33425) := X"8602000C";
        ram_buffer(33426) := X"00000000";
        ram_buffer(33427) := X"34422000";
        ram_buffer(33428) := X"00021400";
        ram_buffer(33429) := X"00021403";
        ram_buffer(33430) := X"A602000C";
        ram_buffer(33431) := X"8E030064";
        ram_buffer(33432) := X"2402DFFF";
        ram_buffer(33433) := X"00621024";
        ram_buffer(33434) := X"AE020064";
        ram_buffer(33435) := X"AE000004";
        ram_buffer(33436) := X"8602000C";
        ram_buffer(33437) := X"00000000";
        ram_buffer(33438) := X"3042FFFF";
        ram_buffer(33439) := X"30420020";
        ram_buffer(33440) := X"10400004";
        ram_buffer(33441) := X"00000000";
        ram_buffer(33442) := X"2402FFFF";
        ram_buffer(33443) := X"100000A5";
        ram_buffer(33444) := X"00000000";
        ram_buffer(33445) := X"8602000C";
        ram_buffer(33446) := X"00000000";
        ram_buffer(33447) := X"3042FFFF";
        ram_buffer(33448) := X"30420004";
        ram_buffer(33449) := X"14400032";
        ram_buffer(33450) := X"00000000";
        ram_buffer(33451) := X"8602000C";
        ram_buffer(33452) := X"00000000";
        ram_buffer(33453) := X"3042FFFF";
        ram_buffer(33454) := X"30420010";
        ram_buffer(33455) := X"1440000D";
        ram_buffer(33456) := X"00000000";
        ram_buffer(33457) := X"8FC20028";
        ram_buffer(33458) := X"24030009";
        ram_buffer(33459) := X"AC430000";
        ram_buffer(33460) := X"8602000C";
        ram_buffer(33461) := X"00000000";
        ram_buffer(33462) := X"34420040";
        ram_buffer(33463) := X"00021400";
        ram_buffer(33464) := X"00021403";
        ram_buffer(33465) := X"A602000C";
        ram_buffer(33466) := X"2402FFFF";
        ram_buffer(33467) := X"1000008D";
        ram_buffer(33468) := X"00000000";
        ram_buffer(33469) := X"8602000C";
        ram_buffer(33470) := X"00000000";
        ram_buffer(33471) := X"3042FFFF";
        ram_buffer(33472) := X"30420008";
        ram_buffer(33473) := X"10400012";
        ram_buffer(33474) := X"00000000";
        ram_buffer(33475) := X"02002821";
        ram_buffer(33476) := X"8FC40028";
        ram_buffer(33477) := X"0C026EE1";
        ram_buffer(33478) := X"00000000";
        ram_buffer(33479) := X"10400004";
        ram_buffer(33480) := X"00000000";
        ram_buffer(33481) := X"2402FFFF";
        ram_buffer(33482) := X"1000007E";
        ram_buffer(33483) := X"00000000";
        ram_buffer(33484) := X"8603000C";
        ram_buffer(33485) := X"2402FFF7";
        ram_buffer(33486) := X"00621024";
        ram_buffer(33487) := X"00021400";
        ram_buffer(33488) := X"00021403";
        ram_buffer(33489) := X"A602000C";
        ram_buffer(33490) := X"AE000008";
        ram_buffer(33491) := X"AE000018";
        ram_buffer(33492) := X"8602000C";
        ram_buffer(33493) := X"00000000";
        ram_buffer(33494) := X"34420004";
        ram_buffer(33495) := X"00021400";
        ram_buffer(33496) := X"00021403";
        ram_buffer(33497) := X"A602000C";
        ram_buffer(33498) := X"1000001D";
        ram_buffer(33499) := X"00000000";
        ram_buffer(33500) := X"8E020030";
        ram_buffer(33501) := X"00000000";
        ram_buffer(33502) := X"10400019";
        ram_buffer(33503) := X"00000000";
        ram_buffer(33504) := X"8E030030";
        ram_buffer(33505) := X"26020040";
        ram_buffer(33506) := X"10620007";
        ram_buffer(33507) := X"00000000";
        ram_buffer(33508) := X"8E020030";
        ram_buffer(33509) := X"00000000";
        ram_buffer(33510) := X"00402821";
        ram_buffer(33511) := X"8FC40028";
        ram_buffer(33512) := X"0C027301";
        ram_buffer(33513) := X"00000000";
        ram_buffer(33514) := X"AE000030";
        ram_buffer(33515) := X"8E02003C";
        ram_buffer(33516) := X"00000000";
        ram_buffer(33517) := X"AE020004";
        ram_buffer(33518) := X"8E020004";
        ram_buffer(33519) := X"00000000";
        ram_buffer(33520) := X"10400007";
        ram_buffer(33521) := X"00000000";
        ram_buffer(33522) := X"8E020038";
        ram_buffer(33523) := X"00000000";
        ram_buffer(33524) := X"AE020000";
        ram_buffer(33525) := X"00001021";
        ram_buffer(33526) := X"10000052";
        ram_buffer(33527) := X"00000000";
        ram_buffer(33528) := X"8E020010";
        ram_buffer(33529) := X"00000000";
        ram_buffer(33530) := X"14400005";
        ram_buffer(33531) := X"00000000";
        ram_buffer(33532) := X"02002821";
        ram_buffer(33533) := X"8FC40028";
        ram_buffer(33534) := X"0C027999";
        ram_buffer(33535) := X"00000000";
        ram_buffer(33536) := X"8602000C";
        ram_buffer(33537) := X"00000000";
        ram_buffer(33538) := X"3042FFFF";
        ram_buffer(33539) := X"30420003";
        ram_buffer(33540) := X"1040001A";
        ram_buffer(33541) := X"00000000";
        ram_buffer(33542) := X"9602000C";
        ram_buffer(33543) := X"00000000";
        ram_buffer(33544) := X"A7C20014";
        ram_buffer(33545) := X"24020001";
        ram_buffer(33546) := X"A602000C";
        ram_buffer(33547) := X"8F83809C";
        ram_buffer(33548) := X"3C02100A";
        ram_buffer(33549) := X"24450968";
        ram_buffer(33550) := X"00602021";
        ram_buffer(33551) := X"0C027803";
        ram_buffer(33552) := X"00000000";
        ram_buffer(33553) := X"97C20014";
        ram_buffer(33554) := X"00000000";
        ram_buffer(33555) := X"A602000C";
        ram_buffer(33556) := X"8602000C";
        ram_buffer(33557) := X"00000000";
        ram_buffer(33558) := X"3042FFFF";
        ram_buffer(33559) := X"30430009";
        ram_buffer(33560) := X"24020009";
        ram_buffer(33561) := X"14620005";
        ram_buffer(33562) := X"00000000";
        ram_buffer(33563) := X"02002821";
        ram_buffer(33564) := X"8FC40028";
        ram_buffer(33565) := X"0C026DCB";
        ram_buffer(33566) := X"00000000";
        ram_buffer(33567) := X"8E020010";
        ram_buffer(33568) := X"00000000";
        ram_buffer(33569) := X"AE020000";
        ram_buffer(33570) := X"8E020020";
        ram_buffer(33571) := X"8E03001C";
        ram_buffer(33572) := X"8E040000";
        ram_buffer(33573) := X"8E050014";
        ram_buffer(33574) := X"00000000";
        ram_buffer(33575) := X"00A03821";
        ram_buffer(33576) := X"00803021";
        ram_buffer(33577) := X"00602821";
        ram_buffer(33578) := X"8FC40028";
        ram_buffer(33579) := X"0040F809";
        ram_buffer(33580) := X"00000000";
        ram_buffer(33581) := X"AE020004";
        ram_buffer(33582) := X"8E020004";
        ram_buffer(33583) := X"00000000";
        ram_buffer(33584) := X"1C400017";
        ram_buffer(33585) := X"00000000";
        ram_buffer(33586) := X"8E020004";
        ram_buffer(33587) := X"00000000";
        ram_buffer(33588) := X"14400009";
        ram_buffer(33589) := X"00000000";
        ram_buffer(33590) := X"8602000C";
        ram_buffer(33591) := X"00000000";
        ram_buffer(33592) := X"34420020";
        ram_buffer(33593) := X"00021400";
        ram_buffer(33594) := X"00021403";
        ram_buffer(33595) := X"A602000C";
        ram_buffer(33596) := X"10000008";
        ram_buffer(33597) := X"00000000";
        ram_buffer(33598) := X"AE000004";
        ram_buffer(33599) := X"8602000C";
        ram_buffer(33600) := X"00000000";
        ram_buffer(33601) := X"34420040";
        ram_buffer(33602) := X"00021400";
        ram_buffer(33603) := X"00021403";
        ram_buffer(33604) := X"A602000C";
        ram_buffer(33605) := X"2402FFFF";
        ram_buffer(33606) := X"10000002";
        ram_buffer(33607) := X"00000000";
        ram_buffer(33608) := X"00001021";
        ram_buffer(33609) := X"03C0E821";
        ram_buffer(33610) := X"8FBF0024";
        ram_buffer(33611) := X"8FBE0020";
        ram_buffer(33612) := X"8FB0001C";
        ram_buffer(33613) := X"27BD0028";
        ram_buffer(33614) := X"03E00008";
        ram_buffer(33615) := X"00000000";
        ram_buffer(33616) := X"27BDFFD8";
        ram_buffer(33617) := X"AFBF0024";
        ram_buffer(33618) := X"AFBE0020";
        ram_buffer(33619) := X"AFB0001C";
        ram_buffer(33620) := X"03A0F021";
        ram_buffer(33621) := X"AFC40028";
        ram_buffer(33622) := X"00A08021";
        ram_buffer(33623) := X"8FC20028";
        ram_buffer(33624) := X"00000000";
        ram_buffer(33625) := X"AFC20010";
        ram_buffer(33626) := X"8FC20010";
        ram_buffer(33627) := X"00000000";
        ram_buffer(33628) := X"1040000A";
        ram_buffer(33629) := X"00000000";
        ram_buffer(33630) := X"8FC20010";
        ram_buffer(33631) := X"00000000";
        ram_buffer(33632) := X"8C420038";
        ram_buffer(33633) := X"00000000";
        ram_buffer(33634) := X"14400004";
        ram_buffer(33635) := X"00000000";
        ram_buffer(33636) := X"8FC40010";
        ram_buffer(33637) := X"0C027069";
        ram_buffer(33638) := X"00000000";
        ram_buffer(33639) := X"02002821";
        ram_buffer(33640) := X"8FC40028";
        ram_buffer(33641) := X"0C028274";
        ram_buffer(33642) := X"00000000";
        ram_buffer(33643) := X"1440000C";
        ram_buffer(33644) := X"00000000";
        ram_buffer(33645) := X"8E020004";
        ram_buffer(33646) := X"00000000";
        ram_buffer(33647) := X"2442FFFF";
        ram_buffer(33648) := X"AE020004";
        ram_buffer(33649) := X"8E020000";
        ram_buffer(33650) := X"00000000";
        ram_buffer(33651) := X"24430001";
        ram_buffer(33652) := X"AE030000";
        ram_buffer(33653) := X"90420000";
        ram_buffer(33654) := X"10000002";
        ram_buffer(33655) := X"00000000";
        ram_buffer(33656) := X"2402FFFF";
        ram_buffer(33657) := X"03C0E821";
        ram_buffer(33658) := X"8FBF0024";
        ram_buffer(33659) := X"8FBE0020";
        ram_buffer(33660) := X"8FB0001C";
        ram_buffer(33661) := X"27BD0028";
        ram_buffer(33662) := X"03E00008";
        ram_buffer(33663) := X"00000000";
        ram_buffer(33664) := X"27BDFFE8";
        ram_buffer(33665) := X"AFBF0014";
        ram_buffer(33666) := X"AFBE0010";
        ram_buffer(33667) := X"03A0F021";
        ram_buffer(33668) := X"00801821";
        ram_buffer(33669) := X"8F828098";
        ram_buffer(33670) := X"00602821";
        ram_buffer(33671) := X"00402021";
        ram_buffer(33672) := X"0C028350";
        ram_buffer(33673) := X"00000000";
        ram_buffer(33674) := X"03C0E821";
        ram_buffer(33675) := X"8FBF0014";
        ram_buffer(33676) := X"8FBE0010";
        ram_buffer(33677) := X"27BD0018";
        ram_buffer(33678) := X"03E00008";
        ram_buffer(33679) := X"00000000";
        ram_buffer(33680) := X"27BDFFE0";
        ram_buffer(33681) := X"AFBF001C";
        ram_buffer(33682) := X"AFBE0018";
        ram_buffer(33683) := X"03A0F021";
        ram_buffer(33684) := X"AFC40020";
        ram_buffer(33685) := X"AFC50024";
        ram_buffer(33686) := X"AF8081EC";
        ram_buffer(33687) := X"8FC40024";
        ram_buffer(33688) := X"0C02FC7B";
        ram_buffer(33689) := X"00000000";
        ram_buffer(33690) := X"AFC20010";
        ram_buffer(33691) := X"8FC30010";
        ram_buffer(33692) := X"2402FFFF";
        ram_buffer(33693) := X"14620009";
        ram_buffer(33694) := X"00000000";
        ram_buffer(33695) := X"8F8281EC";
        ram_buffer(33696) := X"00000000";
        ram_buffer(33697) := X"10400005";
        ram_buffer(33698) := X"00000000";
        ram_buffer(33699) := X"8F8381EC";
        ram_buffer(33700) := X"8FC20020";
        ram_buffer(33701) := X"00000000";
        ram_buffer(33702) := X"AC430000";
        ram_buffer(33703) := X"8FC20010";
        ram_buffer(33704) := X"03C0E821";
        ram_buffer(33705) := X"8FBF001C";
        ram_buffer(33706) := X"8FBE0018";
        ram_buffer(33707) := X"27BD0020";
        ram_buffer(33708) := X"03E00008";
        ram_buffer(33709) := X"00000000";
        ram_buffer(33710) := X"27BDFF78";
        ram_buffer(33711) := X"AFBF0084";
        ram_buffer(33712) := X"AFBE0080";
        ram_buffer(33713) := X"03A0F021";
        ram_buffer(33714) := X"AFC40088";
        ram_buffer(33715) := X"AFC5008C";
        ram_buffer(33716) := X"AFC60090";
        ram_buffer(33717) := X"AFC70094";
        ram_buffer(33718) := X"24020208";
        ram_buffer(33719) := X"A7C20024";
        ram_buffer(33720) := X"8FC2008C";
        ram_buffer(33721) := X"00000000";
        ram_buffer(33722) := X"AFC20018";
        ram_buffer(33723) := X"8FC20018";
        ram_buffer(33724) := X"00000000";
        ram_buffer(33725) := X"AFC20028";
        ram_buffer(33726) := X"3C027FFF";
        ram_buffer(33727) := X"3442FFFF";
        ram_buffer(33728) := X"AFC20020";
        ram_buffer(33729) := X"8FC20020";
        ram_buffer(33730) := X"00000000";
        ram_buffer(33731) := X"AFC2002C";
        ram_buffer(33732) := X"2402FFFF";
        ram_buffer(33733) := X"A7C20026";
        ram_buffer(33734) := X"27C20094";
        ram_buffer(33735) := X"AFC20014";
        ram_buffer(33736) := X"8FC30014";
        ram_buffer(33737) := X"27C20018";
        ram_buffer(33738) := X"00603821";
        ram_buffer(33739) := X"8FC60090";
        ram_buffer(33740) := X"00402821";
        ram_buffer(33741) := X"8FC40088";
        ram_buffer(33742) := X"0C0285AE";
        ram_buffer(33743) := X"00000000";
        ram_buffer(33744) := X"AFC20010";
        ram_buffer(33745) := X"8FC20018";
        ram_buffer(33746) := X"00000000";
        ram_buffer(33747) := X"A0400000";
        ram_buffer(33748) := X"8FC20010";
        ram_buffer(33749) := X"03C0E821";
        ram_buffer(33750) := X"8FBF0084";
        ram_buffer(33751) := X"8FBE0080";
        ram_buffer(33752) := X"27BD0088";
        ram_buffer(33753) := X"03E00008";
        ram_buffer(33754) := X"00000000";
        ram_buffer(33755) := X"27BDFF78";
        ram_buffer(33756) := X"AFBF0084";
        ram_buffer(33757) := X"AFBE0080";
        ram_buffer(33758) := X"03A0F021";
        ram_buffer(33759) := X"AFC40088";
        ram_buffer(33760) := X"AFC5008C";
        ram_buffer(33761) := X"AFC60090";
        ram_buffer(33762) := X"AFC70094";
        ram_buffer(33763) := X"24020208";
        ram_buffer(33764) := X"A7C20024";
        ram_buffer(33765) := X"8FC20088";
        ram_buffer(33766) := X"00000000";
        ram_buffer(33767) := X"AFC20018";
        ram_buffer(33768) := X"8FC20018";
        ram_buffer(33769) := X"00000000";
        ram_buffer(33770) := X"AFC20028";
        ram_buffer(33771) := X"3C027FFF";
        ram_buffer(33772) := X"3442FFFF";
        ram_buffer(33773) := X"AFC20020";
        ram_buffer(33774) := X"8FC20020";
        ram_buffer(33775) := X"00000000";
        ram_buffer(33776) := X"AFC2002C";
        ram_buffer(33777) := X"2402FFFF";
        ram_buffer(33778) := X"A7C20026";
        ram_buffer(33779) := X"27C20090";
        ram_buffer(33780) := X"AFC20014";
        ram_buffer(33781) := X"8F828098";
        ram_buffer(33782) := X"8FC40014";
        ram_buffer(33783) := X"27C30018";
        ram_buffer(33784) := X"00803821";
        ram_buffer(33785) := X"8FC6008C";
        ram_buffer(33786) := X"00602821";
        ram_buffer(33787) := X"00402021";
        ram_buffer(33788) := X"0C0285AE";
        ram_buffer(33789) := X"00000000";
        ram_buffer(33790) := X"AFC20010";
        ram_buffer(33791) := X"8FC20018";
        ram_buffer(33792) := X"00000000";
        ram_buffer(33793) := X"A0400000";
        ram_buffer(33794) := X"8FC20010";
        ram_buffer(33795) := X"03C0E821";
        ram_buffer(33796) := X"8FBF0084";
        ram_buffer(33797) := X"8FBE0080";
        ram_buffer(33798) := X"27BD0088";
        ram_buffer(33799) := X"03E00008";
        ram_buffer(33800) := X"00000000";
        ram_buffer(33801) := X"27BDFF78";
        ram_buffer(33802) := X"AFBF0084";
        ram_buffer(33803) := X"AFBE0080";
        ram_buffer(33804) := X"03A0F021";
        ram_buffer(33805) := X"AFC40088";
        ram_buffer(33806) := X"AFC5008C";
        ram_buffer(33807) := X"AFC60090";
        ram_buffer(33808) := X"AFC70094";
        ram_buffer(33809) := X"24020204";
        ram_buffer(33810) := X"A7C20024";
        ram_buffer(33811) := X"8FC20088";
        ram_buffer(33812) := X"00000000";
        ram_buffer(33813) := X"AFC20018";
        ram_buffer(33814) := X"8FC20018";
        ram_buffer(33815) := X"00000000";
        ram_buffer(33816) := X"AFC20028";
        ram_buffer(33817) := X"8FC40088";
        ram_buffer(33818) := X"0C02851E";
        ram_buffer(33819) := X"00000000";
        ram_buffer(33820) := X"AFC2001C";
        ram_buffer(33821) := X"8FC2001C";
        ram_buffer(33822) := X"00000000";
        ram_buffer(33823) := X"AFC2002C";
        ram_buffer(33824) := X"3C02100A";
        ram_buffer(33825) := X"24421264";
        ram_buffer(33826) := X"AFC20038";
        ram_buffer(33827) := X"AFC00048";
        ram_buffer(33828) := X"AFC0005C";
        ram_buffer(33829) := X"2402FFFF";
        ram_buffer(33830) := X"A7C20026";
        ram_buffer(33831) := X"27C20090";
        ram_buffer(33832) := X"AFC20014";
        ram_buffer(33833) := X"8F828098";
        ram_buffer(33834) := X"8FC40014";
        ram_buffer(33835) := X"27C30018";
        ram_buffer(33836) := X"00803821";
        ram_buffer(33837) := X"8FC6008C";
        ram_buffer(33838) := X"00602821";
        ram_buffer(33839) := X"00402021";
        ram_buffer(33840) := X"0C029456";
        ram_buffer(33841) := X"00000000";
        ram_buffer(33842) := X"AFC20010";
        ram_buffer(33843) := X"8FC20010";
        ram_buffer(33844) := X"03C0E821";
        ram_buffer(33845) := X"8FBF0084";
        ram_buffer(33846) := X"8FBE0080";
        ram_buffer(33847) := X"27BD0088";
        ram_buffer(33848) := X"03E00008";
        ram_buffer(33849) := X"00000000";
        ram_buffer(33850) := X"27BDFF78";
        ram_buffer(33851) := X"AFBF0084";
        ram_buffer(33852) := X"AFBE0080";
        ram_buffer(33853) := X"03A0F021";
        ram_buffer(33854) := X"AFC40088";
        ram_buffer(33855) := X"AFC5008C";
        ram_buffer(33856) := X"AFC60090";
        ram_buffer(33857) := X"AFC70094";
        ram_buffer(33858) := X"24020204";
        ram_buffer(33859) := X"A7C20024";
        ram_buffer(33860) := X"8FC2008C";
        ram_buffer(33861) := X"00000000";
        ram_buffer(33862) := X"AFC20018";
        ram_buffer(33863) := X"8FC20018";
        ram_buffer(33864) := X"00000000";
        ram_buffer(33865) := X"AFC20028";
        ram_buffer(33866) := X"8FC4008C";
        ram_buffer(33867) := X"0C02851E";
        ram_buffer(33868) := X"00000000";
        ram_buffer(33869) := X"AFC2001C";
        ram_buffer(33870) := X"8FC2001C";
        ram_buffer(33871) := X"00000000";
        ram_buffer(33872) := X"AFC2002C";
        ram_buffer(33873) := X"3C02100A";
        ram_buffer(33874) := X"24421264";
        ram_buffer(33875) := X"AFC20038";
        ram_buffer(33876) := X"AFC00048";
        ram_buffer(33877) := X"AFC0005C";
        ram_buffer(33878) := X"2402FFFF";
        ram_buffer(33879) := X"A7C20026";
        ram_buffer(33880) := X"27C20094";
        ram_buffer(33881) := X"AFC20014";
        ram_buffer(33882) := X"8FC30014";
        ram_buffer(33883) := X"27C20018";
        ram_buffer(33884) := X"00603821";
        ram_buffer(33885) := X"8FC60090";
        ram_buffer(33886) := X"00402821";
        ram_buffer(33887) := X"8FC40088";
        ram_buffer(33888) := X"0C029456";
        ram_buffer(33889) := X"00000000";
        ram_buffer(33890) := X"AFC20010";
        ram_buffer(33891) := X"8FC20010";
        ram_buffer(33892) := X"03C0E821";
        ram_buffer(33893) := X"8FBF0084";
        ram_buffer(33894) := X"8FBE0080";
        ram_buffer(33895) := X"27BD0088";
        ram_buffer(33896) := X"03E00008";
        ram_buffer(33897) := X"00000000";
        ram_buffer(33898) := X"27BDFFE0";
        ram_buffer(33899) := X"AFBF001C";
        ram_buffer(33900) := X"AFBE0018";
        ram_buffer(33901) := X"AFB10014";
        ram_buffer(33902) := X"AFB00010";
        ram_buffer(33903) := X"03A0F021";
        ram_buffer(33904) := X"AFC40020";
        ram_buffer(33905) := X"AFC50024";
        ram_buffer(33906) := X"AFC60028";
        ram_buffer(33907) := X"AFC7002C";
        ram_buffer(33908) := X"8FD00024";
        ram_buffer(33909) := X"00000000";
        ram_buffer(33910) := X"8602000E";
        ram_buffer(33911) := X"00000000";
        ram_buffer(33912) := X"00401821";
        ram_buffer(33913) := X"8FC2002C";
        ram_buffer(33914) := X"00000000";
        ram_buffer(33915) := X"00403821";
        ram_buffer(33916) := X"8FC60028";
        ram_buffer(33917) := X"00602821";
        ram_buffer(33918) := X"8FC40020";
        ram_buffer(33919) := X"0C02C685";
        ram_buffer(33920) := X"00000000";
        ram_buffer(33921) := X"00408821";
        ram_buffer(33922) := X"06200007";
        ram_buffer(33923) := X"00000000";
        ram_buffer(33924) := X"8E020050";
        ram_buffer(33925) := X"00000000";
        ram_buffer(33926) := X"00511021";
        ram_buffer(33927) := X"AE020050";
        ram_buffer(33928) := X"10000007";
        ram_buffer(33929) := X"00000000";
        ram_buffer(33930) := X"8603000C";
        ram_buffer(33931) := X"2402EFFF";
        ram_buffer(33932) := X"00621024";
        ram_buffer(33933) := X"00021400";
        ram_buffer(33934) := X"00021403";
        ram_buffer(33935) := X"A602000C";
        ram_buffer(33936) := X"02201021";
        ram_buffer(33937) := X"03C0E821";
        ram_buffer(33938) := X"8FBF001C";
        ram_buffer(33939) := X"8FBE0018";
        ram_buffer(33940) := X"8FB10014";
        ram_buffer(33941) := X"8FB00010";
        ram_buffer(33942) := X"27BD0020";
        ram_buffer(33943) := X"03E00008";
        ram_buffer(33944) := X"00000000";
        ram_buffer(33945) := X"27BDFFF8";
        ram_buffer(33946) := X"AFBE0004";
        ram_buffer(33947) := X"03A0F021";
        ram_buffer(33948) := X"AFC40008";
        ram_buffer(33949) := X"AFC5000C";
        ram_buffer(33950) := X"AFC60010";
        ram_buffer(33951) := X"AFC70014";
        ram_buffer(33952) := X"00001021";
        ram_buffer(33953) := X"03C0E821";
        ram_buffer(33954) := X"8FBE0004";
        ram_buffer(33955) := X"27BD0008";
        ram_buffer(33956) := X"03E00008";
        ram_buffer(33957) := X"00000000";
        ram_buffer(33958) := X"27BDFFD8";
        ram_buffer(33959) := X"AFBF0024";
        ram_buffer(33960) := X"AFBE0020";
        ram_buffer(33961) := X"AFB0001C";
        ram_buffer(33962) := X"03A0F021";
        ram_buffer(33963) := X"AFC40028";
        ram_buffer(33964) := X"AFC5002C";
        ram_buffer(33965) := X"AFC60030";
        ram_buffer(33966) := X"AFC70034";
        ram_buffer(33967) := X"8FD0002C";
        ram_buffer(33968) := X"00000000";
        ram_buffer(33969) := X"8602000C";
        ram_buffer(33970) := X"00000000";
        ram_buffer(33971) := X"3042FFFF";
        ram_buffer(33972) := X"30420100";
        ram_buffer(33973) := X"10400008";
        ram_buffer(33974) := X"00000000";
        ram_buffer(33975) := X"8602000E";
        ram_buffer(33976) := X"24070002";
        ram_buffer(33977) := X"00003021";
        ram_buffer(33978) := X"00402821";
        ram_buffer(33979) := X"8FC40028";
        ram_buffer(33980) := X"0C02BB51";
        ram_buffer(33981) := X"00000000";
        ram_buffer(33982) := X"8603000C";
        ram_buffer(33983) := X"2402EFFF";
        ram_buffer(33984) := X"00621024";
        ram_buffer(33985) := X"00021400";
        ram_buffer(33986) := X"00021403";
        ram_buffer(33987) := X"A602000C";
        ram_buffer(33988) := X"8602000E";
        ram_buffer(33989) := X"00000000";
        ram_buffer(33990) := X"00401821";
        ram_buffer(33991) := X"8FC20034";
        ram_buffer(33992) := X"00000000";
        ram_buffer(33993) := X"00403821";
        ram_buffer(33994) := X"8FC60030";
        ram_buffer(33995) := X"00602821";
        ram_buffer(33996) := X"8FC40028";
        ram_buffer(33997) := X"0C02ACCF";
        ram_buffer(33998) := X"00000000";
        ram_buffer(33999) := X"AFC20010";
        ram_buffer(34000) := X"8FC20010";
        ram_buffer(34001) := X"03C0E821";
        ram_buffer(34002) := X"8FBF0024";
        ram_buffer(34003) := X"8FBE0020";
        ram_buffer(34004) := X"8FB0001C";
        ram_buffer(34005) := X"27BD0028";
        ram_buffer(34006) := X"03E00008";
        ram_buffer(34007) := X"00000000";
        ram_buffer(34008) := X"27BDFFE0";
        ram_buffer(34009) := X"AFBF001C";
        ram_buffer(34010) := X"AFBE0018";
        ram_buffer(34011) := X"AFB10014";
        ram_buffer(34012) := X"AFB00010";
        ram_buffer(34013) := X"03A0F021";
        ram_buffer(34014) := X"AFC40020";
        ram_buffer(34015) := X"AFC50024";
        ram_buffer(34016) := X"AFC60028";
        ram_buffer(34017) := X"AFC7002C";
        ram_buffer(34018) := X"8FD00024";
        ram_buffer(34019) := X"00000000";
        ram_buffer(34020) := X"8602000E";
        ram_buffer(34021) := X"8FC7002C";
        ram_buffer(34022) := X"8FC60028";
        ram_buffer(34023) := X"00402821";
        ram_buffer(34024) := X"8FC40020";
        ram_buffer(34025) := X"0C02BB51";
        ram_buffer(34026) := X"00000000";
        ram_buffer(34027) := X"00408821";
        ram_buffer(34028) := X"2402FFFF";
        ram_buffer(34029) := X"16220009";
        ram_buffer(34030) := X"00000000";
        ram_buffer(34031) := X"8603000C";
        ram_buffer(34032) := X"2402EFFF";
        ram_buffer(34033) := X"00621024";
        ram_buffer(34034) := X"00021400";
        ram_buffer(34035) := X"00021403";
        ram_buffer(34036) := X"A602000C";
        ram_buffer(34037) := X"10000008";
        ram_buffer(34038) := X"00000000";
        ram_buffer(34039) := X"8602000C";
        ram_buffer(34040) := X"00000000";
        ram_buffer(34041) := X"34421000";
        ram_buffer(34042) := X"00021400";
        ram_buffer(34043) := X"00021403";
        ram_buffer(34044) := X"A602000C";
        ram_buffer(34045) := X"AE110050";
        ram_buffer(34046) := X"02201021";
        ram_buffer(34047) := X"03C0E821";
        ram_buffer(34048) := X"8FBF001C";
        ram_buffer(34049) := X"8FBE0018";
        ram_buffer(34050) := X"8FB10014";
        ram_buffer(34051) := X"8FB00010";
        ram_buffer(34052) := X"27BD0020";
        ram_buffer(34053) := X"03E00008";
        ram_buffer(34054) := X"00000000";
        ram_buffer(34055) := X"27BDFFE0";
        ram_buffer(34056) := X"AFBF001C";
        ram_buffer(34057) := X"AFBE0018";
        ram_buffer(34058) := X"03A0F021";
        ram_buffer(34059) := X"AFC40020";
        ram_buffer(34060) := X"AFC50024";
        ram_buffer(34061) := X"8FC20024";
        ram_buffer(34062) := X"00000000";
        ram_buffer(34063) := X"AFC20010";
        ram_buffer(34064) := X"8FC20010";
        ram_buffer(34065) := X"00000000";
        ram_buffer(34066) := X"8442000E";
        ram_buffer(34067) := X"00000000";
        ram_buffer(34068) := X"00402821";
        ram_buffer(34069) := X"8FC40020";
        ram_buffer(34070) := X"0C02AE34";
        ram_buffer(34071) := X"00000000";
        ram_buffer(34072) := X"03C0E821";
        ram_buffer(34073) := X"8FBF001C";
        ram_buffer(34074) := X"8FBE0018";
        ram_buffer(34075) := X"27BD0020";
        ram_buffer(34076) := X"03E00008";
        ram_buffer(34077) := X"00000000";
        ram_buffer(34078) := X"24820001";
        ram_buffer(34079) := X"90830000";
        ram_buffer(34080) := X"00000000";
        ram_buffer(34081) := X"1460FFFD";
        ram_buffer(34082) := X"24840001";
        ram_buffer(34083) := X"03E00008";
        ram_buffer(34084) := X"00821023";
        ram_buffer(34085) := X"27BDFFF0";
        ram_buffer(34086) := X"AFBE000C";
        ram_buffer(34087) := X"03A0F021";
        ram_buffer(34088) := X"AFC40010";
        ram_buffer(34089) := X"AFC50014";
        ram_buffer(34090) := X"AFC60018";
        ram_buffer(34091) := X"8FC20018";
        ram_buffer(34092) := X"00000000";
        ram_buffer(34093) := X"14400004";
        ram_buffer(34094) := X"00000000";
        ram_buffer(34095) := X"00001021";
        ram_buffer(34096) := X"10000078";
        ram_buffer(34097) := X"00000000";
        ram_buffer(34098) := X"8FC30010";
        ram_buffer(34099) := X"8FC20014";
        ram_buffer(34100) := X"00000000";
        ram_buffer(34101) := X"00621025";
        ram_buffer(34102) := X"30420003";
        ram_buffer(34103) := X"14400058";
        ram_buffer(34104) := X"00000000";
        ram_buffer(34105) := X"8FC20010";
        ram_buffer(34106) := X"00000000";
        ram_buffer(34107) := X"AFC20000";
        ram_buffer(34108) := X"8FC20014";
        ram_buffer(34109) := X"00000000";
        ram_buffer(34110) := X"AFC20004";
        ram_buffer(34111) := X"10000025";
        ram_buffer(34112) := X"00000000";
        ram_buffer(34113) := X"8FC20018";
        ram_buffer(34114) := X"00000000";
        ram_buffer(34115) := X"2442FFFC";
        ram_buffer(34116) := X"AFC20018";
        ram_buffer(34117) := X"8FC20018";
        ram_buffer(34118) := X"00000000";
        ram_buffer(34119) := X"10400012";
        ram_buffer(34120) := X"00000000";
        ram_buffer(34121) := X"8FC20000";
        ram_buffer(34122) := X"00000000";
        ram_buffer(34123) := X"8C430000";
        ram_buffer(34124) := X"3C02FEFE";
        ram_buffer(34125) := X"3442FEFF";
        ram_buffer(34126) := X"00621821";
        ram_buffer(34127) := X"8FC20000";
        ram_buffer(34128) := X"00000000";
        ram_buffer(34129) := X"8C420000";
        ram_buffer(34130) := X"00000000";
        ram_buffer(34131) := X"00021027";
        ram_buffer(34132) := X"00621824";
        ram_buffer(34133) := X"3C028080";
        ram_buffer(34134) := X"34428080";
        ram_buffer(34135) := X"00621024";
        ram_buffer(34136) := X"10400004";
        ram_buffer(34137) := X"00000000";
        ram_buffer(34138) := X"00001021";
        ram_buffer(34139) := X"1000004D";
        ram_buffer(34140) := X"00000000";
        ram_buffer(34141) := X"8FC20000";
        ram_buffer(34142) := X"00000000";
        ram_buffer(34143) := X"24420004";
        ram_buffer(34144) := X"AFC20000";
        ram_buffer(34145) := X"8FC20004";
        ram_buffer(34146) := X"00000000";
        ram_buffer(34147) := X"24420004";
        ram_buffer(34148) := X"AFC20004";
        ram_buffer(34149) := X"8FC20018";
        ram_buffer(34150) := X"00000000";
        ram_buffer(34151) := X"2C420004";
        ram_buffer(34152) := X"1440000A";
        ram_buffer(34153) := X"00000000";
        ram_buffer(34154) := X"8FC20000";
        ram_buffer(34155) := X"00000000";
        ram_buffer(34156) := X"8C430000";
        ram_buffer(34157) := X"8FC20004";
        ram_buffer(34158) := X"00000000";
        ram_buffer(34159) := X"8C420000";
        ram_buffer(34160) := X"00000000";
        ram_buffer(34161) := X"1062FFCF";
        ram_buffer(34162) := X"00000000";
        ram_buffer(34163) := X"8FC20000";
        ram_buffer(34164) := X"00000000";
        ram_buffer(34165) := X"AFC20010";
        ram_buffer(34166) := X"8FC20004";
        ram_buffer(34167) := X"00000000";
        ram_buffer(34168) := X"AFC20014";
        ram_buffer(34169) := X"10000016";
        ram_buffer(34170) := X"00000000";
        ram_buffer(34171) := X"8FC20018";
        ram_buffer(34172) := X"00000000";
        ram_buffer(34173) := X"10400007";
        ram_buffer(34174) := X"00000000";
        ram_buffer(34175) := X"8FC20010";
        ram_buffer(34176) := X"00000000";
        ram_buffer(34177) := X"80420000";
        ram_buffer(34178) := X"00000000";
        ram_buffer(34179) := X"14400004";
        ram_buffer(34180) := X"00000000";
        ram_buffer(34181) := X"00001021";
        ram_buffer(34182) := X"10000022";
        ram_buffer(34183) := X"00000000";
        ram_buffer(34184) := X"8FC20010";
        ram_buffer(34185) := X"00000000";
        ram_buffer(34186) := X"24420001";
        ram_buffer(34187) := X"AFC20010";
        ram_buffer(34188) := X"8FC20014";
        ram_buffer(34189) := X"00000000";
        ram_buffer(34190) := X"24420001";
        ram_buffer(34191) := X"AFC20014";
        ram_buffer(34192) := X"8FC20018";
        ram_buffer(34193) := X"00000000";
        ram_buffer(34194) := X"2443FFFF";
        ram_buffer(34195) := X"AFC30018";
        ram_buffer(34196) := X"1040000A";
        ram_buffer(34197) := X"00000000";
        ram_buffer(34198) := X"8FC20010";
        ram_buffer(34199) := X"00000000";
        ram_buffer(34200) := X"80430000";
        ram_buffer(34201) := X"8FC20014";
        ram_buffer(34202) := X"00000000";
        ram_buffer(34203) := X"80420000";
        ram_buffer(34204) := X"00000000";
        ram_buffer(34205) := X"1062FFDD";
        ram_buffer(34206) := X"00000000";
        ram_buffer(34207) := X"8FC20010";
        ram_buffer(34208) := X"00000000";
        ram_buffer(34209) := X"90420000";
        ram_buffer(34210) := X"00000000";
        ram_buffer(34211) := X"00401821";
        ram_buffer(34212) := X"8FC20014";
        ram_buffer(34213) := X"00000000";
        ram_buffer(34214) := X"90420000";
        ram_buffer(34215) := X"00000000";
        ram_buffer(34216) := X"00621023";
        ram_buffer(34217) := X"03C0E821";
        ram_buffer(34218) := X"8FBE000C";
        ram_buffer(34219) := X"27BD0010";
        ram_buffer(34220) := X"03E00008";
        ram_buffer(34221) := X"00000000";
        ram_buffer(34222) := X"27BDFE18";
        ram_buffer(34223) := X"AFBF01E4";
        ram_buffer(34224) := X"AFBE01E0";
        ram_buffer(34225) := X"AFB701DC";
        ram_buffer(34226) := X"AFB601D8";
        ram_buffer(34227) := X"AFB501D4";
        ram_buffer(34228) := X"AFB401D0";
        ram_buffer(34229) := X"AFB301CC";
        ram_buffer(34230) := X"AFB201C8";
        ram_buffer(34231) := X"AFB101C4";
        ram_buffer(34232) := X"AFB001C0";
        ram_buffer(34233) := X"03A0F021";
        ram_buffer(34234) := X"AFC401E8";
        ram_buffer(34235) := X"AFC501EC";
        ram_buffer(34236) := X"AFC601F0";
        ram_buffer(34237) := X"AFC701F4";
        ram_buffer(34238) := X"AFC0003C";
        ram_buffer(34239) := X"AFC00040";
        ram_buffer(34240) := X"AFC00044";
        ram_buffer(34241) := X"8FC401E8";
        ram_buffer(34242) := X"0C02BB25";
        ram_buffer(34243) := X"00000000";
        ram_buffer(34244) := X"8C420000";
        ram_buffer(34245) := X"00000000";
        ram_buffer(34246) := X"AFC20084";
        ram_buffer(34247) := X"8FC40084";
        ram_buffer(34248) := X"0C02851E";
        ram_buffer(34249) := X"00000000";
        ram_buffer(34250) := X"AFC20088";
        ram_buffer(34251) := X"00001821";
        ram_buffer(34252) := X"00001021";
        ram_buffer(34253) := X"AFC300A4";
        ram_buffer(34254) := X"AFC200A0";
        ram_buffer(34255) := X"AFC00048";
        ram_buffer(34256) := X"AFC000B4";
        ram_buffer(34257) := X"AFC00070";
        ram_buffer(34258) := X"AFC00074";
        ram_buffer(34259) := X"8FC201EC";
        ram_buffer(34260) := X"00000000";
        ram_buffer(34261) := X"8442000C";
        ram_buffer(34262) := X"00000000";
        ram_buffer(34263) := X"3042FFFF";
        ram_buffer(34264) := X"30420080";
        ram_buffer(34265) := X"10400024";
        ram_buffer(34266) := X"00000000";
        ram_buffer(34267) := X"8FC201EC";
        ram_buffer(34268) := X"00000000";
        ram_buffer(34269) := X"8C420010";
        ram_buffer(34270) := X"00000000";
        ram_buffer(34271) := X"1440001E";
        ram_buffer(34272) := X"00000000";
        ram_buffer(34273) := X"24050040";
        ram_buffer(34274) := X"8FC401E8";
        ram_buffer(34275) := X"0C027B8F";
        ram_buffer(34276) := X"00000000";
        ram_buffer(34277) := X"00401821";
        ram_buffer(34278) := X"8FC201EC";
        ram_buffer(34279) := X"00000000";
        ram_buffer(34280) := X"AC430000";
        ram_buffer(34281) := X"8FC201EC";
        ram_buffer(34282) := X"00000000";
        ram_buffer(34283) := X"8C430000";
        ram_buffer(34284) := X"8FC201EC";
        ram_buffer(34285) := X"00000000";
        ram_buffer(34286) := X"AC430010";
        ram_buffer(34287) := X"8FC201EC";
        ram_buffer(34288) := X"00000000";
        ram_buffer(34289) := X"8C420000";
        ram_buffer(34290) := X"00000000";
        ram_buffer(34291) := X"14400007";
        ram_buffer(34292) := X"00000000";
        ram_buffer(34293) := X"8FC201E8";
        ram_buffer(34294) := X"2403000C";
        ram_buffer(34295) := X"AC430000";
        ram_buffer(34296) := X"2402FFFF";
        ram_buffer(34297) := X"10000C54";
        ram_buffer(34298) := X"00000000";
        ram_buffer(34299) := X"8FC201EC";
        ram_buffer(34300) := X"24030040";
        ram_buffer(34301) := X"AC430014";
        ram_buffer(34302) := X"8FD501F0";
        ram_buffer(34303) := X"27D000C4";
        ram_buffer(34304) := X"AFD000B8";
        ram_buffer(34305) := X"AFC000C0";
        ram_buffer(34306) := X"AFC000BC";
        ram_buffer(34307) := X"AFC00030";
        ram_buffer(34308) := X"02A09821";
        ram_buffer(34309) := X"10000002";
        ram_buffer(34310) := X"00000000";
        ram_buffer(34311) := X"26B50001";
        ram_buffer(34312) := X"82A20000";
        ram_buffer(34313) := X"00000000";
        ram_buffer(34314) := X"10400005";
        ram_buffer(34315) := X"00000000";
        ram_buffer(34316) := X"82A30000";
        ram_buffer(34317) := X"24020025";
        ram_buffer(34318) := X"1462FFF8";
        ram_buffer(34319) := X"00000000";
        ram_buffer(34320) := X"02A01821";
        ram_buffer(34321) := X"02601021";
        ram_buffer(34322) := X"00628823";
        ram_buffer(34323) := X"1220001F";
        ram_buffer(34324) := X"00000000";
        ram_buffer(34325) := X"AE130000";
        ram_buffer(34326) := X"02201021";
        ram_buffer(34327) := X"AE020004";
        ram_buffer(34328) := X"8FC300C0";
        ram_buffer(34329) := X"02201021";
        ram_buffer(34330) := X"00621021";
        ram_buffer(34331) := X"AFC200C0";
        ram_buffer(34332) := X"26100008";
        ram_buffer(34333) := X"8FC200BC";
        ram_buffer(34334) := X"00000000";
        ram_buffer(34335) := X"24420001";
        ram_buffer(34336) := X"AFC200BC";
        ram_buffer(34337) := X"8FC200BC";
        ram_buffer(34338) := X"00000000";
        ram_buffer(34339) := X"28420008";
        ram_buffer(34340) := X"1440000A";
        ram_buffer(34341) := X"00000000";
        ram_buffer(34342) := X"27C200B8";
        ram_buffer(34343) := X"00403021";
        ram_buffer(34344) := X"8FC501EC";
        ram_buffer(34345) := X"8FC401E8";
        ram_buffer(34346) := X"0C02DCA6";
        ram_buffer(34347) := X"00000000";
        ram_buffer(34348) := X"14400B93";
        ram_buffer(34349) := X"00000000";
        ram_buffer(34350) := X"27D000C4";
        ram_buffer(34351) := X"8FC20030";
        ram_buffer(34352) := X"00000000";
        ram_buffer(34353) := X"00511021";
        ram_buffer(34354) := X"AFC20030";
        ram_buffer(34355) := X"82A20000";
        ram_buffer(34356) := X"00000000";
        ram_buffer(34357) := X"10400B76";
        ram_buffer(34358) := X"00000000";
        ram_buffer(34359) := X"AFD5008C";
        ram_buffer(34360) := X"26B50001";
        ram_buffer(34361) := X"00009021";
        ram_buffer(34362) := X"AFC00064";
        ram_buffer(34363) := X"AFC00034";
        ram_buffer(34364) := X"2402FFFF";
        ram_buffer(34365) := X"AFC20038";
        ram_buffer(34366) := X"A3C00098";
        ram_buffer(34367) := X"AFC0004C";
        ram_buffer(34368) := X"AFC00054";
        ram_buffer(34369) := X"8FC20054";
        ram_buffer(34370) := X"00000000";
        ram_buffer(34371) := X"AFC20050";
        ram_buffer(34372) := X"02A01021";
        ram_buffer(34373) := X"24550001";
        ram_buffer(34374) := X"80420000";
        ram_buffer(34375) := X"00000000";
        ram_buffer(34376) := X"0040A021";
        ram_buffer(34377) := X"2683FFE0";
        ram_buffer(34378) := X"2C62005B";
        ram_buffer(34379) := X"1040055B";
        ram_buffer(34380) := X"00000000";
        ram_buffer(34381) := X"00031880";
        ram_buffer(34382) := X"3C02100D";
        ram_buffer(34383) := X"2442A0D8";
        ram_buffer(34384) := X"00621021";
        ram_buffer(34385) := X"8C420000";
        ram_buffer(34386) := X"00000000";
        ram_buffer(34387) := X"00400008";
        ram_buffer(34388) := X"00000000";
        ram_buffer(34389) := X"8FC401E8";
        ram_buffer(34390) := X"0C02BB25";
        ram_buffer(34391) := X"00000000";
        ram_buffer(34392) := X"8C420004";
        ram_buffer(34393) := X"00000000";
        ram_buffer(34394) := X"AFC2003C";
        ram_buffer(34395) := X"8FC4003C";
        ram_buffer(34396) := X"0C02851E";
        ram_buffer(34397) := X"00000000";
        ram_buffer(34398) := X"AFC20040";
        ram_buffer(34399) := X"8FC401E8";
        ram_buffer(34400) := X"0C02BB25";
        ram_buffer(34401) := X"00000000";
        ram_buffer(34402) := X"8C420008";
        ram_buffer(34403) := X"00000000";
        ram_buffer(34404) := X"AFC20044";
        ram_buffer(34405) := X"8FC20040";
        ram_buffer(34406) := X"00000000";
        ram_buffer(34407) := X"1040FFDC";
        ram_buffer(34408) := X"00000000";
        ram_buffer(34409) := X"8FC20044";
        ram_buffer(34410) := X"00000000";
        ram_buffer(34411) := X"1040FFD8";
        ram_buffer(34412) := X"00000000";
        ram_buffer(34413) := X"8FC20044";
        ram_buffer(34414) := X"00000000";
        ram_buffer(34415) := X"80420000";
        ram_buffer(34416) := X"00000000";
        ram_buffer(34417) := X"1040FFD2";
        ram_buffer(34418) := X"00000000";
        ram_buffer(34419) := X"36520400";
        ram_buffer(34420) := X"1000FFCF";
        ram_buffer(34421) := X"00000000";
        ram_buffer(34422) := X"83C20098";
        ram_buffer(34423) := X"00000000";
        ram_buffer(34424) := X"1440FFCB";
        ram_buffer(34425) := X"00000000";
        ram_buffer(34426) := X"24020020";
        ram_buffer(34427) := X"A3C20098";
        ram_buffer(34428) := X"1000FFC7";
        ram_buffer(34429) := X"00000000";
        ram_buffer(34430) := X"36520001";
        ram_buffer(34431) := X"1000FFC4";
        ram_buffer(34432) := X"00000000";
        ram_buffer(34433) := X"8FC301F4";
        ram_buffer(34434) := X"00000000";
        ram_buffer(34435) := X"24620004";
        ram_buffer(34436) := X"AFC201F4";
        ram_buffer(34437) := X"8C620000";
        ram_buffer(34438) := X"00000000";
        ram_buffer(34439) := X"AFC20034";
        ram_buffer(34440) := X"8FC20034";
        ram_buffer(34441) := X"00000000";
        ram_buffer(34442) := X"04400003";
        ram_buffer(34443) := X"00000000";
        ram_buffer(34444) := X"1000FFB7";
        ram_buffer(34445) := X"00000000";
        ram_buffer(34446) := X"8FC20034";
        ram_buffer(34447) := X"00000000";
        ram_buffer(34448) := X"00021023";
        ram_buffer(34449) := X"AFC20034";
        ram_buffer(34450) := X"36520004";
        ram_buffer(34451) := X"1000FFB0";
        ram_buffer(34452) := X"00000000";
        ram_buffer(34453) := X"2402002B";
        ram_buffer(34454) := X"A3C20098";
        ram_buffer(34455) := X"1000FFAC";
        ram_buffer(34456) := X"00000000";
        ram_buffer(34457) := X"02A01021";
        ram_buffer(34458) := X"24550001";
        ram_buffer(34459) := X"80420000";
        ram_buffer(34460) := X"00000000";
        ram_buffer(34461) := X"0040A021";
        ram_buffer(34462) := X"2402002A";
        ram_buffer(34463) := X"16820010";
        ram_buffer(34464) := X"00000000";
        ram_buffer(34465) := X"8FC301F4";
        ram_buffer(34466) := X"00000000";
        ram_buffer(34467) := X"24620004";
        ram_buffer(34468) := X"AFC201F4";
        ram_buffer(34469) := X"8C620000";
        ram_buffer(34470) := X"00000000";
        ram_buffer(34471) := X"AFC20038";
        ram_buffer(34472) := X"8FC20038";
        ram_buffer(34473) := X"00000000";
        ram_buffer(34474) := X"0441FF99";
        ram_buffer(34475) := X"00000000";
        ram_buffer(34476) := X"2402FFFF";
        ram_buffer(34477) := X"AFC20038";
        ram_buffer(34478) := X"1000FF95";
        ram_buffer(34479) := X"00000000";
        ram_buffer(34480) := X"00008821";
        ram_buffer(34481) := X"1000000D";
        ram_buffer(34482) := X"00000000";
        ram_buffer(34483) := X"02201821";
        ram_buffer(34484) := X"00031040";
        ram_buffer(34485) := X"00401821";
        ram_buffer(34486) := X"00031080";
        ram_buffer(34487) := X"00621821";
        ram_buffer(34488) := X"2682FFD0";
        ram_buffer(34489) := X"00628821";
        ram_buffer(34490) := X"02A01021";
        ram_buffer(34491) := X"24550001";
        ram_buffer(34492) := X"80420000";
        ram_buffer(34493) := X"00000000";
        ram_buffer(34494) := X"0040A021";
        ram_buffer(34495) := X"2682FFD0";
        ram_buffer(34496) := X"2C42000A";
        ram_buffer(34497) := X"1440FFF1";
        ram_buffer(34498) := X"00000000";
        ram_buffer(34499) := X"02201021";
        ram_buffer(34500) := X"04410002";
        ram_buffer(34501) := X"00000000";
        ram_buffer(34502) := X"2402FFFF";
        ram_buffer(34503) := X"AFC20038";
        ram_buffer(34504) := X"1000FF80";
        ram_buffer(34505) := X"00000000";
        ram_buffer(34506) := X"36520080";
        ram_buffer(34507) := X"1000FF78";
        ram_buffer(34508) := X"00000000";
        ram_buffer(34509) := X"00008821";
        ram_buffer(34510) := X"02201821";
        ram_buffer(34511) := X"00031040";
        ram_buffer(34512) := X"00401821";
        ram_buffer(34513) := X"00031080";
        ram_buffer(34514) := X"00621821";
        ram_buffer(34515) := X"2682FFD0";
        ram_buffer(34516) := X"00628821";
        ram_buffer(34517) := X"02A01021";
        ram_buffer(34518) := X"24550001";
        ram_buffer(34519) := X"80420000";
        ram_buffer(34520) := X"00000000";
        ram_buffer(34521) := X"0040A021";
        ram_buffer(34522) := X"2682FFD0";
        ram_buffer(34523) := X"2C42000A";
        ram_buffer(34524) := X"1440FFF1";
        ram_buffer(34525) := X"00000000";
        ram_buffer(34526) := X"AFD10034";
        ram_buffer(34527) := X"1000FF69";
        ram_buffer(34528) := X"00000000";
        ram_buffer(34529) := X"36520008";
        ram_buffer(34530) := X"1000FF61";
        ram_buffer(34531) := X"00000000";
        ram_buffer(34532) := X"82A30000";
        ram_buffer(34533) := X"24020068";
        ram_buffer(34534) := X"14620005";
        ram_buffer(34535) := X"00000000";
        ram_buffer(34536) := X"26B50001";
        ram_buffer(34537) := X"36520200";
        ram_buffer(34538) := X"1000FF59";
        ram_buffer(34539) := X"00000000";
        ram_buffer(34540) := X"36520040";
        ram_buffer(34541) := X"1000FF56";
        ram_buffer(34542) := X"00000000";
        ram_buffer(34543) := X"82A30000";
        ram_buffer(34544) := X"2402006C";
        ram_buffer(34545) := X"14620005";
        ram_buffer(34546) := X"00000000";
        ram_buffer(34547) := X"26B50001";
        ram_buffer(34548) := X"36520020";
        ram_buffer(34549) := X"1000FF4E";
        ram_buffer(34550) := X"00000000";
        ram_buffer(34551) := X"36520010";
        ram_buffer(34552) := X"1000FF4B";
        ram_buffer(34553) := X"00000000";
        ram_buffer(34554) := X"36520020";
        ram_buffer(34555) := X"1000FF48";
        ram_buffer(34556) := X"00000000";
        ram_buffer(34557) := X"36520020";
        ram_buffer(34558) := X"1000FF45";
        ram_buffer(34559) := X"00000000";
        ram_buffer(34560) := X"27D30104";
        ram_buffer(34561) := X"8FC301F4";
        ram_buffer(34562) := X"00000000";
        ram_buffer(34563) := X"24620004";
        ram_buffer(34564) := X"AFC201F4";
        ram_buffer(34565) := X"8C620000";
        ram_buffer(34566) := X"00000000";
        ram_buffer(34567) := X"00021600";
        ram_buffer(34568) := X"00021603";
        ram_buffer(34569) := X"A2620000";
        ram_buffer(34570) := X"24020001";
        ram_buffer(34571) := X"AFC2006C";
        ram_buffer(34572) := X"A3C00098";
        ram_buffer(34573) := X"100004A5";
        ram_buffer(34574) := X"00000000";
        ram_buffer(34575) := X"36520010";
        ram_buffer(34576) := X"32420020";
        ram_buffer(34577) := X"1040000E";
        ram_buffer(34578) := X"00000000";
        ram_buffer(34579) := X"8FC201F4";
        ram_buffer(34580) := X"00000000";
        ram_buffer(34581) := X"24430007";
        ram_buffer(34582) := X"2402FFF8";
        ram_buffer(34583) := X"00621024";
        ram_buffer(34584) := X"24430008";
        ram_buffer(34585) := X"AFC301F4";
        ram_buffer(34586) := X"8C430004";
        ram_buffer(34587) := X"8C420000";
        ram_buffer(34588) := X"AFC30174";
        ram_buffer(34589) := X"AFC20170";
        ram_buffer(34590) := X"10000038";
        ram_buffer(34591) := X"00000000";
        ram_buffer(34592) := X"32420010";
        ram_buffer(34593) := X"1040000C";
        ram_buffer(34594) := X"00000000";
        ram_buffer(34595) := X"8FC301F4";
        ram_buffer(34596) := X"00000000";
        ram_buffer(34597) := X"24620004";
        ram_buffer(34598) := X"AFC201F4";
        ram_buffer(34599) := X"8C620000";
        ram_buffer(34600) := X"00000000";
        ram_buffer(34601) := X"AFC20174";
        ram_buffer(34602) := X"000217C3";
        ram_buffer(34603) := X"AFC20170";
        ram_buffer(34604) := X"1000002A";
        ram_buffer(34605) := X"00000000";
        ram_buffer(34606) := X"32420040";
        ram_buffer(34607) := X"1040000E";
        ram_buffer(34608) := X"00000000";
        ram_buffer(34609) := X"8FC301F4";
        ram_buffer(34610) := X"00000000";
        ram_buffer(34611) := X"24620004";
        ram_buffer(34612) := X"AFC201F4";
        ram_buffer(34613) := X"8C620000";
        ram_buffer(34614) := X"00000000";
        ram_buffer(34615) := X"00021400";
        ram_buffer(34616) := X"00021403";
        ram_buffer(34617) := X"AFC20174";
        ram_buffer(34618) := X"000217C3";
        ram_buffer(34619) := X"AFC20170";
        ram_buffer(34620) := X"1000001A";
        ram_buffer(34621) := X"00000000";
        ram_buffer(34622) := X"32420200";
        ram_buffer(34623) := X"1040000E";
        ram_buffer(34624) := X"00000000";
        ram_buffer(34625) := X"8FC301F4";
        ram_buffer(34626) := X"00000000";
        ram_buffer(34627) := X"24620004";
        ram_buffer(34628) := X"AFC201F4";
        ram_buffer(34629) := X"8C620000";
        ram_buffer(34630) := X"00000000";
        ram_buffer(34631) := X"00021600";
        ram_buffer(34632) := X"00021603";
        ram_buffer(34633) := X"AFC20174";
        ram_buffer(34634) := X"000217C3";
        ram_buffer(34635) := X"AFC20170";
        ram_buffer(34636) := X"1000000A";
        ram_buffer(34637) := X"00000000";
        ram_buffer(34638) := X"8FC301F4";
        ram_buffer(34639) := X"00000000";
        ram_buffer(34640) := X"24620004";
        ram_buffer(34641) := X"AFC201F4";
        ram_buffer(34642) := X"8C620000";
        ram_buffer(34643) := X"00000000";
        ram_buffer(34644) := X"AFC20174";
        ram_buffer(34645) := X"000217C3";
        ram_buffer(34646) := X"AFC20170";
        ram_buffer(34647) := X"8FC30174";
        ram_buffer(34648) := X"8FC20170";
        ram_buffer(34649) := X"AFC3005C";
        ram_buffer(34650) := X"AFC20058";
        ram_buffer(34651) := X"8FC3005C";
        ram_buffer(34652) := X"8FC20058";
        ram_buffer(34653) := X"00000000";
        ram_buffer(34654) := X"0441000E";
        ram_buffer(34655) := X"00000000";
        ram_buffer(34656) := X"00001821";
        ram_buffer(34657) := X"00001021";
        ram_buffer(34658) := X"8FC5005C";
        ram_buffer(34659) := X"8FC40058";
        ram_buffer(34660) := X"00653823";
        ram_buffer(34661) := X"0067402B";
        ram_buffer(34662) := X"00443023";
        ram_buffer(34663) := X"00C81023";
        ram_buffer(34664) := X"00403021";
        ram_buffer(34665) := X"AFC7005C";
        ram_buffer(34666) := X"AFC60058";
        ram_buffer(34667) := X"2402002D";
        ram_buffer(34668) := X"A3C20098";
        ram_buffer(34669) := X"24020001";
        ram_buffer(34670) := X"A3C20060";
        ram_buffer(34671) := X"10000344";
        ram_buffer(34672) := X"00000000";
        ram_buffer(34673) := X"32420008";
        ram_buffer(34674) := X"1040000F";
        ram_buffer(34675) := X"00000000";
        ram_buffer(34676) := X"8FC201F4";
        ram_buffer(34677) := X"00000000";
        ram_buffer(34678) := X"24430007";
        ram_buffer(34679) := X"2402FFF8";
        ram_buffer(34680) := X"00621824";
        ram_buffer(34681) := X"24620008";
        ram_buffer(34682) := X"AFC201F4";
        ram_buffer(34683) := X"8C620000";
        ram_buffer(34684) := X"8C630004";
        ram_buffer(34685) := X"00000000";
        ram_buffer(34686) := X"AFC300A4";
        ram_buffer(34687) := X"AFC200A0";
        ram_buffer(34688) := X"1000000D";
        ram_buffer(34689) := X"00000000";
        ram_buffer(34690) := X"8FC201F4";
        ram_buffer(34691) := X"00000000";
        ram_buffer(34692) := X"24430007";
        ram_buffer(34693) := X"2402FFF8";
        ram_buffer(34694) := X"00621824";
        ram_buffer(34695) := X"24620008";
        ram_buffer(34696) := X"AFC201F4";
        ram_buffer(34697) := X"8C620000";
        ram_buffer(34698) := X"8C630004";
        ram_buffer(34699) := X"00000000";
        ram_buffer(34700) := X"AFC300A4";
        ram_buffer(34701) := X"AFC200A0";
        ram_buffer(34702) := X"8FC300A4";
        ram_buffer(34703) := X"8FC200A0";
        ram_buffer(34704) := X"00602821";
        ram_buffer(34705) := X"00402021";
        ram_buffer(34706) := X"0C02CAED";
        ram_buffer(34707) := X"00000000";
        ram_buffer(34708) := X"00401821";
        ram_buffer(34709) := X"24020001";
        ram_buffer(34710) := X"1462001C";
        ram_buffer(34711) := X"00000000";
        ram_buffer(34712) := X"8FC300A4";
        ram_buffer(34713) := X"8FC200A0";
        ram_buffer(34714) := X"00003821";
        ram_buffer(34715) := X"00003021";
        ram_buffer(34716) := X"00602821";
        ram_buffer(34717) := X"00402021";
        ram_buffer(34718) := X"0C0316F7";
        ram_buffer(34719) := X"00000000";
        ram_buffer(34720) := X"04410003";
        ram_buffer(34721) := X"00000000";
        ram_buffer(34722) := X"2402002D";
        ram_buffer(34723) := X"A3C20098";
        ram_buffer(34724) := X"2A820048";
        ram_buffer(34725) := X"10400005";
        ram_buffer(34726) := X"00000000";
        ram_buffer(34727) := X"3C02100D";
        ram_buffer(34728) := X"2453A078";
        ram_buffer(34729) := X"10000003";
        ram_buffer(34730) := X"00000000";
        ram_buffer(34731) := X"3C02100D";
        ram_buffer(34732) := X"2453A07C";
        ram_buffer(34733) := X"24020003";
        ram_buffer(34734) := X"AFC2006C";
        ram_buffer(34735) := X"2402FF7F";
        ram_buffer(34736) := X"02429024";
        ram_buffer(34737) := X"10000401";
        ram_buffer(34738) := X"00000000";
        ram_buffer(34739) := X"8FC300A4";
        ram_buffer(34740) := X"8FC200A0";
        ram_buffer(34741) := X"00602821";
        ram_buffer(34742) := X"00402021";
        ram_buffer(34743) := X"0C02CAED";
        ram_buffer(34744) := X"00000000";
        ram_buffer(34745) := X"14400010";
        ram_buffer(34746) := X"00000000";
        ram_buffer(34747) := X"2A820048";
        ram_buffer(34748) := X"10400005";
        ram_buffer(34749) := X"00000000";
        ram_buffer(34750) := X"3C02100D";
        ram_buffer(34751) := X"2453A080";
        ram_buffer(34752) := X"10000003";
        ram_buffer(34753) := X"00000000";
        ram_buffer(34754) := X"3C02100D";
        ram_buffer(34755) := X"2453A084";
        ram_buffer(34756) := X"24020003";
        ram_buffer(34757) := X"AFC2006C";
        ram_buffer(34758) := X"2402FF7F";
        ram_buffer(34759) := X"02429024";
        ram_buffer(34760) := X"100003EA";
        ram_buffer(34761) := X"00000000";
        ram_buffer(34762) := X"24020061";
        ram_buffer(34763) := X"12820004";
        ram_buffer(34764) := X"00000000";
        ram_buffer(34765) := X"24020041";
        ram_buffer(34766) := X"1682002F";
        ram_buffer(34767) := X"00000000";
        ram_buffer(34768) := X"24020030";
        ram_buffer(34769) := X"A3C20168";
        ram_buffer(34770) := X"24020061";
        ram_buffer(34771) := X"16820004";
        ram_buffer(34772) := X"00000000";
        ram_buffer(34773) := X"24020078";
        ram_buffer(34774) := X"10000002";
        ram_buffer(34775) := X"00000000";
        ram_buffer(34776) := X"24020058";
        ram_buffer(34777) := X"A3C20169";
        ram_buffer(34778) := X"36520002";
        ram_buffer(34779) := X"8FC20038";
        ram_buffer(34780) := X"00000000";
        ram_buffer(34781) := X"28420064";
        ram_buffer(34782) := X"1440001C";
        ram_buffer(34783) := X"00000000";
        ram_buffer(34784) := X"8FC20038";
        ram_buffer(34785) := X"00000000";
        ram_buffer(34786) := X"24420001";
        ram_buffer(34787) := X"00402821";
        ram_buffer(34788) := X"8FC401E8";
        ram_buffer(34789) := X"0C027B8F";
        ram_buffer(34790) := X"00000000";
        ram_buffer(34791) := X"AFC20074";
        ram_buffer(34792) := X"8FC20074";
        ram_buffer(34793) := X"00000000";
        ram_buffer(34794) := X"1440000D";
        ram_buffer(34795) := X"00000000";
        ram_buffer(34796) := X"8FC201EC";
        ram_buffer(34797) := X"00000000";
        ram_buffer(34798) := X"8442000C";
        ram_buffer(34799) := X"00000000";
        ram_buffer(34800) := X"34420040";
        ram_buffer(34801) := X"00021C00";
        ram_buffer(34802) := X"00031C03";
        ram_buffer(34803) := X"8FC201EC";
        ram_buffer(34804) := X"00000000";
        ram_buffer(34805) := X"A443000C";
        ram_buffer(34806) := X"10000A42";
        ram_buffer(34807) := X"00000000";
        ram_buffer(34808) := X"8FD30074";
        ram_buffer(34809) := X"10000018";
        ram_buffer(34810) := X"00000000";
        ram_buffer(34811) := X"27D30104";
        ram_buffer(34812) := X"10000015";
        ram_buffer(34813) := X"00000000";
        ram_buffer(34814) := X"8FC30038";
        ram_buffer(34815) := X"2402FFFF";
        ram_buffer(34816) := X"14620005";
        ram_buffer(34817) := X"00000000";
        ram_buffer(34818) := X"24020006";
        ram_buffer(34819) := X"AFC20038";
        ram_buffer(34820) := X"1000000D";
        ram_buffer(34821) := X"00000000";
        ram_buffer(34822) := X"24020067";
        ram_buffer(34823) := X"12820004";
        ram_buffer(34824) := X"00000000";
        ram_buffer(34825) := X"24020047";
        ram_buffer(34826) := X"16820007";
        ram_buffer(34827) := X"00000000";
        ram_buffer(34828) := X"8FC20038";
        ram_buffer(34829) := X"00000000";
        ram_buffer(34830) := X"14400003";
        ram_buffer(34831) := X"00000000";
        ram_buffer(34832) := X"24020001";
        ram_buffer(34833) := X"AFC20038";
        ram_buffer(34834) := X"36520100";
        ram_buffer(34835) := X"8FC500A4";
        ram_buffer(34836) := X"8FC400A0";
        ram_buffer(34837) := X"AFB30028";
        ram_buffer(34838) := X"27C200B4";
        ram_buffer(34839) := X"AFA20024";
        ram_buffer(34840) := X"AFB40020";
        ram_buffer(34841) := X"27C200A8";
        ram_buffer(34842) := X"AFA2001C";
        ram_buffer(34843) := X"27C20099";
        ram_buffer(34844) := X"AFA20018";
        ram_buffer(34845) := X"AFB20014";
        ram_buffer(34846) := X"8FC20038";
        ram_buffer(34847) := X"00000000";
        ram_buffer(34848) := X"AFA20010";
        ram_buffer(34849) := X"00A03821";
        ram_buffer(34850) := X"00803021";
        ram_buffer(34851) := X"8FC401E8";
        ram_buffer(34852) := X"0C02925C";
        ram_buffer(34853) := X"00000000";
        ram_buffer(34854) := X"00409821";
        ram_buffer(34855) := X"24020067";
        ram_buffer(34856) := X"12820004";
        ram_buffer(34857) := X"00000000";
        ram_buffer(34858) := X"24020047";
        ram_buffer(34859) := X"16820012";
        ram_buffer(34860) := X"00000000";
        ram_buffer(34861) := X"8FC200A8";
        ram_buffer(34862) := X"00000000";
        ram_buffer(34863) := X"2842FFFD";
        ram_buffer(34864) := X"14400007";
        ram_buffer(34865) := X"00000000";
        ram_buffer(34866) := X"8FC300A8";
        ram_buffer(34867) := X"8FC20038";
        ram_buffer(34868) := X"00000000";
        ram_buffer(34869) := X"0043102A";
        ram_buffer(34870) := X"10400004";
        ram_buffer(34871) := X"00000000";
        ram_buffer(34872) := X"2694FFFE";
        ram_buffer(34873) := X"10000008";
        ram_buffer(34874) := X"00000000";
        ram_buffer(34875) := X"24140067";
        ram_buffer(34876) := X"10000005";
        ram_buffer(34877) := X"00000000";
        ram_buffer(34878) := X"24020046";
        ram_buffer(34879) := X"16820002";
        ram_buffer(34880) := X"00000000";
        ram_buffer(34881) := X"24140066";
        ram_buffer(34882) := X"2A820066";
        ram_buffer(34883) := X"10400022";
        ram_buffer(34884) := X"00000000";
        ram_buffer(34885) := X"8FC200A8";
        ram_buffer(34886) := X"00000000";
        ram_buffer(34887) := X"2442FFFF";
        ram_buffer(34888) := X"AFC200A8";
        ram_buffer(34889) := X"8FC300A8";
        ram_buffer(34890) := X"27C200AC";
        ram_buffer(34891) := X"02803021";
        ram_buffer(34892) := X"00602821";
        ram_buffer(34893) := X"00402021";
        ram_buffer(34894) := X"0C0293C2";
        ram_buffer(34895) := X"00000000";
        ram_buffer(34896) := X"AFC20048";
        ram_buffer(34897) := X"8FC300B4";
        ram_buffer(34898) := X"8FC20048";
        ram_buffer(34899) := X"00000000";
        ram_buffer(34900) := X"00431021";
        ram_buffer(34901) := X"AFC2006C";
        ram_buffer(34902) := X"8FC200B4";
        ram_buffer(34903) := X"00000000";
        ram_buffer(34904) := X"28420002";
        ram_buffer(34905) := X"10400004";
        ram_buffer(34906) := X"00000000";
        ram_buffer(34907) := X"32420001";
        ram_buffer(34908) := X"10400005";
        ram_buffer(34909) := X"00000000";
        ram_buffer(34910) := X"8FC2006C";
        ram_buffer(34911) := X"00000000";
        ram_buffer(34912) := X"24420001";
        ram_buffer(34913) := X"AFC2006C";
        ram_buffer(34914) := X"2402FBFF";
        ram_buffer(34915) := X"02429024";
        ram_buffer(34916) := X"1000009D";
        ram_buffer(34917) := X"00000000";
        ram_buffer(34918) := X"24020066";
        ram_buffer(34919) := X"16820028";
        ram_buffer(34920) := X"00000000";
        ram_buffer(34921) := X"8FC200A8";
        ram_buffer(34922) := X"00000000";
        ram_buffer(34923) := X"18400014";
        ram_buffer(34924) := X"00000000";
        ram_buffer(34925) := X"8FC200A8";
        ram_buffer(34926) := X"00000000";
        ram_buffer(34927) := X"AFC2006C";
        ram_buffer(34928) := X"8FC20038";
        ram_buffer(34929) := X"00000000";
        ram_buffer(34930) := X"14400004";
        ram_buffer(34931) := X"00000000";
        ram_buffer(34932) := X"32420001";
        ram_buffer(34933) := X"1040003A";
        ram_buffer(34934) := X"00000000";
        ram_buffer(34935) := X"8FC20038";
        ram_buffer(34936) := X"00000000";
        ram_buffer(34937) := X"24430001";
        ram_buffer(34938) := X"8FC2006C";
        ram_buffer(34939) := X"00000000";
        ram_buffer(34940) := X"00431021";
        ram_buffer(34941) := X"AFC2006C";
        ram_buffer(34942) := X"10000031";
        ram_buffer(34943) := X"00000000";
        ram_buffer(34944) := X"8FC20038";
        ram_buffer(34945) := X"00000000";
        ram_buffer(34946) := X"14400004";
        ram_buffer(34947) := X"00000000";
        ram_buffer(34948) := X"32420001";
        ram_buffer(34949) := X"10400006";
        ram_buffer(34950) := X"00000000";
        ram_buffer(34951) := X"8FC20038";
        ram_buffer(34952) := X"00000000";
        ram_buffer(34953) := X"24420002";
        ram_buffer(34954) := X"10000002";
        ram_buffer(34955) := X"00000000";
        ram_buffer(34956) := X"24020001";
        ram_buffer(34957) := X"AFC2006C";
        ram_buffer(34958) := X"10000021";
        ram_buffer(34959) := X"00000000";
        ram_buffer(34960) := X"8FC300A8";
        ram_buffer(34961) := X"8FC200B4";
        ram_buffer(34962) := X"00000000";
        ram_buffer(34963) := X"0062102A";
        ram_buffer(34964) := X"1440000D";
        ram_buffer(34965) := X"00000000";
        ram_buffer(34966) := X"8FC200A8";
        ram_buffer(34967) := X"00000000";
        ram_buffer(34968) := X"AFC2006C";
        ram_buffer(34969) := X"32420001";
        ram_buffer(34970) := X"10400015";
        ram_buffer(34971) := X"00000000";
        ram_buffer(34972) := X"8FC2006C";
        ram_buffer(34973) := X"00000000";
        ram_buffer(34974) := X"24420001";
        ram_buffer(34975) := X"AFC2006C";
        ram_buffer(34976) := X"1000000F";
        ram_buffer(34977) := X"00000000";
        ram_buffer(34978) := X"8FC200A8";
        ram_buffer(34979) := X"00000000";
        ram_buffer(34980) := X"1C400006";
        ram_buffer(34981) := X"00000000";
        ram_buffer(34982) := X"8FC300A8";
        ram_buffer(34983) := X"24020002";
        ram_buffer(34984) := X"00431823";
        ram_buffer(34985) := X"10000002";
        ram_buffer(34986) := X"00000000";
        ram_buffer(34987) := X"24030001";
        ram_buffer(34988) := X"8FC200B4";
        ram_buffer(34989) := X"00000000";
        ram_buffer(34990) := X"00621021";
        ram_buffer(34991) := X"AFC2006C";
        ram_buffer(34992) := X"32420400";
        ram_buffer(34993) := X"1040004D";
        ram_buffer(34994) := X"00000000";
        ram_buffer(34995) := X"8FC200A8";
        ram_buffer(34996) := X"00000000";
        ram_buffer(34997) := X"18400049";
        ram_buffer(34998) := X"00000000";
        ram_buffer(34999) := X"AFC00054";
        ram_buffer(35000) := X"8FC20054";
        ram_buffer(35001) := X"00000000";
        ram_buffer(35002) := X"AFC20050";
        ram_buffer(35003) := X"8FC200A8";
        ram_buffer(35004) := X"00000000";
        ram_buffer(35005) := X"AFC2004C";
        ram_buffer(35006) := X"10000029";
        ram_buffer(35007) := X"00000000";
        ram_buffer(35008) := X"8FC20044";
        ram_buffer(35009) := X"00000000";
        ram_buffer(35010) := X"80420000";
        ram_buffer(35011) := X"00000000";
        ram_buffer(35012) := X"00401821";
        ram_buffer(35013) := X"8FC2004C";
        ram_buffer(35014) := X"00000000";
        ram_buffer(35015) := X"0062102A";
        ram_buffer(35016) := X"10400027";
        ram_buffer(35017) := X"00000000";
        ram_buffer(35018) := X"8FC20044";
        ram_buffer(35019) := X"00000000";
        ram_buffer(35020) := X"80420000";
        ram_buffer(35021) := X"00000000";
        ram_buffer(35022) := X"00401821";
        ram_buffer(35023) := X"8FC2004C";
        ram_buffer(35024) := X"00000000";
        ram_buffer(35025) := X"00431023";
        ram_buffer(35026) := X"AFC2004C";
        ram_buffer(35027) := X"8FC20044";
        ram_buffer(35028) := X"00000000";
        ram_buffer(35029) := X"24420001";
        ram_buffer(35030) := X"80420000";
        ram_buffer(35031) := X"00000000";
        ram_buffer(35032) := X"1040000B";
        ram_buffer(35033) := X"00000000";
        ram_buffer(35034) := X"8FC20050";
        ram_buffer(35035) := X"00000000";
        ram_buffer(35036) := X"24420001";
        ram_buffer(35037) := X"AFC20050";
        ram_buffer(35038) := X"8FC20044";
        ram_buffer(35039) := X"00000000";
        ram_buffer(35040) := X"24420001";
        ram_buffer(35041) := X"AFC20044";
        ram_buffer(35042) := X"10000005";
        ram_buffer(35043) := X"00000000";
        ram_buffer(35044) := X"8FC20054";
        ram_buffer(35045) := X"00000000";
        ram_buffer(35046) := X"24420001";
        ram_buffer(35047) := X"AFC20054";
        ram_buffer(35048) := X"8FC20044";
        ram_buffer(35049) := X"00000000";
        ram_buffer(35050) := X"80430000";
        ram_buffer(35051) := X"2402007F";
        ram_buffer(35052) := X"1462FFD3";
        ram_buffer(35053) := X"00000000";
        ram_buffer(35054) := X"10000002";
        ram_buffer(35055) := X"00000000";
        ram_buffer(35056) := X"00000000";
        ram_buffer(35057) := X"8FC30050";
        ram_buffer(35058) := X"8FC20054";
        ram_buffer(35059) := X"00000000";
        ram_buffer(35060) := X"00621021";
        ram_buffer(35061) := X"00401821";
        ram_buffer(35062) := X"8FC20040";
        ram_buffer(35063) := X"00000000";
        ram_buffer(35064) := X"00620018";
        ram_buffer(35065) := X"8FC2006C";
        ram_buffer(35066) := X"00001812";
        ram_buffer(35067) := X"00621021";
        ram_buffer(35068) := X"AFC2006C";
        ram_buffer(35069) := X"10000004";
        ram_buffer(35070) := X"00000000";
        ram_buffer(35071) := X"8FC200A8";
        ram_buffer(35072) := X"00000000";
        ram_buffer(35073) := X"AFC2004C";
        ram_buffer(35074) := X"83C20099";
        ram_buffer(35075) := X"00000000";
        ram_buffer(35076) := X"104002AD";
        ram_buffer(35077) := X"00000000";
        ram_buffer(35078) := X"2402002D";
        ram_buffer(35079) := X"A3C20098";
        ram_buffer(35080) := X"100002A9";
        ram_buffer(35081) := X"00000000";
        ram_buffer(35082) := X"32420020";
        ram_buffer(35083) := X"10400011";
        ram_buffer(35084) := X"00000000";
        ram_buffer(35085) := X"8FC201F4";
        ram_buffer(35086) := X"00000000";
        ram_buffer(35087) := X"24430004";
        ram_buffer(35088) := X"AFC301F4";
        ram_buffer(35089) := X"8C430000";
        ram_buffer(35090) := X"8FC20030";
        ram_buffer(35091) := X"00000000";
        ram_buffer(35092) := X"AFC2018C";
        ram_buffer(35093) := X"000217C3";
        ram_buffer(35094) := X"AFC20188";
        ram_buffer(35095) := X"8FC5018C";
        ram_buffer(35096) := X"8FC40188";
        ram_buffer(35097) := X"AC650004";
        ram_buffer(35098) := X"AC640000";
        ram_buffer(35099) := X"1000088E";
        ram_buffer(35100) := X"00000000";
        ram_buffer(35101) := X"32420010";
        ram_buffer(35102) := X"1040000B";
        ram_buffer(35103) := X"00000000";
        ram_buffer(35104) := X"8FC201F4";
        ram_buffer(35105) := X"00000000";
        ram_buffer(35106) := X"24430004";
        ram_buffer(35107) := X"AFC301F4";
        ram_buffer(35108) := X"8C420000";
        ram_buffer(35109) := X"8FC30030";
        ram_buffer(35110) := X"00000000";
        ram_buffer(35111) := X"AC430000";
        ram_buffer(35112) := X"10000881";
        ram_buffer(35113) := X"00000000";
        ram_buffer(35114) := X"32420040";
        ram_buffer(35115) := X"1040000D";
        ram_buffer(35116) := X"00000000";
        ram_buffer(35117) := X"8FC201F4";
        ram_buffer(35118) := X"00000000";
        ram_buffer(35119) := X"24430004";
        ram_buffer(35120) := X"AFC301F4";
        ram_buffer(35121) := X"8C420000";
        ram_buffer(35122) := X"8FC30030";
        ram_buffer(35123) := X"00000000";
        ram_buffer(35124) := X"00031C00";
        ram_buffer(35125) := X"00031C03";
        ram_buffer(35126) := X"A4430000";
        ram_buffer(35127) := X"10000872";
        ram_buffer(35128) := X"00000000";
        ram_buffer(35129) := X"32420200";
        ram_buffer(35130) := X"1040000D";
        ram_buffer(35131) := X"00000000";
        ram_buffer(35132) := X"8FC201F4";
        ram_buffer(35133) := X"00000000";
        ram_buffer(35134) := X"24430004";
        ram_buffer(35135) := X"AFC301F4";
        ram_buffer(35136) := X"8C420000";
        ram_buffer(35137) := X"8FC30030";
        ram_buffer(35138) := X"00000000";
        ram_buffer(35139) := X"00031E00";
        ram_buffer(35140) := X"00031E03";
        ram_buffer(35141) := X"A0430000";
        ram_buffer(35142) := X"10000863";
        ram_buffer(35143) := X"00000000";
        ram_buffer(35144) := X"8FC201F4";
        ram_buffer(35145) := X"00000000";
        ram_buffer(35146) := X"24430004";
        ram_buffer(35147) := X"AFC301F4";
        ram_buffer(35148) := X"8C420000";
        ram_buffer(35149) := X"8FC30030";
        ram_buffer(35150) := X"00000000";
        ram_buffer(35151) := X"AC430000";
        ram_buffer(35152) := X"10000859";
        ram_buffer(35153) := X"00000000";
        ram_buffer(35154) := X"36520010";
        ram_buffer(35155) := X"32420020";
        ram_buffer(35156) := X"1040000C";
        ram_buffer(35157) := X"00000000";
        ram_buffer(35158) := X"8FC201F4";
        ram_buffer(35159) := X"00000000";
        ram_buffer(35160) := X"24430007";
        ram_buffer(35161) := X"2402FFF8";
        ram_buffer(35162) := X"00621024";
        ram_buffer(35163) := X"24430008";
        ram_buffer(35164) := X"AFC301F4";
        ram_buffer(35165) := X"8C570004";
        ram_buffer(35166) := X"8C560000";
        ram_buffer(35167) := X"1000003C";
        ram_buffer(35168) := X"00000000";
        ram_buffer(35169) := X"32420010";
        ram_buffer(35170) := X"1040000B";
        ram_buffer(35171) := X"00000000";
        ram_buffer(35172) := X"8FC301F4";
        ram_buffer(35173) := X"00000000";
        ram_buffer(35174) := X"24620004";
        ram_buffer(35175) := X"AFC201F4";
        ram_buffer(35176) := X"8C620000";
        ram_buffer(35177) := X"00000000";
        ram_buffer(35178) := X"0040B821";
        ram_buffer(35179) := X"0000B021";
        ram_buffer(35180) := X"1000002F";
        ram_buffer(35181) := X"00000000";
        ram_buffer(35182) := X"32420040";
        ram_buffer(35183) := X"10400011";
        ram_buffer(35184) := X"00000000";
        ram_buffer(35185) := X"8FC301F4";
        ram_buffer(35186) := X"00000000";
        ram_buffer(35187) := X"24620004";
        ram_buffer(35188) := X"AFC201F4";
        ram_buffer(35189) := X"8C620000";
        ram_buffer(35190) := X"00000000";
        ram_buffer(35191) := X"AFC20194";
        ram_buffer(35192) := X"AFC00190";
        ram_buffer(35193) := X"8FC30194";
        ram_buffer(35194) := X"8FC20190";
        ram_buffer(35195) := X"00000000";
        ram_buffer(35196) := X"00402021";
        ram_buffer(35197) := X"30960000";
        ram_buffer(35198) := X"3077FFFF";
        ram_buffer(35199) := X"1000001C";
        ram_buffer(35200) := X"00000000";
        ram_buffer(35201) := X"32420200";
        ram_buffer(35202) := X"10400011";
        ram_buffer(35203) := X"00000000";
        ram_buffer(35204) := X"8FC301F4";
        ram_buffer(35205) := X"00000000";
        ram_buffer(35206) := X"24620004";
        ram_buffer(35207) := X"AFC201F4";
        ram_buffer(35208) := X"8C620000";
        ram_buffer(35209) := X"00000000";
        ram_buffer(35210) := X"AFC2019C";
        ram_buffer(35211) := X"AFC00198";
        ram_buffer(35212) := X"8FC3019C";
        ram_buffer(35213) := X"8FC20198";
        ram_buffer(35214) := X"00000000";
        ram_buffer(35215) := X"00402021";
        ram_buffer(35216) := X"30960000";
        ram_buffer(35217) := X"307700FF";
        ram_buffer(35218) := X"10000009";
        ram_buffer(35219) := X"00000000";
        ram_buffer(35220) := X"8FC301F4";
        ram_buffer(35221) := X"00000000";
        ram_buffer(35222) := X"24620004";
        ram_buffer(35223) := X"AFC201F4";
        ram_buffer(35224) := X"8C620000";
        ram_buffer(35225) := X"00000000";
        ram_buffer(35226) := X"0040B821";
        ram_buffer(35227) := X"0000B021";
        ram_buffer(35228) := X"AFD7005C";
        ram_buffer(35229) := X"AFD60058";
        ram_buffer(35230) := X"A3C00060";
        ram_buffer(35231) := X"2402FBFF";
        ram_buffer(35232) := X"02429024";
        ram_buffer(35233) := X"10000111";
        ram_buffer(35234) := X"00000000";
        ram_buffer(35235) := X"8FC201F4";
        ram_buffer(35236) := X"00000000";
        ram_buffer(35237) := X"24430004";
        ram_buffer(35238) := X"AFC301F4";
        ram_buffer(35239) := X"8C420000";
        ram_buffer(35240) := X"00000000";
        ram_buffer(35241) := X"AFC2005C";
        ram_buffer(35242) := X"AFC00058";
        ram_buffer(35243) := X"24020002";
        ram_buffer(35244) := X"A3C20060";
        ram_buffer(35245) := X"3C02100D";
        ram_buffer(35246) := X"2442A088";
        ram_buffer(35247) := X"AFC20070";
        ram_buffer(35248) := X"36520002";
        ram_buffer(35249) := X"24020030";
        ram_buffer(35250) := X"A3C20168";
        ram_buffer(35251) := X"24140078";
        ram_buffer(35252) := X"24020078";
        ram_buffer(35253) := X"A3C20169";
        ram_buffer(35254) := X"100000FC";
        ram_buffer(35255) := X"00000000";
        ram_buffer(35256) := X"8FC301F4";
        ram_buffer(35257) := X"00000000";
        ram_buffer(35258) := X"24620004";
        ram_buffer(35259) := X"AFC201F4";
        ram_buffer(35260) := X"8C730000";
        ram_buffer(35261) := X"A3C00098";
        ram_buffer(35262) := X"1660000D";
        ram_buffer(35263) := X"00000000";
        ram_buffer(35264) := X"3C02100D";
        ram_buffer(35265) := X"2453A09C";
        ram_buffer(35266) := X"8FC20038";
        ram_buffer(35267) := X"00000000";
        ram_buffer(35268) := X"00401821";
        ram_buffer(35269) := X"2C620007";
        ram_buffer(35270) := X"14400002";
        ram_buffer(35271) := X"00000000";
        ram_buffer(35272) := X"24030006";
        ram_buffer(35273) := X"AFC3006C";
        ram_buffer(35274) := X"100001E8";
        ram_buffer(35275) := X"00000000";
        ram_buffer(35276) := X"8FC20038";
        ram_buffer(35277) := X"00000000";
        ram_buffer(35278) := X"04400018";
        ram_buffer(35279) := X"00000000";
        ram_buffer(35280) := X"8FC20038";
        ram_buffer(35281) := X"00000000";
        ram_buffer(35282) := X"00403021";
        ram_buffer(35283) := X"00002821";
        ram_buffer(35284) := X"02602021";
        ram_buffer(35285) := X"0C02BC51";
        ram_buffer(35286) := X"00000000";
        ram_buffer(35287) := X"AFC20090";
        ram_buffer(35288) := X"8FC20090";
        ram_buffer(35289) := X"00000000";
        ram_buffer(35290) := X"10400007";
        ram_buffer(35291) := X"00000000";
        ram_buffer(35292) := X"8FC30090";
        ram_buffer(35293) := X"02601021";
        ram_buffer(35294) := X"00621023";
        ram_buffer(35295) := X"AFC2006C";
        ram_buffer(35296) := X"100001D2";
        ram_buffer(35297) := X"00000000";
        ram_buffer(35298) := X"8FC20038";
        ram_buffer(35299) := X"00000000";
        ram_buffer(35300) := X"AFC2006C";
        ram_buffer(35301) := X"100001CD";
        ram_buffer(35302) := X"00000000";
        ram_buffer(35303) := X"02602021";
        ram_buffer(35304) := X"0C02851E";
        ram_buffer(35305) := X"00000000";
        ram_buffer(35306) := X"AFC2006C";
        ram_buffer(35307) := X"100001C7";
        ram_buffer(35308) := X"00000000";
        ram_buffer(35309) := X"36520010";
        ram_buffer(35310) := X"32420020";
        ram_buffer(35311) := X"1040000E";
        ram_buffer(35312) := X"00000000";
        ram_buffer(35313) := X"8FC201F4";
        ram_buffer(35314) := X"00000000";
        ram_buffer(35315) := X"24430007";
        ram_buffer(35316) := X"2402FFF8";
        ram_buffer(35317) := X"00621024";
        ram_buffer(35318) := X"24430008";
        ram_buffer(35319) := X"AFC301F4";
        ram_buffer(35320) := X"8C430004";
        ram_buffer(35321) := X"8C420000";
        ram_buffer(35322) := X"AFC3017C";
        ram_buffer(35323) := X"AFC20178";
        ram_buffer(35324) := X"10000040";
        ram_buffer(35325) := X"00000000";
        ram_buffer(35326) := X"32420010";
        ram_buffer(35327) := X"1040000B";
        ram_buffer(35328) := X"00000000";
        ram_buffer(35329) := X"8FC301F4";
        ram_buffer(35330) := X"00000000";
        ram_buffer(35331) := X"24620004";
        ram_buffer(35332) := X"AFC201F4";
        ram_buffer(35333) := X"8C620000";
        ram_buffer(35334) := X"00000000";
        ram_buffer(35335) := X"AFC2017C";
        ram_buffer(35336) := X"AFC00178";
        ram_buffer(35337) := X"10000033";
        ram_buffer(35338) := X"00000000";
        ram_buffer(35339) := X"32420040";
        ram_buffer(35340) := X"10400013";
        ram_buffer(35341) := X"00000000";
        ram_buffer(35342) := X"8FC301F4";
        ram_buffer(35343) := X"00000000";
        ram_buffer(35344) := X"24620004";
        ram_buffer(35345) := X"AFC201F4";
        ram_buffer(35346) := X"8C620000";
        ram_buffer(35347) := X"00000000";
        ram_buffer(35348) := X"AFC201A4";
        ram_buffer(35349) := X"AFC001A0";
        ram_buffer(35350) := X"8FC301A4";
        ram_buffer(35351) := X"8FC201A0";
        ram_buffer(35352) := X"00000000";
        ram_buffer(35353) := X"00402021";
        ram_buffer(35354) := X"30840000";
        ram_buffer(35355) := X"AFC40178";
        ram_buffer(35356) := X"3062FFFF";
        ram_buffer(35357) := X"AFC2017C";
        ram_buffer(35358) := X"1000001E";
        ram_buffer(35359) := X"00000000";
        ram_buffer(35360) := X"32420200";
        ram_buffer(35361) := X"10400013";
        ram_buffer(35362) := X"00000000";
        ram_buffer(35363) := X"8FC301F4";
        ram_buffer(35364) := X"00000000";
        ram_buffer(35365) := X"24620004";
        ram_buffer(35366) := X"AFC201F4";
        ram_buffer(35367) := X"8C620000";
        ram_buffer(35368) := X"00000000";
        ram_buffer(35369) := X"AFC201AC";
        ram_buffer(35370) := X"AFC001A8";
        ram_buffer(35371) := X"8FC301AC";
        ram_buffer(35372) := X"8FC201A8";
        ram_buffer(35373) := X"00000000";
        ram_buffer(35374) := X"00402021";
        ram_buffer(35375) := X"30840000";
        ram_buffer(35376) := X"AFC40178";
        ram_buffer(35377) := X"306200FF";
        ram_buffer(35378) := X"AFC2017C";
        ram_buffer(35379) := X"10000009";
        ram_buffer(35380) := X"00000000";
        ram_buffer(35381) := X"8FC301F4";
        ram_buffer(35382) := X"00000000";
        ram_buffer(35383) := X"24620004";
        ram_buffer(35384) := X"AFC201F4";
        ram_buffer(35385) := X"8C620000";
        ram_buffer(35386) := X"00000000";
        ram_buffer(35387) := X"AFC2017C";
        ram_buffer(35388) := X"AFC00178";
        ram_buffer(35389) := X"8FC3017C";
        ram_buffer(35390) := X"8FC20178";
        ram_buffer(35391) := X"AFC3005C";
        ram_buffer(35392) := X"AFC20058";
        ram_buffer(35393) := X"24020001";
        ram_buffer(35394) := X"A3C20060";
        ram_buffer(35395) := X"1000006F";
        ram_buffer(35396) := X"00000000";
        ram_buffer(35397) := X"3C02100D";
        ram_buffer(35398) := X"2442A0A4";
        ram_buffer(35399) := X"AFC20070";
        ram_buffer(35400) := X"10000004";
        ram_buffer(35401) := X"00000000";
        ram_buffer(35402) := X"3C02100D";
        ram_buffer(35403) := X"2442A088";
        ram_buffer(35404) := X"AFC20070";
        ram_buffer(35405) := X"32420020";
        ram_buffer(35406) := X"1040000E";
        ram_buffer(35407) := X"00000000";
        ram_buffer(35408) := X"8FC201F4";
        ram_buffer(35409) := X"00000000";
        ram_buffer(35410) := X"24430007";
        ram_buffer(35411) := X"2402FFF8";
        ram_buffer(35412) := X"00621024";
        ram_buffer(35413) := X"24430008";
        ram_buffer(35414) := X"AFC301F4";
        ram_buffer(35415) := X"8C430004";
        ram_buffer(35416) := X"8C420000";
        ram_buffer(35417) := X"AFC30184";
        ram_buffer(35418) := X"AFC20180";
        ram_buffer(35419) := X"10000040";
        ram_buffer(35420) := X"00000000";
        ram_buffer(35421) := X"32420010";
        ram_buffer(35422) := X"1040000B";
        ram_buffer(35423) := X"00000000";
        ram_buffer(35424) := X"8FC301F4";
        ram_buffer(35425) := X"00000000";
        ram_buffer(35426) := X"24620004";
        ram_buffer(35427) := X"AFC201F4";
        ram_buffer(35428) := X"8C620000";
        ram_buffer(35429) := X"00000000";
        ram_buffer(35430) := X"AFC20184";
        ram_buffer(35431) := X"AFC00180";
        ram_buffer(35432) := X"10000033";
        ram_buffer(35433) := X"00000000";
        ram_buffer(35434) := X"32420040";
        ram_buffer(35435) := X"10400013";
        ram_buffer(35436) := X"00000000";
        ram_buffer(35437) := X"8FC301F4";
        ram_buffer(35438) := X"00000000";
        ram_buffer(35439) := X"24620004";
        ram_buffer(35440) := X"AFC201F4";
        ram_buffer(35441) := X"8C620000";
        ram_buffer(35442) := X"00000000";
        ram_buffer(35443) := X"AFC201B4";
        ram_buffer(35444) := X"AFC001B0";
        ram_buffer(35445) := X"8FC301B4";
        ram_buffer(35446) := X"8FC201B0";
        ram_buffer(35447) := X"00000000";
        ram_buffer(35448) := X"00402021";
        ram_buffer(35449) := X"30840000";
        ram_buffer(35450) := X"AFC40180";
        ram_buffer(35451) := X"3062FFFF";
        ram_buffer(35452) := X"AFC20184";
        ram_buffer(35453) := X"1000001E";
        ram_buffer(35454) := X"00000000";
        ram_buffer(35455) := X"32420200";
        ram_buffer(35456) := X"10400013";
        ram_buffer(35457) := X"00000000";
        ram_buffer(35458) := X"8FC301F4";
        ram_buffer(35459) := X"00000000";
        ram_buffer(35460) := X"24620004";
        ram_buffer(35461) := X"AFC201F4";
        ram_buffer(35462) := X"8C620000";
        ram_buffer(35463) := X"00000000";
        ram_buffer(35464) := X"AFC201BC";
        ram_buffer(35465) := X"AFC001B8";
        ram_buffer(35466) := X"8FC301BC";
        ram_buffer(35467) := X"8FC201B8";
        ram_buffer(35468) := X"00000000";
        ram_buffer(35469) := X"00402021";
        ram_buffer(35470) := X"30840000";
        ram_buffer(35471) := X"AFC40180";
        ram_buffer(35472) := X"306200FF";
        ram_buffer(35473) := X"AFC20184";
        ram_buffer(35474) := X"10000009";
        ram_buffer(35475) := X"00000000";
        ram_buffer(35476) := X"8FC301F4";
        ram_buffer(35477) := X"00000000";
        ram_buffer(35478) := X"24620004";
        ram_buffer(35479) := X"AFC201F4";
        ram_buffer(35480) := X"8C620000";
        ram_buffer(35481) := X"00000000";
        ram_buffer(35482) := X"AFC20184";
        ram_buffer(35483) := X"AFC00180";
        ram_buffer(35484) := X"8FC30184";
        ram_buffer(35485) := X"8FC20180";
        ram_buffer(35486) := X"AFC3005C";
        ram_buffer(35487) := X"AFC20058";
        ram_buffer(35488) := X"24020002";
        ram_buffer(35489) := X"A3C20060";
        ram_buffer(35490) := X"32420001";
        ram_buffer(35491) := X"1040000D";
        ram_buffer(35492) := X"00000000";
        ram_buffer(35493) := X"8FC20058";
        ram_buffer(35494) := X"8FC3005C";
        ram_buffer(35495) := X"00000000";
        ram_buffer(35496) := X"00431025";
        ram_buffer(35497) := X"10400007";
        ram_buffer(35498) := X"00000000";
        ram_buffer(35499) := X"24020030";
        ram_buffer(35500) := X"A3C20168";
        ram_buffer(35501) := X"00141600";
        ram_buffer(35502) := X"00021603";
        ram_buffer(35503) := X"A3C20169";
        ram_buffer(35504) := X"36520002";
        ram_buffer(35505) := X"2402FBFF";
        ram_buffer(35506) := X"02429024";
        ram_buffer(35507) := X"A3C00098";
        ram_buffer(35508) := X"8FC20038";
        ram_buffer(35509) := X"00000000";
        ram_buffer(35510) := X"AFC20064";
        ram_buffer(35511) := X"8FC20064";
        ram_buffer(35512) := X"00000000";
        ram_buffer(35513) := X"04400003";
        ram_buffer(35514) := X"00000000";
        ram_buffer(35515) := X"2402FF7F";
        ram_buffer(35516) := X"02429024";
        ram_buffer(35517) := X"27D30104";
        ram_buffer(35518) := X"26730064";
        ram_buffer(35519) := X"8FC30058";
        ram_buffer(35520) := X"8FC2005C";
        ram_buffer(35521) := X"00000000";
        ram_buffer(35522) := X"00621825";
        ram_buffer(35523) := X"14600005";
        ram_buffer(35524) := X"00000000";
        ram_buffer(35525) := X"8FC20038";
        ram_buffer(35526) := X"00000000";
        ram_buffer(35527) := X"104000CD";
        ram_buffer(35528) := X"00000000";
        ram_buffer(35529) := X"93C30060";
        ram_buffer(35530) := X"24020001";
        ram_buffer(35531) := X"1062002E";
        ram_buffer(35532) := X"00000000";
        ram_buffer(35533) := X"24020002";
        ram_buffer(35534) := X"1062009C";
        ram_buffer(35535) := X"00000000";
        ram_buffer(35536) := X"146000B8";
        ram_buffer(35537) := X"00000000";
        ram_buffer(35538) := X"2673FFFF";
        ram_buffer(35539) := X"93C2005F";
        ram_buffer(35540) := X"00000000";
        ram_buffer(35541) := X"30420007";
        ram_buffer(35542) := X"304200FF";
        ram_buffer(35543) := X"24420030";
        ram_buffer(35544) := X"304200FF";
        ram_buffer(35545) := X"00021600";
        ram_buffer(35546) := X"00021603";
        ram_buffer(35547) := X"A2620000";
        ram_buffer(35548) := X"8FC20058";
        ram_buffer(35549) := X"00000000";
        ram_buffer(35550) := X"00021F40";
        ram_buffer(35551) := X"8FC2005C";
        ram_buffer(35552) := X"00000000";
        ram_buffer(35553) := X"000210C2";
        ram_buffer(35554) := X"00431025";
        ram_buffer(35555) := X"AFC2005C";
        ram_buffer(35556) := X"8FC20058";
        ram_buffer(35557) := X"00000000";
        ram_buffer(35558) := X"000210C2";
        ram_buffer(35559) := X"AFC20058";
        ram_buffer(35560) := X"8FC30058";
        ram_buffer(35561) := X"8FC2005C";
        ram_buffer(35562) := X"00000000";
        ram_buffer(35563) := X"00621825";
        ram_buffer(35564) := X"1460FFE5";
        ram_buffer(35565) := X"00000000";
        ram_buffer(35566) := X"32420001";
        ram_buffer(35567) := X"104000A2";
        ram_buffer(35568) := X"00000000";
        ram_buffer(35569) := X"82630000";
        ram_buffer(35570) := X"24020030";
        ram_buffer(35571) := X"1062009E";
        ram_buffer(35572) := X"00000000";
        ram_buffer(35573) := X"2673FFFF";
        ram_buffer(35574) := X"24020030";
        ram_buffer(35575) := X"A2620000";
        ram_buffer(35576) := X"10000099";
        ram_buffer(35577) := X"00000000";
        ram_buffer(35578) := X"8FC20058";
        ram_buffer(35579) := X"00000000";
        ram_buffer(35580) := X"14400014";
        ram_buffer(35581) := X"00000000";
        ram_buffer(35582) := X"8FC20058";
        ram_buffer(35583) := X"00000000";
        ram_buffer(35584) := X"14400006";
        ram_buffer(35585) := X"00000000";
        ram_buffer(35586) := X"8FC2005C";
        ram_buffer(35587) := X"00000000";
        ram_buffer(35588) := X"2C42000A";
        ram_buffer(35589) := X"1040000B";
        ram_buffer(35590) := X"00000000";
        ram_buffer(35591) := X"2673FFFF";
        ram_buffer(35592) := X"93C2005F";
        ram_buffer(35593) := X"00000000";
        ram_buffer(35594) := X"24420030";
        ram_buffer(35595) := X"304200FF";
        ram_buffer(35596) := X"00021600";
        ram_buffer(35597) := X"00021603";
        ram_buffer(35598) := X"A2620000";
        ram_buffer(35599) := X"10000083";
        ram_buffer(35600) := X"00000000";
        ram_buffer(35601) := X"AFC000B4";
        ram_buffer(35602) := X"2673FFFF";
        ram_buffer(35603) := X"8FC3005C";
        ram_buffer(35604) := X"8FC20058";
        ram_buffer(35605) := X"2407000A";
        ram_buffer(35606) := X"00003021";
        ram_buffer(35607) := X"00602821";
        ram_buffer(35608) := X"00402021";
        ram_buffer(35609) := X"0C030BFE";
        ram_buffer(35610) := X"00000000";
        ram_buffer(35611) := X"306200FF";
        ram_buffer(35612) := X"24420030";
        ram_buffer(35613) := X"304200FF";
        ram_buffer(35614) := X"00021600";
        ram_buffer(35615) := X"00021603";
        ram_buffer(35616) := X"A2620000";
        ram_buffer(35617) := X"8FC200B4";
        ram_buffer(35618) := X"00000000";
        ram_buffer(35619) := X"24420001";
        ram_buffer(35620) := X"AFC200B4";
        ram_buffer(35621) := X"32420400";
        ram_buffer(35622) := X"10400032";
        ram_buffer(35623) := X"00000000";
        ram_buffer(35624) := X"8FC20044";
        ram_buffer(35625) := X"00000000";
        ram_buffer(35626) := X"80420000";
        ram_buffer(35627) := X"00000000";
        ram_buffer(35628) := X"00401821";
        ram_buffer(35629) := X"8FC200B4";
        ram_buffer(35630) := X"00000000";
        ram_buffer(35631) := X"14620029";
        ram_buffer(35632) := X"00000000";
        ram_buffer(35633) := X"8FC20044";
        ram_buffer(35634) := X"00000000";
        ram_buffer(35635) := X"80430000";
        ram_buffer(35636) := X"2402007F";
        ram_buffer(35637) := X"10620023";
        ram_buffer(35638) := X"00000000";
        ram_buffer(35639) := X"8FC20058";
        ram_buffer(35640) := X"00000000";
        ram_buffer(35641) := X"1440000A";
        ram_buffer(35642) := X"00000000";
        ram_buffer(35643) := X"8FC20058";
        ram_buffer(35644) := X"00000000";
        ram_buffer(35645) := X"1440001B";
        ram_buffer(35646) := X"00000000";
        ram_buffer(35647) := X"8FC2005C";
        ram_buffer(35648) := X"00000000";
        ram_buffer(35649) := X"2C42000A";
        ram_buffer(35650) := X"14400016";
        ram_buffer(35651) := X"00000000";
        ram_buffer(35652) := X"8FC20040";
        ram_buffer(35653) := X"00000000";
        ram_buffer(35654) := X"00021023";
        ram_buffer(35655) := X"02629821";
        ram_buffer(35656) := X"8FC60040";
        ram_buffer(35657) := X"8FC5003C";
        ram_buffer(35658) := X"02602021";
        ram_buffer(35659) := X"0C02CCBF";
        ram_buffer(35660) := X"00000000";
        ram_buffer(35661) := X"AFC000B4";
        ram_buffer(35662) := X"8FC20044";
        ram_buffer(35663) := X"00000000";
        ram_buffer(35664) := X"24420001";
        ram_buffer(35665) := X"80420000";
        ram_buffer(35666) := X"00000000";
        ram_buffer(35667) := X"10400005";
        ram_buffer(35668) := X"00000000";
        ram_buffer(35669) := X"8FC20044";
        ram_buffer(35670) := X"00000000";
        ram_buffer(35671) := X"24420001";
        ram_buffer(35672) := X"AFC20044";
        ram_buffer(35673) := X"8FC3005C";
        ram_buffer(35674) := X"8FC20058";
        ram_buffer(35675) := X"2407000A";
        ram_buffer(35676) := X"00003021";
        ram_buffer(35677) := X"00602821";
        ram_buffer(35678) := X"00402021";
        ram_buffer(35679) := X"0C030A67";
        ram_buffer(35680) := X"00000000";
        ram_buffer(35681) := X"AFC3005C";
        ram_buffer(35682) := X"AFC20058";
        ram_buffer(35683) := X"8FC30058";
        ram_buffer(35684) := X"8FC2005C";
        ram_buffer(35685) := X"00000000";
        ram_buffer(35686) := X"00621825";
        ram_buffer(35687) := X"1460FFAA";
        ram_buffer(35688) := X"00000000";
        ram_buffer(35689) := X"10000029";
        ram_buffer(35690) := X"00000000";
        ram_buffer(35691) := X"2673FFFF";
        ram_buffer(35692) := X"8FC2005C";
        ram_buffer(35693) := X"00000000";
        ram_buffer(35694) := X"3043000F";
        ram_buffer(35695) := X"8FC20070";
        ram_buffer(35696) := X"00000000";
        ram_buffer(35697) := X"00431021";
        ram_buffer(35698) := X"80420000";
        ram_buffer(35699) := X"00000000";
        ram_buffer(35700) := X"A2620000";
        ram_buffer(35701) := X"8FC20058";
        ram_buffer(35702) := X"00000000";
        ram_buffer(35703) := X"00021F00";
        ram_buffer(35704) := X"8FC2005C";
        ram_buffer(35705) := X"00000000";
        ram_buffer(35706) := X"00021102";
        ram_buffer(35707) := X"00431025";
        ram_buffer(35708) := X"AFC2005C";
        ram_buffer(35709) := X"8FC20058";
        ram_buffer(35710) := X"00000000";
        ram_buffer(35711) := X"00021102";
        ram_buffer(35712) := X"AFC20058";
        ram_buffer(35713) := X"8FC30058";
        ram_buffer(35714) := X"8FC2005C";
        ram_buffer(35715) := X"00000000";
        ram_buffer(35716) := X"00621825";
        ram_buffer(35717) := X"1460FFE5";
        ram_buffer(35718) := X"00000000";
        ram_buffer(35719) := X"1000000B";
        ram_buffer(35720) := X"00000000";
        ram_buffer(35721) := X"3C02100D";
        ram_buffer(35722) := X"2453A0B8";
        ram_buffer(35723) := X"02602021";
        ram_buffer(35724) := X"0C02851E";
        ram_buffer(35725) := X"00000000";
        ram_buffer(35726) := X"AFC2006C";
        ram_buffer(35727) := X"00000000";
        ram_buffer(35728) := X"10000022";
        ram_buffer(35729) := X"00000000";
        ram_buffer(35730) := X"00000000";
        ram_buffer(35731) := X"1000000B";
        ram_buffer(35732) := X"00000000";
        ram_buffer(35733) := X"93C20060";
        ram_buffer(35734) := X"00000000";
        ram_buffer(35735) := X"14400007";
        ram_buffer(35736) := X"00000000";
        ram_buffer(35737) := X"32420001";
        ram_buffer(35738) := X"10400004";
        ram_buffer(35739) := X"00000000";
        ram_buffer(35740) := X"2673FFFF";
        ram_buffer(35741) := X"24020030";
        ram_buffer(35742) := X"A2620000";
        ram_buffer(35743) := X"27C20104";
        ram_buffer(35744) := X"24420064";
        ram_buffer(35745) := X"00401821";
        ram_buffer(35746) := X"02601021";
        ram_buffer(35747) := X"00621023";
        ram_buffer(35748) := X"AFC2006C";
        ram_buffer(35749) := X"1000000D";
        ram_buffer(35750) := X"00000000";
        ram_buffer(35751) := X"12800607";
        ram_buffer(35752) := X"00000000";
        ram_buffer(35753) := X"27D30104";
        ram_buffer(35754) := X"00141600";
        ram_buffer(35755) := X"00021603";
        ram_buffer(35756) := X"A2620000";
        ram_buffer(35757) := X"24020001";
        ram_buffer(35758) := X"AFC2006C";
        ram_buffer(35759) := X"A3C00098";
        ram_buffer(35760) := X"10000002";
        ram_buffer(35761) := X"00000000";
        ram_buffer(35762) := X"00000000";
        ram_buffer(35763) := X"8FC40064";
        ram_buffer(35764) := X"8FC3006C";
        ram_buffer(35765) := X"00000000";
        ram_buffer(35766) := X"0064102A";
        ram_buffer(35767) := X"10400002";
        ram_buffer(35768) := X"00000000";
        ram_buffer(35769) := X"00801821";
        ram_buffer(35770) := X"AFC30068";
        ram_buffer(35771) := X"83C20098";
        ram_buffer(35772) := X"00000000";
        ram_buffer(35773) := X"10400005";
        ram_buffer(35774) := X"00000000";
        ram_buffer(35775) := X"8FC20068";
        ram_buffer(35776) := X"00000000";
        ram_buffer(35777) := X"24420001";
        ram_buffer(35778) := X"AFC20068";
        ram_buffer(35779) := X"32420002";
        ram_buffer(35780) := X"10400005";
        ram_buffer(35781) := X"00000000";
        ram_buffer(35782) := X"8FC20068";
        ram_buffer(35783) := X"00000000";
        ram_buffer(35784) := X"24420002";
        ram_buffer(35785) := X"AFC20068";
        ram_buffer(35786) := X"32420084";
        ram_buffer(35787) := X"14400045";
        ram_buffer(35788) := X"00000000";
        ram_buffer(35789) := X"8FC30034";
        ram_buffer(35790) := X"8FC20068";
        ram_buffer(35791) := X"00000000";
        ram_buffer(35792) := X"00628823";
        ram_buffer(35793) := X"1A20003F";
        ram_buffer(35794) := X"00000000";
        ram_buffer(35795) := X"1000001E";
        ram_buffer(35796) := X"00000000";
        ram_buffer(35797) := X"3C02100D";
        ram_buffer(35798) := X"2442A244";
        ram_buffer(35799) := X"AE020000";
        ram_buffer(35800) := X"24020010";
        ram_buffer(35801) := X"AE020004";
        ram_buffer(35802) := X"8FC200C0";
        ram_buffer(35803) := X"00000000";
        ram_buffer(35804) := X"24420010";
        ram_buffer(35805) := X"AFC200C0";
        ram_buffer(35806) := X"26100008";
        ram_buffer(35807) := X"8FC200BC";
        ram_buffer(35808) := X"00000000";
        ram_buffer(35809) := X"24420001";
        ram_buffer(35810) := X"AFC200BC";
        ram_buffer(35811) := X"8FC200BC";
        ram_buffer(35812) := X"00000000";
        ram_buffer(35813) := X"28420008";
        ram_buffer(35814) := X"1440000A";
        ram_buffer(35815) := X"00000000";
        ram_buffer(35816) := X"27C200B8";
        ram_buffer(35817) := X"00403021";
        ram_buffer(35818) := X"8FC501EC";
        ram_buffer(35819) := X"8FC401E8";
        ram_buffer(35820) := X"0C02DCA6";
        ram_buffer(35821) := X"00000000";
        ram_buffer(35822) := X"144005D4";
        ram_buffer(35823) := X"00000000";
        ram_buffer(35824) := X"27D000C4";
        ram_buffer(35825) := X"2631FFF0";
        ram_buffer(35826) := X"2A220011";
        ram_buffer(35827) := X"1040FFE1";
        ram_buffer(35828) := X"00000000";
        ram_buffer(35829) := X"3C02100D";
        ram_buffer(35830) := X"2442A244";
        ram_buffer(35831) := X"AE020000";
        ram_buffer(35832) := X"02201021";
        ram_buffer(35833) := X"AE020004";
        ram_buffer(35834) := X"8FC300C0";
        ram_buffer(35835) := X"02201021";
        ram_buffer(35836) := X"00621021";
        ram_buffer(35837) := X"AFC200C0";
        ram_buffer(35838) := X"26100008";
        ram_buffer(35839) := X"8FC200BC";
        ram_buffer(35840) := X"00000000";
        ram_buffer(35841) := X"24420001";
        ram_buffer(35842) := X"AFC200BC";
        ram_buffer(35843) := X"8FC200BC";
        ram_buffer(35844) := X"00000000";
        ram_buffer(35845) := X"28420008";
        ram_buffer(35846) := X"1440000A";
        ram_buffer(35847) := X"00000000";
        ram_buffer(35848) := X"27C200B8";
        ram_buffer(35849) := X"00403021";
        ram_buffer(35850) := X"8FC501EC";
        ram_buffer(35851) := X"8FC401E8";
        ram_buffer(35852) := X"0C02DCA6";
        ram_buffer(35853) := X"00000000";
        ram_buffer(35854) := X"144005B7";
        ram_buffer(35855) := X"00000000";
        ram_buffer(35856) := X"27D000C4";
        ram_buffer(35857) := X"83C20098";
        ram_buffer(35858) := X"00000000";
        ram_buffer(35859) := X"1040001C";
        ram_buffer(35860) := X"00000000";
        ram_buffer(35861) := X"27C20098";
        ram_buffer(35862) := X"AE020000";
        ram_buffer(35863) := X"24020001";
        ram_buffer(35864) := X"AE020004";
        ram_buffer(35865) := X"8FC200C0";
        ram_buffer(35866) := X"00000000";
        ram_buffer(35867) := X"24420001";
        ram_buffer(35868) := X"AFC200C0";
        ram_buffer(35869) := X"26100008";
        ram_buffer(35870) := X"8FC200BC";
        ram_buffer(35871) := X"00000000";
        ram_buffer(35872) := X"24420001";
        ram_buffer(35873) := X"AFC200BC";
        ram_buffer(35874) := X"8FC200BC";
        ram_buffer(35875) := X"00000000";
        ram_buffer(35876) := X"28420008";
        ram_buffer(35877) := X"1440000A";
        ram_buffer(35878) := X"00000000";
        ram_buffer(35879) := X"27C200B8";
        ram_buffer(35880) := X"00403021";
        ram_buffer(35881) := X"8FC501EC";
        ram_buffer(35882) := X"8FC401E8";
        ram_buffer(35883) := X"0C02DCA6";
        ram_buffer(35884) := X"00000000";
        ram_buffer(35885) := X"1440059B";
        ram_buffer(35886) := X"00000000";
        ram_buffer(35887) := X"27D000C4";
        ram_buffer(35888) := X"32420002";
        ram_buffer(35889) := X"1040001C";
        ram_buffer(35890) := X"00000000";
        ram_buffer(35891) := X"27C20168";
        ram_buffer(35892) := X"AE020000";
        ram_buffer(35893) := X"24020002";
        ram_buffer(35894) := X"AE020004";
        ram_buffer(35895) := X"8FC200C0";
        ram_buffer(35896) := X"00000000";
        ram_buffer(35897) := X"24420002";
        ram_buffer(35898) := X"AFC200C0";
        ram_buffer(35899) := X"26100008";
        ram_buffer(35900) := X"8FC200BC";
        ram_buffer(35901) := X"00000000";
        ram_buffer(35902) := X"24420001";
        ram_buffer(35903) := X"AFC200BC";
        ram_buffer(35904) := X"8FC200BC";
        ram_buffer(35905) := X"00000000";
        ram_buffer(35906) := X"28420008";
        ram_buffer(35907) := X"1440000A";
        ram_buffer(35908) := X"00000000";
        ram_buffer(35909) := X"27C200B8";
        ram_buffer(35910) := X"00403021";
        ram_buffer(35911) := X"8FC501EC";
        ram_buffer(35912) := X"8FC401E8";
        ram_buffer(35913) := X"0C02DCA6";
        ram_buffer(35914) := X"00000000";
        ram_buffer(35915) := X"14400580";
        ram_buffer(35916) := X"00000000";
        ram_buffer(35917) := X"27D000C4";
        ram_buffer(35918) := X"32430084";
        ram_buffer(35919) := X"24020080";
        ram_buffer(35920) := X"14620045";
        ram_buffer(35921) := X"00000000";
        ram_buffer(35922) := X"8FC30034";
        ram_buffer(35923) := X"8FC20068";
        ram_buffer(35924) := X"00000000";
        ram_buffer(35925) := X"00628823";
        ram_buffer(35926) := X"1A20003F";
        ram_buffer(35927) := X"00000000";
        ram_buffer(35928) := X"1000001E";
        ram_buffer(35929) := X"00000000";
        ram_buffer(35930) := X"3C02100D";
        ram_buffer(35931) := X"2442A254";
        ram_buffer(35932) := X"AE020000";
        ram_buffer(35933) := X"24020010";
        ram_buffer(35934) := X"AE020004";
        ram_buffer(35935) := X"8FC200C0";
        ram_buffer(35936) := X"00000000";
        ram_buffer(35937) := X"24420010";
        ram_buffer(35938) := X"AFC200C0";
        ram_buffer(35939) := X"26100008";
        ram_buffer(35940) := X"8FC200BC";
        ram_buffer(35941) := X"00000000";
        ram_buffer(35942) := X"24420001";
        ram_buffer(35943) := X"AFC200BC";
        ram_buffer(35944) := X"8FC200BC";
        ram_buffer(35945) := X"00000000";
        ram_buffer(35946) := X"28420008";
        ram_buffer(35947) := X"1440000A";
        ram_buffer(35948) := X"00000000";
        ram_buffer(35949) := X"27C200B8";
        ram_buffer(35950) := X"00403021";
        ram_buffer(35951) := X"8FC501EC";
        ram_buffer(35952) := X"8FC401E8";
        ram_buffer(35953) := X"0C02DCA6";
        ram_buffer(35954) := X"00000000";
        ram_buffer(35955) := X"1440055B";
        ram_buffer(35956) := X"00000000";
        ram_buffer(35957) := X"27D000C4";
        ram_buffer(35958) := X"2631FFF0";
        ram_buffer(35959) := X"2A220011";
        ram_buffer(35960) := X"1040FFE1";
        ram_buffer(35961) := X"00000000";
        ram_buffer(35962) := X"3C02100D";
        ram_buffer(35963) := X"2442A254";
        ram_buffer(35964) := X"AE020000";
        ram_buffer(35965) := X"02201021";
        ram_buffer(35966) := X"AE020004";
        ram_buffer(35967) := X"8FC300C0";
        ram_buffer(35968) := X"02201021";
        ram_buffer(35969) := X"00621021";
        ram_buffer(35970) := X"AFC200C0";
        ram_buffer(35971) := X"26100008";
        ram_buffer(35972) := X"8FC200BC";
        ram_buffer(35973) := X"00000000";
        ram_buffer(35974) := X"24420001";
        ram_buffer(35975) := X"AFC200BC";
        ram_buffer(35976) := X"8FC200BC";
        ram_buffer(35977) := X"00000000";
        ram_buffer(35978) := X"28420008";
        ram_buffer(35979) := X"1440000A";
        ram_buffer(35980) := X"00000000";
        ram_buffer(35981) := X"27C200B8";
        ram_buffer(35982) := X"00403021";
        ram_buffer(35983) := X"8FC501EC";
        ram_buffer(35984) := X"8FC401E8";
        ram_buffer(35985) := X"0C02DCA6";
        ram_buffer(35986) := X"00000000";
        ram_buffer(35987) := X"1440053E";
        ram_buffer(35988) := X"00000000";
        ram_buffer(35989) := X"27D000C4";
        ram_buffer(35990) := X"8FC30064";
        ram_buffer(35991) := X"8FC2006C";
        ram_buffer(35992) := X"00000000";
        ram_buffer(35993) := X"00628823";
        ram_buffer(35994) := X"1A20003F";
        ram_buffer(35995) := X"00000000";
        ram_buffer(35996) := X"1000001E";
        ram_buffer(35997) := X"00000000";
        ram_buffer(35998) := X"3C02100D";
        ram_buffer(35999) := X"2442A254";
        ram_buffer(36000) := X"AE020000";
        ram_buffer(36001) := X"24020010";
        ram_buffer(36002) := X"AE020004";
        ram_buffer(36003) := X"8FC200C0";
        ram_buffer(36004) := X"00000000";
        ram_buffer(36005) := X"24420010";
        ram_buffer(36006) := X"AFC200C0";
        ram_buffer(36007) := X"26100008";
        ram_buffer(36008) := X"8FC200BC";
        ram_buffer(36009) := X"00000000";
        ram_buffer(36010) := X"24420001";
        ram_buffer(36011) := X"AFC200BC";
        ram_buffer(36012) := X"8FC200BC";
        ram_buffer(36013) := X"00000000";
        ram_buffer(36014) := X"28420008";
        ram_buffer(36015) := X"1440000A";
        ram_buffer(36016) := X"00000000";
        ram_buffer(36017) := X"27C200B8";
        ram_buffer(36018) := X"00403021";
        ram_buffer(36019) := X"8FC501EC";
        ram_buffer(36020) := X"8FC401E8";
        ram_buffer(36021) := X"0C02DCA6";
        ram_buffer(36022) := X"00000000";
        ram_buffer(36023) := X"1440051D";
        ram_buffer(36024) := X"00000000";
        ram_buffer(36025) := X"27D000C4";
        ram_buffer(36026) := X"2631FFF0";
        ram_buffer(36027) := X"2A220011";
        ram_buffer(36028) := X"1040FFE1";
        ram_buffer(36029) := X"00000000";
        ram_buffer(36030) := X"3C02100D";
        ram_buffer(36031) := X"2442A254";
        ram_buffer(36032) := X"AE020000";
        ram_buffer(36033) := X"02201021";
        ram_buffer(36034) := X"AE020004";
        ram_buffer(36035) := X"8FC300C0";
        ram_buffer(36036) := X"02201021";
        ram_buffer(36037) := X"00621021";
        ram_buffer(36038) := X"AFC200C0";
        ram_buffer(36039) := X"26100008";
        ram_buffer(36040) := X"8FC200BC";
        ram_buffer(36041) := X"00000000";
        ram_buffer(36042) := X"24420001";
        ram_buffer(36043) := X"AFC200BC";
        ram_buffer(36044) := X"8FC200BC";
        ram_buffer(36045) := X"00000000";
        ram_buffer(36046) := X"28420008";
        ram_buffer(36047) := X"1440000A";
        ram_buffer(36048) := X"00000000";
        ram_buffer(36049) := X"27C200B8";
        ram_buffer(36050) := X"00403021";
        ram_buffer(36051) := X"8FC501EC";
        ram_buffer(36052) := X"8FC401E8";
        ram_buffer(36053) := X"0C02DCA6";
        ram_buffer(36054) := X"00000000";
        ram_buffer(36055) := X"14400500";
        ram_buffer(36056) := X"00000000";
        ram_buffer(36057) := X"27D000C4";
        ram_buffer(36058) := X"32420100";
        ram_buffer(36059) := X"1440001F";
        ram_buffer(36060) := X"00000000";
        ram_buffer(36061) := X"AE130000";
        ram_buffer(36062) := X"8FC2006C";
        ram_buffer(36063) := X"00000000";
        ram_buffer(36064) := X"AE020004";
        ram_buffer(36065) := X"8FC300C0";
        ram_buffer(36066) := X"8FC2006C";
        ram_buffer(36067) := X"00000000";
        ram_buffer(36068) := X"00621021";
        ram_buffer(36069) := X"AFC200C0";
        ram_buffer(36070) := X"26100008";
        ram_buffer(36071) := X"8FC200BC";
        ram_buffer(36072) := X"00000000";
        ram_buffer(36073) := X"24420001";
        ram_buffer(36074) := X"AFC200BC";
        ram_buffer(36075) := X"8FC200BC";
        ram_buffer(36076) := X"00000000";
        ram_buffer(36077) := X"28420008";
        ram_buffer(36078) := X"14400452";
        ram_buffer(36079) := X"00000000";
        ram_buffer(36080) := X"27C200B8";
        ram_buffer(36081) := X"00403021";
        ram_buffer(36082) := X"8FC501EC";
        ram_buffer(36083) := X"8FC401E8";
        ram_buffer(36084) := X"0C02DCA6";
        ram_buffer(36085) := X"00000000";
        ram_buffer(36086) := X"144004E4";
        ram_buffer(36087) := X"00000000";
        ram_buffer(36088) := X"27D000C4";
        ram_buffer(36089) := X"10000447";
        ram_buffer(36090) := X"00000000";
        ram_buffer(36091) := X"2A820066";
        ram_buffer(36092) := X"1440035A";
        ram_buffer(36093) := X"00000000";
        ram_buffer(36094) := X"8FC300A4";
        ram_buffer(36095) := X"8FC200A0";
        ram_buffer(36096) := X"00003821";
        ram_buffer(36097) := X"00003021";
        ram_buffer(36098) := X"00602821";
        ram_buffer(36099) := X"00402021";
        ram_buffer(36100) := X"0C03167F";
        ram_buffer(36101) := X"00000000";
        ram_buffer(36102) := X"14400089";
        ram_buffer(36103) := X"00000000";
        ram_buffer(36104) := X"3C02100D";
        ram_buffer(36105) := X"2442A0D4";
        ram_buffer(36106) := X"AE020000";
        ram_buffer(36107) := X"24020001";
        ram_buffer(36108) := X"AE020004";
        ram_buffer(36109) := X"8FC200C0";
        ram_buffer(36110) := X"00000000";
        ram_buffer(36111) := X"24420001";
        ram_buffer(36112) := X"AFC200C0";
        ram_buffer(36113) := X"26100008";
        ram_buffer(36114) := X"8FC200BC";
        ram_buffer(36115) := X"00000000";
        ram_buffer(36116) := X"24420001";
        ram_buffer(36117) := X"AFC200BC";
        ram_buffer(36118) := X"8FC200BC";
        ram_buffer(36119) := X"00000000";
        ram_buffer(36120) := X"28420008";
        ram_buffer(36121) := X"1440000A";
        ram_buffer(36122) := X"00000000";
        ram_buffer(36123) := X"27C200B8";
        ram_buffer(36124) := X"00403021";
        ram_buffer(36125) := X"8FC501EC";
        ram_buffer(36126) := X"8FC401E8";
        ram_buffer(36127) := X"0C02DCA6";
        ram_buffer(36128) := X"00000000";
        ram_buffer(36129) := X"144004BC";
        ram_buffer(36130) := X"00000000";
        ram_buffer(36131) := X"27D000C4";
        ram_buffer(36132) := X"8FC300A8";
        ram_buffer(36133) := X"8FC200B4";
        ram_buffer(36134) := X"00000000";
        ram_buffer(36135) := X"0062102A";
        ram_buffer(36136) := X"14400004";
        ram_buffer(36137) := X"00000000";
        ram_buffer(36138) := X"32420001";
        ram_buffer(36139) := X"10400415";
        ram_buffer(36140) := X"00000000";
        ram_buffer(36141) := X"8FC20084";
        ram_buffer(36142) := X"00000000";
        ram_buffer(36143) := X"AE020000";
        ram_buffer(36144) := X"8FC20088";
        ram_buffer(36145) := X"00000000";
        ram_buffer(36146) := X"AE020004";
        ram_buffer(36147) := X"8FC300C0";
        ram_buffer(36148) := X"8FC20088";
        ram_buffer(36149) := X"00000000";
        ram_buffer(36150) := X"00621021";
        ram_buffer(36151) := X"AFC200C0";
        ram_buffer(36152) := X"26100008";
        ram_buffer(36153) := X"8FC200BC";
        ram_buffer(36154) := X"00000000";
        ram_buffer(36155) := X"24420001";
        ram_buffer(36156) := X"AFC200BC";
        ram_buffer(36157) := X"8FC200BC";
        ram_buffer(36158) := X"00000000";
        ram_buffer(36159) := X"28420008";
        ram_buffer(36160) := X"1440000A";
        ram_buffer(36161) := X"00000000";
        ram_buffer(36162) := X"27C200B8";
        ram_buffer(36163) := X"00403021";
        ram_buffer(36164) := X"8FC501EC";
        ram_buffer(36165) := X"8FC401E8";
        ram_buffer(36166) := X"0C02DCA6";
        ram_buffer(36167) := X"00000000";
        ram_buffer(36168) := X"14400498";
        ram_buffer(36169) := X"00000000";
        ram_buffer(36170) := X"27D000C4";
        ram_buffer(36171) := X"8FC200B4";
        ram_buffer(36172) := X"00000000";
        ram_buffer(36173) := X"2451FFFF";
        ram_buffer(36174) := X"1A2003F2";
        ram_buffer(36175) := X"00000000";
        ram_buffer(36176) := X"1000001E";
        ram_buffer(36177) := X"00000000";
        ram_buffer(36178) := X"3C02100D";
        ram_buffer(36179) := X"2442A254";
        ram_buffer(36180) := X"AE020000";
        ram_buffer(36181) := X"24020010";
        ram_buffer(36182) := X"AE020004";
        ram_buffer(36183) := X"8FC200C0";
        ram_buffer(36184) := X"00000000";
        ram_buffer(36185) := X"24420010";
        ram_buffer(36186) := X"AFC200C0";
        ram_buffer(36187) := X"26100008";
        ram_buffer(36188) := X"8FC200BC";
        ram_buffer(36189) := X"00000000";
        ram_buffer(36190) := X"24420001";
        ram_buffer(36191) := X"AFC200BC";
        ram_buffer(36192) := X"8FC200BC";
        ram_buffer(36193) := X"00000000";
        ram_buffer(36194) := X"28420008";
        ram_buffer(36195) := X"1440000A";
        ram_buffer(36196) := X"00000000";
        ram_buffer(36197) := X"27C200B8";
        ram_buffer(36198) := X"00403021";
        ram_buffer(36199) := X"8FC501EC";
        ram_buffer(36200) := X"8FC401E8";
        ram_buffer(36201) := X"0C02DCA6";
        ram_buffer(36202) := X"00000000";
        ram_buffer(36203) := X"14400478";
        ram_buffer(36204) := X"00000000";
        ram_buffer(36205) := X"27D000C4";
        ram_buffer(36206) := X"2631FFF0";
        ram_buffer(36207) := X"2A220011";
        ram_buffer(36208) := X"1040FFE1";
        ram_buffer(36209) := X"00000000";
        ram_buffer(36210) := X"3C02100D";
        ram_buffer(36211) := X"2442A254";
        ram_buffer(36212) := X"AE020000";
        ram_buffer(36213) := X"02201021";
        ram_buffer(36214) := X"AE020004";
        ram_buffer(36215) := X"8FC300C0";
        ram_buffer(36216) := X"02201021";
        ram_buffer(36217) := X"00621021";
        ram_buffer(36218) := X"AFC200C0";
        ram_buffer(36219) := X"26100008";
        ram_buffer(36220) := X"8FC200BC";
        ram_buffer(36221) := X"00000000";
        ram_buffer(36222) := X"24420001";
        ram_buffer(36223) := X"AFC200BC";
        ram_buffer(36224) := X"8FC200BC";
        ram_buffer(36225) := X"00000000";
        ram_buffer(36226) := X"28420008";
        ram_buffer(36227) := X"144003BD";
        ram_buffer(36228) := X"00000000";
        ram_buffer(36229) := X"27C200B8";
        ram_buffer(36230) := X"00403021";
        ram_buffer(36231) := X"8FC501EC";
        ram_buffer(36232) := X"8FC401E8";
        ram_buffer(36233) := X"0C02DCA6";
        ram_buffer(36234) := X"00000000";
        ram_buffer(36235) := X"1440045B";
        ram_buffer(36236) := X"00000000";
        ram_buffer(36237) := X"27D000C4";
        ram_buffer(36238) := X"100003B2";
        ram_buffer(36239) := X"00000000";
        ram_buffer(36240) := X"8FC200A8";
        ram_buffer(36241) := X"00000000";
        ram_buffer(36242) := X"1C4000A7";
        ram_buffer(36243) := X"00000000";
        ram_buffer(36244) := X"3C02100D";
        ram_buffer(36245) := X"2442A0D4";
        ram_buffer(36246) := X"AE020000";
        ram_buffer(36247) := X"24020001";
        ram_buffer(36248) := X"AE020004";
        ram_buffer(36249) := X"8FC200C0";
        ram_buffer(36250) := X"00000000";
        ram_buffer(36251) := X"24420001";
        ram_buffer(36252) := X"AFC200C0";
        ram_buffer(36253) := X"26100008";
        ram_buffer(36254) := X"8FC200BC";
        ram_buffer(36255) := X"00000000";
        ram_buffer(36256) := X"24420001";
        ram_buffer(36257) := X"AFC200BC";
        ram_buffer(36258) := X"8FC200BC";
        ram_buffer(36259) := X"00000000";
        ram_buffer(36260) := X"28420008";
        ram_buffer(36261) := X"1440000A";
        ram_buffer(36262) := X"00000000";
        ram_buffer(36263) := X"27C200B8";
        ram_buffer(36264) := X"00403021";
        ram_buffer(36265) := X"8FC501EC";
        ram_buffer(36266) := X"8FC401E8";
        ram_buffer(36267) := X"0C02DCA6";
        ram_buffer(36268) := X"00000000";
        ram_buffer(36269) := X"1440043C";
        ram_buffer(36270) := X"00000000";
        ram_buffer(36271) := X"27D000C4";
        ram_buffer(36272) := X"8FC200A8";
        ram_buffer(36273) := X"00000000";
        ram_buffer(36274) := X"14400008";
        ram_buffer(36275) := X"00000000";
        ram_buffer(36276) := X"8FC200B4";
        ram_buffer(36277) := X"00000000";
        ram_buffer(36278) := X"14400004";
        ram_buffer(36279) := X"00000000";
        ram_buffer(36280) := X"32420001";
        ram_buffer(36281) := X"10400387";
        ram_buffer(36282) := X"00000000";
        ram_buffer(36283) := X"8FC20084";
        ram_buffer(36284) := X"00000000";
        ram_buffer(36285) := X"AE020000";
        ram_buffer(36286) := X"8FC20088";
        ram_buffer(36287) := X"00000000";
        ram_buffer(36288) := X"AE020004";
        ram_buffer(36289) := X"8FC300C0";
        ram_buffer(36290) := X"8FC20088";
        ram_buffer(36291) := X"00000000";
        ram_buffer(36292) := X"00621021";
        ram_buffer(36293) := X"AFC200C0";
        ram_buffer(36294) := X"26100008";
        ram_buffer(36295) := X"8FC200BC";
        ram_buffer(36296) := X"00000000";
        ram_buffer(36297) := X"24420001";
        ram_buffer(36298) := X"AFC200BC";
        ram_buffer(36299) := X"8FC200BC";
        ram_buffer(36300) := X"00000000";
        ram_buffer(36301) := X"28420008";
        ram_buffer(36302) := X"1440000A";
        ram_buffer(36303) := X"00000000";
        ram_buffer(36304) := X"27C200B8";
        ram_buffer(36305) := X"00403021";
        ram_buffer(36306) := X"8FC501EC";
        ram_buffer(36307) := X"8FC401E8";
        ram_buffer(36308) := X"0C02DCA6";
        ram_buffer(36309) := X"00000000";
        ram_buffer(36310) := X"14400416";
        ram_buffer(36311) := X"00000000";
        ram_buffer(36312) := X"27D000C4";
        ram_buffer(36313) := X"8FC200A8";
        ram_buffer(36314) := X"00000000";
        ram_buffer(36315) := X"00028823";
        ram_buffer(36316) := X"1A20003F";
        ram_buffer(36317) := X"00000000";
        ram_buffer(36318) := X"1000001E";
        ram_buffer(36319) := X"00000000";
        ram_buffer(36320) := X"3C02100D";
        ram_buffer(36321) := X"2442A254";
        ram_buffer(36322) := X"AE020000";
        ram_buffer(36323) := X"24020010";
        ram_buffer(36324) := X"AE020004";
        ram_buffer(36325) := X"8FC200C0";
        ram_buffer(36326) := X"00000000";
        ram_buffer(36327) := X"24420010";
        ram_buffer(36328) := X"AFC200C0";
        ram_buffer(36329) := X"26100008";
        ram_buffer(36330) := X"8FC200BC";
        ram_buffer(36331) := X"00000000";
        ram_buffer(36332) := X"24420001";
        ram_buffer(36333) := X"AFC200BC";
        ram_buffer(36334) := X"8FC200BC";
        ram_buffer(36335) := X"00000000";
        ram_buffer(36336) := X"28420008";
        ram_buffer(36337) := X"1440000A";
        ram_buffer(36338) := X"00000000";
        ram_buffer(36339) := X"27C200B8";
        ram_buffer(36340) := X"00403021";
        ram_buffer(36341) := X"8FC501EC";
        ram_buffer(36342) := X"8FC401E8";
        ram_buffer(36343) := X"0C02DCA6";
        ram_buffer(36344) := X"00000000";
        ram_buffer(36345) := X"144003F6";
        ram_buffer(36346) := X"00000000";
        ram_buffer(36347) := X"27D000C4";
        ram_buffer(36348) := X"2631FFF0";
        ram_buffer(36349) := X"2A220011";
        ram_buffer(36350) := X"1040FFE1";
        ram_buffer(36351) := X"00000000";
        ram_buffer(36352) := X"3C02100D";
        ram_buffer(36353) := X"2442A254";
        ram_buffer(36354) := X"AE020000";
        ram_buffer(36355) := X"02201021";
        ram_buffer(36356) := X"AE020004";
        ram_buffer(36357) := X"8FC300C0";
        ram_buffer(36358) := X"02201021";
        ram_buffer(36359) := X"00621021";
        ram_buffer(36360) := X"AFC200C0";
        ram_buffer(36361) := X"26100008";
        ram_buffer(36362) := X"8FC200BC";
        ram_buffer(36363) := X"00000000";
        ram_buffer(36364) := X"24420001";
        ram_buffer(36365) := X"AFC200BC";
        ram_buffer(36366) := X"8FC200BC";
        ram_buffer(36367) := X"00000000";
        ram_buffer(36368) := X"28420008";
        ram_buffer(36369) := X"1440000A";
        ram_buffer(36370) := X"00000000";
        ram_buffer(36371) := X"27C200B8";
        ram_buffer(36372) := X"00403021";
        ram_buffer(36373) := X"8FC501EC";
        ram_buffer(36374) := X"8FC401E8";
        ram_buffer(36375) := X"0C02DCA6";
        ram_buffer(36376) := X"00000000";
        ram_buffer(36377) := X"144003D9";
        ram_buffer(36378) := X"00000000";
        ram_buffer(36379) := X"27D000C4";
        ram_buffer(36380) := X"AE130000";
        ram_buffer(36381) := X"8FC200B4";
        ram_buffer(36382) := X"00000000";
        ram_buffer(36383) := X"AE020004";
        ram_buffer(36384) := X"8FC300C0";
        ram_buffer(36385) := X"8FC200B4";
        ram_buffer(36386) := X"00000000";
        ram_buffer(36387) := X"00621021";
        ram_buffer(36388) := X"AFC200C0";
        ram_buffer(36389) := X"26100008";
        ram_buffer(36390) := X"8FC200BC";
        ram_buffer(36391) := X"00000000";
        ram_buffer(36392) := X"24420001";
        ram_buffer(36393) := X"AFC200BC";
        ram_buffer(36394) := X"8FC200BC";
        ram_buffer(36395) := X"00000000";
        ram_buffer(36396) := X"28420008";
        ram_buffer(36397) := X"14400313";
        ram_buffer(36398) := X"00000000";
        ram_buffer(36399) := X"27C200B8";
        ram_buffer(36400) := X"00403021";
        ram_buffer(36401) := X"8FC501EC";
        ram_buffer(36402) := X"8FC401E8";
        ram_buffer(36403) := X"0C02DCA6";
        ram_buffer(36404) := X"00000000";
        ram_buffer(36405) := X"144003C0";
        ram_buffer(36406) := X"00000000";
        ram_buffer(36407) := X"27D000C4";
        ram_buffer(36408) := X"10000308";
        ram_buffer(36409) := X"00000000";
        ram_buffer(36410) := X"AFD30094";
        ram_buffer(36411) := X"8FC200B4";
        ram_buffer(36412) := X"00000000";
        ram_buffer(36413) := X"00401821";
        ram_buffer(36414) := X"8FC20094";
        ram_buffer(36415) := X"00000000";
        ram_buffer(36416) := X"00431021";
        ram_buffer(36417) := X"00401821";
        ram_buffer(36418) := X"02601021";
        ram_buffer(36419) := X"00621023";
        ram_buffer(36420) := X"AFC20078";
        ram_buffer(36421) := X"8FC30078";
        ram_buffer(36422) := X"8FC2004C";
        ram_buffer(36423) := X"00000000";
        ram_buffer(36424) := X"0043102A";
        ram_buffer(36425) := X"10400004";
        ram_buffer(36426) := X"00000000";
        ram_buffer(36427) := X"8FC2004C";
        ram_buffer(36428) := X"00000000";
        ram_buffer(36429) := X"AFC20078";
        ram_buffer(36430) := X"8FC20078";
        ram_buffer(36431) := X"00000000";
        ram_buffer(36432) := X"1840001D";
        ram_buffer(36433) := X"00000000";
        ram_buffer(36434) := X"AE130000";
        ram_buffer(36435) := X"8FC20078";
        ram_buffer(36436) := X"00000000";
        ram_buffer(36437) := X"AE020004";
        ram_buffer(36438) := X"8FC300C0";
        ram_buffer(36439) := X"8FC20078";
        ram_buffer(36440) := X"00000000";
        ram_buffer(36441) := X"00621021";
        ram_buffer(36442) := X"AFC200C0";
        ram_buffer(36443) := X"26100008";
        ram_buffer(36444) := X"8FC200BC";
        ram_buffer(36445) := X"00000000";
        ram_buffer(36446) := X"24420001";
        ram_buffer(36447) := X"AFC200BC";
        ram_buffer(36448) := X"8FC200BC";
        ram_buffer(36449) := X"00000000";
        ram_buffer(36450) := X"28420008";
        ram_buffer(36451) := X"1440000A";
        ram_buffer(36452) := X"00000000";
        ram_buffer(36453) := X"27C200B8";
        ram_buffer(36454) := X"00403021";
        ram_buffer(36455) := X"8FC501EC";
        ram_buffer(36456) := X"8FC401E8";
        ram_buffer(36457) := X"0C02DCA6";
        ram_buffer(36458) := X"00000000";
        ram_buffer(36459) := X"1440038D";
        ram_buffer(36460) := X"00000000";
        ram_buffer(36461) := X"27D000C4";
        ram_buffer(36462) := X"8FC30078";
        ram_buffer(36463) := X"00000000";
        ram_buffer(36464) := X"04610002";
        ram_buffer(36465) := X"00000000";
        ram_buffer(36466) := X"00001821";
        ram_buffer(36467) := X"8FC2004C";
        ram_buffer(36468) := X"00000000";
        ram_buffer(36469) := X"00431023";
        ram_buffer(36470) := X"AFC20078";
        ram_buffer(36471) := X"8FC20078";
        ram_buffer(36472) := X"00000000";
        ram_buffer(36473) := X"18400046";
        ram_buffer(36474) := X"00000000";
        ram_buffer(36475) := X"10000021";
        ram_buffer(36476) := X"00000000";
        ram_buffer(36477) := X"3C02100D";
        ram_buffer(36478) := X"2442A254";
        ram_buffer(36479) := X"AE020000";
        ram_buffer(36480) := X"24020010";
        ram_buffer(36481) := X"AE020004";
        ram_buffer(36482) := X"8FC200C0";
        ram_buffer(36483) := X"00000000";
        ram_buffer(36484) := X"24420010";
        ram_buffer(36485) := X"AFC200C0";
        ram_buffer(36486) := X"26100008";
        ram_buffer(36487) := X"8FC200BC";
        ram_buffer(36488) := X"00000000";
        ram_buffer(36489) := X"24420001";
        ram_buffer(36490) := X"AFC200BC";
        ram_buffer(36491) := X"8FC200BC";
        ram_buffer(36492) := X"00000000";
        ram_buffer(36493) := X"28420008";
        ram_buffer(36494) := X"1440000A";
        ram_buffer(36495) := X"00000000";
        ram_buffer(36496) := X"27C200B8";
        ram_buffer(36497) := X"00403021";
        ram_buffer(36498) := X"8FC501EC";
        ram_buffer(36499) := X"8FC401E8";
        ram_buffer(36500) := X"0C02DCA6";
        ram_buffer(36501) := X"00000000";
        ram_buffer(36502) := X"14400365";
        ram_buffer(36503) := X"00000000";
        ram_buffer(36504) := X"27D000C4";
        ram_buffer(36505) := X"8FC20078";
        ram_buffer(36506) := X"00000000";
        ram_buffer(36507) := X"2442FFF0";
        ram_buffer(36508) := X"AFC20078";
        ram_buffer(36509) := X"8FC20078";
        ram_buffer(36510) := X"00000000";
        ram_buffer(36511) := X"28420011";
        ram_buffer(36512) := X"1040FFDC";
        ram_buffer(36513) := X"00000000";
        ram_buffer(36514) := X"3C02100D";
        ram_buffer(36515) := X"2442A254";
        ram_buffer(36516) := X"AE020000";
        ram_buffer(36517) := X"8FC20078";
        ram_buffer(36518) := X"00000000";
        ram_buffer(36519) := X"AE020004";
        ram_buffer(36520) := X"8FC300C0";
        ram_buffer(36521) := X"8FC20078";
        ram_buffer(36522) := X"00000000";
        ram_buffer(36523) := X"00621021";
        ram_buffer(36524) := X"AFC200C0";
        ram_buffer(36525) := X"26100008";
        ram_buffer(36526) := X"8FC200BC";
        ram_buffer(36527) := X"00000000";
        ram_buffer(36528) := X"24420001";
        ram_buffer(36529) := X"AFC200BC";
        ram_buffer(36530) := X"8FC200BC";
        ram_buffer(36531) := X"00000000";
        ram_buffer(36532) := X"28420008";
        ram_buffer(36533) := X"1440000A";
        ram_buffer(36534) := X"00000000";
        ram_buffer(36535) := X"27C200B8";
        ram_buffer(36536) := X"00403021";
        ram_buffer(36537) := X"8FC501EC";
        ram_buffer(36538) := X"8FC401E8";
        ram_buffer(36539) := X"0C02DCA6";
        ram_buffer(36540) := X"00000000";
        ram_buffer(36541) := X"14400341";
        ram_buffer(36542) := X"00000000";
        ram_buffer(36543) := X"27D000C4";
        ram_buffer(36544) := X"8FC2004C";
        ram_buffer(36545) := X"00000000";
        ram_buffer(36546) := X"02629821";
        ram_buffer(36547) := X"32420400";
        ram_buffer(36548) := X"104000DD";
        ram_buffer(36549) := X"00000000";
        ram_buffer(36550) := X"100000C4";
        ram_buffer(36551) := X"00000000";
        ram_buffer(36552) := X"8FC20054";
        ram_buffer(36553) := X"00000000";
        ram_buffer(36554) := X"18400007";
        ram_buffer(36555) := X"00000000";
        ram_buffer(36556) := X"8FC20054";
        ram_buffer(36557) := X"00000000";
        ram_buffer(36558) := X"2442FFFF";
        ram_buffer(36559) := X"AFC20054";
        ram_buffer(36560) := X"10000009";
        ram_buffer(36561) := X"00000000";
        ram_buffer(36562) := X"8FC20044";
        ram_buffer(36563) := X"00000000";
        ram_buffer(36564) := X"2442FFFF";
        ram_buffer(36565) := X"AFC20044";
        ram_buffer(36566) := X"8FC20050";
        ram_buffer(36567) := X"00000000";
        ram_buffer(36568) := X"2442FFFF";
        ram_buffer(36569) := X"AFC20050";
        ram_buffer(36570) := X"8FC2003C";
        ram_buffer(36571) := X"00000000";
        ram_buffer(36572) := X"AE020000";
        ram_buffer(36573) := X"8FC20040";
        ram_buffer(36574) := X"00000000";
        ram_buffer(36575) := X"AE020004";
        ram_buffer(36576) := X"8FC300C0";
        ram_buffer(36577) := X"8FC20040";
        ram_buffer(36578) := X"00000000";
        ram_buffer(36579) := X"00621021";
        ram_buffer(36580) := X"AFC200C0";
        ram_buffer(36581) := X"26100008";
        ram_buffer(36582) := X"8FC200BC";
        ram_buffer(36583) := X"00000000";
        ram_buffer(36584) := X"24420001";
        ram_buffer(36585) := X"AFC200BC";
        ram_buffer(36586) := X"8FC200BC";
        ram_buffer(36587) := X"00000000";
        ram_buffer(36588) := X"28420008";
        ram_buffer(36589) := X"1440000A";
        ram_buffer(36590) := X"00000000";
        ram_buffer(36591) := X"27C200B8";
        ram_buffer(36592) := X"00403021";
        ram_buffer(36593) := X"8FC501EC";
        ram_buffer(36594) := X"8FC401E8";
        ram_buffer(36595) := X"0C02DCA6";
        ram_buffer(36596) := X"00000000";
        ram_buffer(36597) := X"1440030C";
        ram_buffer(36598) := X"00000000";
        ram_buffer(36599) := X"27D000C4";
        ram_buffer(36600) := X"8FC200B4";
        ram_buffer(36601) := X"00000000";
        ram_buffer(36602) := X"00401821";
        ram_buffer(36603) := X"8FC20094";
        ram_buffer(36604) := X"00000000";
        ram_buffer(36605) := X"00431021";
        ram_buffer(36606) := X"00401821";
        ram_buffer(36607) := X"02601021";
        ram_buffer(36608) := X"00621023";
        ram_buffer(36609) := X"AFC2007C";
        ram_buffer(36610) := X"8FC20044";
        ram_buffer(36611) := X"00000000";
        ram_buffer(36612) := X"80420000";
        ram_buffer(36613) := X"00000000";
        ram_buffer(36614) := X"00401821";
        ram_buffer(36615) := X"8FC2007C";
        ram_buffer(36616) := X"00000000";
        ram_buffer(36617) := X"0062102A";
        ram_buffer(36618) := X"10400006";
        ram_buffer(36619) := X"00000000";
        ram_buffer(36620) := X"8FC20044";
        ram_buffer(36621) := X"00000000";
        ram_buffer(36622) := X"80420000";
        ram_buffer(36623) := X"00000000";
        ram_buffer(36624) := X"AFC2007C";
        ram_buffer(36625) := X"8FC2007C";
        ram_buffer(36626) := X"00000000";
        ram_buffer(36627) := X"1840001D";
        ram_buffer(36628) := X"00000000";
        ram_buffer(36629) := X"AE130000";
        ram_buffer(36630) := X"8FC2007C";
        ram_buffer(36631) := X"00000000";
        ram_buffer(36632) := X"AE020004";
        ram_buffer(36633) := X"8FC300C0";
        ram_buffer(36634) := X"8FC2007C";
        ram_buffer(36635) := X"00000000";
        ram_buffer(36636) := X"00621021";
        ram_buffer(36637) := X"AFC200C0";
        ram_buffer(36638) := X"26100008";
        ram_buffer(36639) := X"8FC200BC";
        ram_buffer(36640) := X"00000000";
        ram_buffer(36641) := X"24420001";
        ram_buffer(36642) := X"AFC200BC";
        ram_buffer(36643) := X"8FC200BC";
        ram_buffer(36644) := X"00000000";
        ram_buffer(36645) := X"28420008";
        ram_buffer(36646) := X"1440000A";
        ram_buffer(36647) := X"00000000";
        ram_buffer(36648) := X"27C200B8";
        ram_buffer(36649) := X"00403021";
        ram_buffer(36650) := X"8FC501EC";
        ram_buffer(36651) := X"8FC401E8";
        ram_buffer(36652) := X"0C02DCA6";
        ram_buffer(36653) := X"00000000";
        ram_buffer(36654) := X"144002D6";
        ram_buffer(36655) := X"00000000";
        ram_buffer(36656) := X"27D000C4";
        ram_buffer(36657) := X"8FC20044";
        ram_buffer(36658) := X"00000000";
        ram_buffer(36659) := X"80420000";
        ram_buffer(36660) := X"00000000";
        ram_buffer(36661) := X"00401821";
        ram_buffer(36662) := X"8FC2007C";
        ram_buffer(36663) := X"00000000";
        ram_buffer(36664) := X"04410002";
        ram_buffer(36665) := X"00000000";
        ram_buffer(36666) := X"00001021";
        ram_buffer(36667) := X"00621023";
        ram_buffer(36668) := X"AFC2007C";
        ram_buffer(36669) := X"8FC2007C";
        ram_buffer(36670) := X"00000000";
        ram_buffer(36671) := X"18400046";
        ram_buffer(36672) := X"00000000";
        ram_buffer(36673) := X"10000021";
        ram_buffer(36674) := X"00000000";
        ram_buffer(36675) := X"3C02100D";
        ram_buffer(36676) := X"2442A254";
        ram_buffer(36677) := X"AE020000";
        ram_buffer(36678) := X"24020010";
        ram_buffer(36679) := X"AE020004";
        ram_buffer(36680) := X"8FC200C0";
        ram_buffer(36681) := X"00000000";
        ram_buffer(36682) := X"24420010";
        ram_buffer(36683) := X"AFC200C0";
        ram_buffer(36684) := X"26100008";
        ram_buffer(36685) := X"8FC200BC";
        ram_buffer(36686) := X"00000000";
        ram_buffer(36687) := X"24420001";
        ram_buffer(36688) := X"AFC200BC";
        ram_buffer(36689) := X"8FC200BC";
        ram_buffer(36690) := X"00000000";
        ram_buffer(36691) := X"28420008";
        ram_buffer(36692) := X"1440000A";
        ram_buffer(36693) := X"00000000";
        ram_buffer(36694) := X"27C200B8";
        ram_buffer(36695) := X"00403021";
        ram_buffer(36696) := X"8FC501EC";
        ram_buffer(36697) := X"8FC401E8";
        ram_buffer(36698) := X"0C02DCA6";
        ram_buffer(36699) := X"00000000";
        ram_buffer(36700) := X"144002AB";
        ram_buffer(36701) := X"00000000";
        ram_buffer(36702) := X"27D000C4";
        ram_buffer(36703) := X"8FC2007C";
        ram_buffer(36704) := X"00000000";
        ram_buffer(36705) := X"2442FFF0";
        ram_buffer(36706) := X"AFC2007C";
        ram_buffer(36707) := X"8FC2007C";
        ram_buffer(36708) := X"00000000";
        ram_buffer(36709) := X"28420011";
        ram_buffer(36710) := X"1040FFDC";
        ram_buffer(36711) := X"00000000";
        ram_buffer(36712) := X"3C02100D";
        ram_buffer(36713) := X"2442A254";
        ram_buffer(36714) := X"AE020000";
        ram_buffer(36715) := X"8FC2007C";
        ram_buffer(36716) := X"00000000";
        ram_buffer(36717) := X"AE020004";
        ram_buffer(36718) := X"8FC300C0";
        ram_buffer(36719) := X"8FC2007C";
        ram_buffer(36720) := X"00000000";
        ram_buffer(36721) := X"00621021";
        ram_buffer(36722) := X"AFC200C0";
        ram_buffer(36723) := X"26100008";
        ram_buffer(36724) := X"8FC200BC";
        ram_buffer(36725) := X"00000000";
        ram_buffer(36726) := X"24420001";
        ram_buffer(36727) := X"AFC200BC";
        ram_buffer(36728) := X"8FC200BC";
        ram_buffer(36729) := X"00000000";
        ram_buffer(36730) := X"28420008";
        ram_buffer(36731) := X"1440000A";
        ram_buffer(36732) := X"00000000";
        ram_buffer(36733) := X"27C200B8";
        ram_buffer(36734) := X"00403021";
        ram_buffer(36735) := X"8FC501EC";
        ram_buffer(36736) := X"8FC401E8";
        ram_buffer(36737) := X"0C02DCA6";
        ram_buffer(36738) := X"00000000";
        ram_buffer(36739) := X"14400287";
        ram_buffer(36740) := X"00000000";
        ram_buffer(36741) := X"27D000C4";
        ram_buffer(36742) := X"8FC20044";
        ram_buffer(36743) := X"00000000";
        ram_buffer(36744) := X"80420000";
        ram_buffer(36745) := X"00000000";
        ram_buffer(36746) := X"02629821";
        ram_buffer(36747) := X"8FC20050";
        ram_buffer(36748) := X"00000000";
        ram_buffer(36749) := X"1C40FF3A";
        ram_buffer(36750) := X"00000000";
        ram_buffer(36751) := X"8FC20054";
        ram_buffer(36752) := X"00000000";
        ram_buffer(36753) := X"1C40FF36";
        ram_buffer(36754) := X"00000000";
        ram_buffer(36755) := X"8FC200B4";
        ram_buffer(36756) := X"00000000";
        ram_buffer(36757) := X"00401821";
        ram_buffer(36758) := X"8FC20094";
        ram_buffer(36759) := X"00000000";
        ram_buffer(36760) := X"00431021";
        ram_buffer(36761) := X"0053102B";
        ram_buffer(36762) := X"10400007";
        ram_buffer(36763) := X"00000000";
        ram_buffer(36764) := X"8FC200B4";
        ram_buffer(36765) := X"00000000";
        ram_buffer(36766) := X"00401821";
        ram_buffer(36767) := X"8FC20094";
        ram_buffer(36768) := X"00000000";
        ram_buffer(36769) := X"00439821";
        ram_buffer(36770) := X"8FC300A8";
        ram_buffer(36771) := X"8FC200B4";
        ram_buffer(36772) := X"00000000";
        ram_buffer(36773) := X"0062102A";
        ram_buffer(36774) := X"14400004";
        ram_buffer(36775) := X"00000000";
        ram_buffer(36776) := X"32420001";
        ram_buffer(36777) := X"1040001F";
        ram_buffer(36778) := X"00000000";
        ram_buffer(36779) := X"8FC20084";
        ram_buffer(36780) := X"00000000";
        ram_buffer(36781) := X"AE020000";
        ram_buffer(36782) := X"8FC20088";
        ram_buffer(36783) := X"00000000";
        ram_buffer(36784) := X"AE020004";
        ram_buffer(36785) := X"8FC300C0";
        ram_buffer(36786) := X"8FC20088";
        ram_buffer(36787) := X"00000000";
        ram_buffer(36788) := X"00621021";
        ram_buffer(36789) := X"AFC200C0";
        ram_buffer(36790) := X"26100008";
        ram_buffer(36791) := X"8FC200BC";
        ram_buffer(36792) := X"00000000";
        ram_buffer(36793) := X"24420001";
        ram_buffer(36794) := X"AFC200BC";
        ram_buffer(36795) := X"8FC200BC";
        ram_buffer(36796) := X"00000000";
        ram_buffer(36797) := X"28420008";
        ram_buffer(36798) := X"1440000A";
        ram_buffer(36799) := X"00000000";
        ram_buffer(36800) := X"27C200B8";
        ram_buffer(36801) := X"00403021";
        ram_buffer(36802) := X"8FC501EC";
        ram_buffer(36803) := X"8FC401E8";
        ram_buffer(36804) := X"0C02DCA6";
        ram_buffer(36805) := X"00000000";
        ram_buffer(36806) := X"14400247";
        ram_buffer(36807) := X"00000000";
        ram_buffer(36808) := X"27D000C4";
        ram_buffer(36809) := X"8FC200B4";
        ram_buffer(36810) := X"00000000";
        ram_buffer(36811) := X"00401821";
        ram_buffer(36812) := X"8FC20094";
        ram_buffer(36813) := X"00000000";
        ram_buffer(36814) := X"00431021";
        ram_buffer(36815) := X"00401821";
        ram_buffer(36816) := X"02601021";
        ram_buffer(36817) := X"00621023";
        ram_buffer(36818) := X"AFC20080";
        ram_buffer(36819) := X"8FC300B4";
        ram_buffer(36820) := X"8FC200A8";
        ram_buffer(36821) := X"00000000";
        ram_buffer(36822) := X"00621823";
        ram_buffer(36823) := X"8FC20080";
        ram_buffer(36824) := X"00000000";
        ram_buffer(36825) := X"0062102A";
        ram_buffer(36826) := X"10400006";
        ram_buffer(36827) := X"00000000";
        ram_buffer(36828) := X"8FC300B4";
        ram_buffer(36829) := X"8FC200A8";
        ram_buffer(36830) := X"00000000";
        ram_buffer(36831) := X"00621023";
        ram_buffer(36832) := X"AFC20080";
        ram_buffer(36833) := X"8FC20080";
        ram_buffer(36834) := X"00000000";
        ram_buffer(36835) := X"1840001D";
        ram_buffer(36836) := X"00000000";
        ram_buffer(36837) := X"AE130000";
        ram_buffer(36838) := X"8FC20080";
        ram_buffer(36839) := X"00000000";
        ram_buffer(36840) := X"AE020004";
        ram_buffer(36841) := X"8FC300C0";
        ram_buffer(36842) := X"8FC20080";
        ram_buffer(36843) := X"00000000";
        ram_buffer(36844) := X"00621021";
        ram_buffer(36845) := X"AFC200C0";
        ram_buffer(36846) := X"26100008";
        ram_buffer(36847) := X"8FC200BC";
        ram_buffer(36848) := X"00000000";
        ram_buffer(36849) := X"24420001";
        ram_buffer(36850) := X"AFC200BC";
        ram_buffer(36851) := X"8FC200BC";
        ram_buffer(36852) := X"00000000";
        ram_buffer(36853) := X"28420008";
        ram_buffer(36854) := X"1440000A";
        ram_buffer(36855) := X"00000000";
        ram_buffer(36856) := X"27C200B8";
        ram_buffer(36857) := X"00403021";
        ram_buffer(36858) := X"8FC501EC";
        ram_buffer(36859) := X"8FC401E8";
        ram_buffer(36860) := X"0C02DCA6";
        ram_buffer(36861) := X"00000000";
        ram_buffer(36862) := X"14400212";
        ram_buffer(36863) := X"00000000";
        ram_buffer(36864) := X"27D000C4";
        ram_buffer(36865) := X"8FC300B4";
        ram_buffer(36866) := X"8FC200A8";
        ram_buffer(36867) := X"00000000";
        ram_buffer(36868) := X"00621823";
        ram_buffer(36869) := X"8FC20080";
        ram_buffer(36870) := X"00000000";
        ram_buffer(36871) := X"04410002";
        ram_buffer(36872) := X"00000000";
        ram_buffer(36873) := X"00001021";
        ram_buffer(36874) := X"00621023";
        ram_buffer(36875) := X"AFC20080";
        ram_buffer(36876) := X"8FC20080";
        ram_buffer(36877) := X"00000000";
        ram_buffer(36878) := X"18400132";
        ram_buffer(36879) := X"00000000";
        ram_buffer(36880) := X"10000021";
        ram_buffer(36881) := X"00000000";
        ram_buffer(36882) := X"3C02100D";
        ram_buffer(36883) := X"2442A254";
        ram_buffer(36884) := X"AE020000";
        ram_buffer(36885) := X"24020010";
        ram_buffer(36886) := X"AE020004";
        ram_buffer(36887) := X"8FC200C0";
        ram_buffer(36888) := X"00000000";
        ram_buffer(36889) := X"24420010";
        ram_buffer(36890) := X"AFC200C0";
        ram_buffer(36891) := X"26100008";
        ram_buffer(36892) := X"8FC200BC";
        ram_buffer(36893) := X"00000000";
        ram_buffer(36894) := X"24420001";
        ram_buffer(36895) := X"AFC200BC";
        ram_buffer(36896) := X"8FC200BC";
        ram_buffer(36897) := X"00000000";
        ram_buffer(36898) := X"28420008";
        ram_buffer(36899) := X"1440000A";
        ram_buffer(36900) := X"00000000";
        ram_buffer(36901) := X"27C200B8";
        ram_buffer(36902) := X"00403021";
        ram_buffer(36903) := X"8FC501EC";
        ram_buffer(36904) := X"8FC401E8";
        ram_buffer(36905) := X"0C02DCA6";
        ram_buffer(36906) := X"00000000";
        ram_buffer(36907) := X"144001E8";
        ram_buffer(36908) := X"00000000";
        ram_buffer(36909) := X"27D000C4";
        ram_buffer(36910) := X"8FC20080";
        ram_buffer(36911) := X"00000000";
        ram_buffer(36912) := X"2442FFF0";
        ram_buffer(36913) := X"AFC20080";
        ram_buffer(36914) := X"8FC20080";
        ram_buffer(36915) := X"00000000";
        ram_buffer(36916) := X"28420011";
        ram_buffer(36917) := X"1040FFDC";
        ram_buffer(36918) := X"00000000";
        ram_buffer(36919) := X"3C02100D";
        ram_buffer(36920) := X"2442A254";
        ram_buffer(36921) := X"AE020000";
        ram_buffer(36922) := X"8FC20080";
        ram_buffer(36923) := X"00000000";
        ram_buffer(36924) := X"AE020004";
        ram_buffer(36925) := X"8FC300C0";
        ram_buffer(36926) := X"8FC20080";
        ram_buffer(36927) := X"00000000";
        ram_buffer(36928) := X"00621021";
        ram_buffer(36929) := X"AFC200C0";
        ram_buffer(36930) := X"26100008";
        ram_buffer(36931) := X"8FC200BC";
        ram_buffer(36932) := X"00000000";
        ram_buffer(36933) := X"24420001";
        ram_buffer(36934) := X"AFC200BC";
        ram_buffer(36935) := X"8FC200BC";
        ram_buffer(36936) := X"00000000";
        ram_buffer(36937) := X"28420008";
        ram_buffer(36938) := X"144000F6";
        ram_buffer(36939) := X"00000000";
        ram_buffer(36940) := X"27C200B8";
        ram_buffer(36941) := X"00403021";
        ram_buffer(36942) := X"8FC501EC";
        ram_buffer(36943) := X"8FC401E8";
        ram_buffer(36944) := X"0C02DCA6";
        ram_buffer(36945) := X"00000000";
        ram_buffer(36946) := X"144001C4";
        ram_buffer(36947) := X"00000000";
        ram_buffer(36948) := X"27D000C4";
        ram_buffer(36949) := X"100000EB";
        ram_buffer(36950) := X"00000000";
        ram_buffer(36951) := X"8FC200B4";
        ram_buffer(36952) := X"00000000";
        ram_buffer(36953) := X"28420002";
        ram_buffer(36954) := X"10400004";
        ram_buffer(36955) := X"00000000";
        ram_buffer(36956) := X"32420001";
        ram_buffer(36957) := X"104000A9";
        ram_buffer(36958) := X"00000000";
        ram_buffer(36959) := X"AE130000";
        ram_buffer(36960) := X"24020001";
        ram_buffer(36961) := X"AE020004";
        ram_buffer(36962) := X"8FC200C0";
        ram_buffer(36963) := X"00000000";
        ram_buffer(36964) := X"24420001";
        ram_buffer(36965) := X"AFC200C0";
        ram_buffer(36966) := X"26100008";
        ram_buffer(36967) := X"8FC200BC";
        ram_buffer(36968) := X"00000000";
        ram_buffer(36969) := X"24420001";
        ram_buffer(36970) := X"AFC200BC";
        ram_buffer(36971) := X"8FC200BC";
        ram_buffer(36972) := X"00000000";
        ram_buffer(36973) := X"28420008";
        ram_buffer(36974) := X"1440000A";
        ram_buffer(36975) := X"00000000";
        ram_buffer(36976) := X"27C200B8";
        ram_buffer(36977) := X"00403021";
        ram_buffer(36978) := X"8FC501EC";
        ram_buffer(36979) := X"8FC401E8";
        ram_buffer(36980) := X"0C02DCA6";
        ram_buffer(36981) := X"00000000";
        ram_buffer(36982) := X"144001A3";
        ram_buffer(36983) := X"00000000";
        ram_buffer(36984) := X"27D000C4";
        ram_buffer(36985) := X"26730001";
        ram_buffer(36986) := X"8FC20084";
        ram_buffer(36987) := X"00000000";
        ram_buffer(36988) := X"AE020000";
        ram_buffer(36989) := X"8FC20088";
        ram_buffer(36990) := X"00000000";
        ram_buffer(36991) := X"AE020004";
        ram_buffer(36992) := X"8FC300C0";
        ram_buffer(36993) := X"8FC20088";
        ram_buffer(36994) := X"00000000";
        ram_buffer(36995) := X"00621021";
        ram_buffer(36996) := X"AFC200C0";
        ram_buffer(36997) := X"26100008";
        ram_buffer(36998) := X"8FC200BC";
        ram_buffer(36999) := X"00000000";
        ram_buffer(37000) := X"24420001";
        ram_buffer(37001) := X"AFC200BC";
        ram_buffer(37002) := X"8FC200BC";
        ram_buffer(37003) := X"00000000";
        ram_buffer(37004) := X"28420008";
        ram_buffer(37005) := X"1440000A";
        ram_buffer(37006) := X"00000000";
        ram_buffer(37007) := X"27C200B8";
        ram_buffer(37008) := X"00403021";
        ram_buffer(37009) := X"8FC501EC";
        ram_buffer(37010) := X"8FC401E8";
        ram_buffer(37011) := X"0C02DCA6";
        ram_buffer(37012) := X"00000000";
        ram_buffer(37013) := X"14400187";
        ram_buffer(37014) := X"00000000";
        ram_buffer(37015) := X"27D000C4";
        ram_buffer(37016) := X"8FC300A4";
        ram_buffer(37017) := X"8FC200A0";
        ram_buffer(37018) := X"00003821";
        ram_buffer(37019) := X"00003021";
        ram_buffer(37020) := X"00602821";
        ram_buffer(37021) := X"00402021";
        ram_buffer(37022) := X"0C03167F";
        ram_buffer(37023) := X"00000000";
        ram_buffer(37024) := X"10400021";
        ram_buffer(37025) := X"00000000";
        ram_buffer(37026) := X"AE130000";
        ram_buffer(37027) := X"8FC200B4";
        ram_buffer(37028) := X"00000000";
        ram_buffer(37029) := X"2442FFFF";
        ram_buffer(37030) := X"AE020004";
        ram_buffer(37031) := X"8FC300C0";
        ram_buffer(37032) := X"8FC200B4";
        ram_buffer(37033) := X"00000000";
        ram_buffer(37034) := X"00621021";
        ram_buffer(37035) := X"2442FFFF";
        ram_buffer(37036) := X"AFC200C0";
        ram_buffer(37037) := X"26100008";
        ram_buffer(37038) := X"8FC200BC";
        ram_buffer(37039) := X"00000000";
        ram_buffer(37040) := X"24420001";
        ram_buffer(37041) := X"AFC200BC";
        ram_buffer(37042) := X"8FC200BC";
        ram_buffer(37043) := X"00000000";
        ram_buffer(37044) := X"28420008";
        ram_buffer(37045) := X"1440006D";
        ram_buffer(37046) := X"00000000";
        ram_buffer(37047) := X"27C200B8";
        ram_buffer(37048) := X"00403021";
        ram_buffer(37049) := X"8FC501EC";
        ram_buffer(37050) := X"8FC401E8";
        ram_buffer(37051) := X"0C02DCA6";
        ram_buffer(37052) := X"00000000";
        ram_buffer(37053) := X"14400162";
        ram_buffer(37054) := X"00000000";
        ram_buffer(37055) := X"27D000C4";
        ram_buffer(37056) := X"10000062";
        ram_buffer(37057) := X"00000000";
        ram_buffer(37058) := X"8FC200B4";
        ram_buffer(37059) := X"00000000";
        ram_buffer(37060) := X"2451FFFF";
        ram_buffer(37061) := X"1A20005D";
        ram_buffer(37062) := X"00000000";
        ram_buffer(37063) := X"1000001E";
        ram_buffer(37064) := X"00000000";
        ram_buffer(37065) := X"3C02100D";
        ram_buffer(37066) := X"2442A254";
        ram_buffer(37067) := X"AE020000";
        ram_buffer(37068) := X"24020010";
        ram_buffer(37069) := X"AE020004";
        ram_buffer(37070) := X"8FC200C0";
        ram_buffer(37071) := X"00000000";
        ram_buffer(37072) := X"24420010";
        ram_buffer(37073) := X"AFC200C0";
        ram_buffer(37074) := X"26100008";
        ram_buffer(37075) := X"8FC200BC";
        ram_buffer(37076) := X"00000000";
        ram_buffer(37077) := X"24420001";
        ram_buffer(37078) := X"AFC200BC";
        ram_buffer(37079) := X"8FC200BC";
        ram_buffer(37080) := X"00000000";
        ram_buffer(37081) := X"28420008";
        ram_buffer(37082) := X"1440000A";
        ram_buffer(37083) := X"00000000";
        ram_buffer(37084) := X"27C200B8";
        ram_buffer(37085) := X"00403021";
        ram_buffer(37086) := X"8FC501EC";
        ram_buffer(37087) := X"8FC401E8";
        ram_buffer(37088) := X"0C02DCA6";
        ram_buffer(37089) := X"00000000";
        ram_buffer(37090) := X"14400140";
        ram_buffer(37091) := X"00000000";
        ram_buffer(37092) := X"27D000C4";
        ram_buffer(37093) := X"2631FFF0";
        ram_buffer(37094) := X"2A220011";
        ram_buffer(37095) := X"1040FFE1";
        ram_buffer(37096) := X"00000000";
        ram_buffer(37097) := X"3C02100D";
        ram_buffer(37098) := X"2442A254";
        ram_buffer(37099) := X"AE020000";
        ram_buffer(37100) := X"02201021";
        ram_buffer(37101) := X"AE020004";
        ram_buffer(37102) := X"8FC300C0";
        ram_buffer(37103) := X"02201021";
        ram_buffer(37104) := X"00621021";
        ram_buffer(37105) := X"AFC200C0";
        ram_buffer(37106) := X"26100008";
        ram_buffer(37107) := X"8FC200BC";
        ram_buffer(37108) := X"00000000";
        ram_buffer(37109) := X"24420001";
        ram_buffer(37110) := X"AFC200BC";
        ram_buffer(37111) := X"8FC200BC";
        ram_buffer(37112) := X"00000000";
        ram_buffer(37113) := X"28420008";
        ram_buffer(37114) := X"14400028";
        ram_buffer(37115) := X"00000000";
        ram_buffer(37116) := X"27C200B8";
        ram_buffer(37117) := X"00403021";
        ram_buffer(37118) := X"8FC501EC";
        ram_buffer(37119) := X"8FC401E8";
        ram_buffer(37120) := X"0C02DCA6";
        ram_buffer(37121) := X"00000000";
        ram_buffer(37122) := X"14400123";
        ram_buffer(37123) := X"00000000";
        ram_buffer(37124) := X"27D000C4";
        ram_buffer(37125) := X"1000001D";
        ram_buffer(37126) := X"00000000";
        ram_buffer(37127) := X"AE130000";
        ram_buffer(37128) := X"24020001";
        ram_buffer(37129) := X"AE020004";
        ram_buffer(37130) := X"8FC200C0";
        ram_buffer(37131) := X"00000000";
        ram_buffer(37132) := X"24420001";
        ram_buffer(37133) := X"AFC200C0";
        ram_buffer(37134) := X"26100008";
        ram_buffer(37135) := X"8FC200BC";
        ram_buffer(37136) := X"00000000";
        ram_buffer(37137) := X"24420001";
        ram_buffer(37138) := X"AFC200BC";
        ram_buffer(37139) := X"8FC200BC";
        ram_buffer(37140) := X"00000000";
        ram_buffer(37141) := X"28420008";
        ram_buffer(37142) := X"1440000D";
        ram_buffer(37143) := X"00000000";
        ram_buffer(37144) := X"27C200B8";
        ram_buffer(37145) := X"00403021";
        ram_buffer(37146) := X"8FC501EC";
        ram_buffer(37147) := X"8FC401E8";
        ram_buffer(37148) := X"0C02DCA6";
        ram_buffer(37149) := X"00000000";
        ram_buffer(37150) := X"1440010A";
        ram_buffer(37151) := X"00000000";
        ram_buffer(37152) := X"27D000C4";
        ram_buffer(37153) := X"10000002";
        ram_buffer(37154) := X"00000000";
        ram_buffer(37155) := X"00000000";
        ram_buffer(37156) := X"27C200AC";
        ram_buffer(37157) := X"AE020000";
        ram_buffer(37158) := X"8FC20048";
        ram_buffer(37159) := X"00000000";
        ram_buffer(37160) := X"AE020004";
        ram_buffer(37161) := X"8FC300C0";
        ram_buffer(37162) := X"8FC20048";
        ram_buffer(37163) := X"00000000";
        ram_buffer(37164) := X"00621021";
        ram_buffer(37165) := X"AFC200C0";
        ram_buffer(37166) := X"26100008";
        ram_buffer(37167) := X"8FC200BC";
        ram_buffer(37168) := X"00000000";
        ram_buffer(37169) := X"24420001";
        ram_buffer(37170) := X"AFC200BC";
        ram_buffer(37171) := X"8FC200BC";
        ram_buffer(37172) := X"00000000";
        ram_buffer(37173) := X"28420008";
        ram_buffer(37174) := X"1440000A";
        ram_buffer(37175) := X"00000000";
        ram_buffer(37176) := X"27C200B8";
        ram_buffer(37177) := X"00403021";
        ram_buffer(37178) := X"8FC501EC";
        ram_buffer(37179) := X"8FC401E8";
        ram_buffer(37180) := X"0C02DCA6";
        ram_buffer(37181) := X"00000000";
        ram_buffer(37182) := X"144000ED";
        ram_buffer(37183) := X"00000000";
        ram_buffer(37184) := X"27D000C4";
        ram_buffer(37185) := X"32420004";
        ram_buffer(37186) := X"10400045";
        ram_buffer(37187) := X"00000000";
        ram_buffer(37188) := X"8FC30034";
        ram_buffer(37189) := X"8FC20068";
        ram_buffer(37190) := X"00000000";
        ram_buffer(37191) := X"00628823";
        ram_buffer(37192) := X"1A20003F";
        ram_buffer(37193) := X"00000000";
        ram_buffer(37194) := X"1000001E";
        ram_buffer(37195) := X"00000000";
        ram_buffer(37196) := X"3C02100D";
        ram_buffer(37197) := X"2442A244";
        ram_buffer(37198) := X"AE020000";
        ram_buffer(37199) := X"24020010";
        ram_buffer(37200) := X"AE020004";
        ram_buffer(37201) := X"8FC200C0";
        ram_buffer(37202) := X"00000000";
        ram_buffer(37203) := X"24420010";
        ram_buffer(37204) := X"AFC200C0";
        ram_buffer(37205) := X"26100008";
        ram_buffer(37206) := X"8FC200BC";
        ram_buffer(37207) := X"00000000";
        ram_buffer(37208) := X"24420001";
        ram_buffer(37209) := X"AFC200BC";
        ram_buffer(37210) := X"8FC200BC";
        ram_buffer(37211) := X"00000000";
        ram_buffer(37212) := X"28420008";
        ram_buffer(37213) := X"1440000A";
        ram_buffer(37214) := X"00000000";
        ram_buffer(37215) := X"27C200B8";
        ram_buffer(37216) := X"00403021";
        ram_buffer(37217) := X"8FC501EC";
        ram_buffer(37218) := X"8FC401E8";
        ram_buffer(37219) := X"0C02DCA6";
        ram_buffer(37220) := X"00000000";
        ram_buffer(37221) := X"144000C9";
        ram_buffer(37222) := X"00000000";
        ram_buffer(37223) := X"27D000C4";
        ram_buffer(37224) := X"2631FFF0";
        ram_buffer(37225) := X"2A220011";
        ram_buffer(37226) := X"1040FFE1";
        ram_buffer(37227) := X"00000000";
        ram_buffer(37228) := X"3C02100D";
        ram_buffer(37229) := X"2442A244";
        ram_buffer(37230) := X"AE020000";
        ram_buffer(37231) := X"02201021";
        ram_buffer(37232) := X"AE020004";
        ram_buffer(37233) := X"8FC200C0";
        ram_buffer(37234) := X"02201821";
        ram_buffer(37235) := X"00431021";
        ram_buffer(37236) := X"AFC200C0";
        ram_buffer(37237) := X"26100008";
        ram_buffer(37238) := X"8FC200BC";
        ram_buffer(37239) := X"00000000";
        ram_buffer(37240) := X"24420001";
        ram_buffer(37241) := X"AFC200BC";
        ram_buffer(37242) := X"8FC200BC";
        ram_buffer(37243) := X"00000000";
        ram_buffer(37244) := X"28420008";
        ram_buffer(37245) := X"1440000A";
        ram_buffer(37246) := X"00000000";
        ram_buffer(37247) := X"27C200B8";
        ram_buffer(37248) := X"00403021";
        ram_buffer(37249) := X"8FC501EC";
        ram_buffer(37250) := X"8FC401E8";
        ram_buffer(37251) := X"0C02DCA6";
        ram_buffer(37252) := X"00000000";
        ram_buffer(37253) := X"144000AC";
        ram_buffer(37254) := X"00000000";
        ram_buffer(37255) := X"27D000C4";
        ram_buffer(37256) := X"8FC30034";
        ram_buffer(37257) := X"8FC20068";
        ram_buffer(37258) := X"00000000";
        ram_buffer(37259) := X"0043202A";
        ram_buffer(37260) := X"10800002";
        ram_buffer(37261) := X"00000000";
        ram_buffer(37262) := X"00601021";
        ram_buffer(37263) := X"8FC30030";
        ram_buffer(37264) := X"00000000";
        ram_buffer(37265) := X"00621021";
        ram_buffer(37266) := X"AFC20030";
        ram_buffer(37267) := X"8FC200C0";
        ram_buffer(37268) := X"00000000";
        ram_buffer(37269) := X"10400009";
        ram_buffer(37270) := X"00000000";
        ram_buffer(37271) := X"27C200B8";
        ram_buffer(37272) := X"00403021";
        ram_buffer(37273) := X"8FC501EC";
        ram_buffer(37274) := X"8FC401E8";
        ram_buffer(37275) := X"0C02DCA6";
        ram_buffer(37276) := X"00000000";
        ram_buffer(37277) := X"14400097";
        ram_buffer(37278) := X"00000000";
        ram_buffer(37279) := X"AFC000BC";
        ram_buffer(37280) := X"27D000C4";
        ram_buffer(37281) := X"8FC20074";
        ram_buffer(37282) := X"00000000";
        ram_buffer(37283) := X"1040F460";
        ram_buffer(37284) := X"00000000";
        ram_buffer(37285) := X"8FC50074";
        ram_buffer(37286) := X"8FC401E8";
        ram_buffer(37287) := X"0C027301";
        ram_buffer(37288) := X"00000000";
        ram_buffer(37289) := X"AFC00074";
        ram_buffer(37290) := X"1000F459";
        ram_buffer(37291) := X"00000000";
        ram_buffer(37292) := X"00000000";
        ram_buffer(37293) := X"10000002";
        ram_buffer(37294) := X"00000000";
        ram_buffer(37295) := X"00000000";
        ram_buffer(37296) := X"8FC200C0";
        ram_buffer(37297) := X"00000000";
        ram_buffer(37298) := X"10400009";
        ram_buffer(37299) := X"00000000";
        ram_buffer(37300) := X"27C200B8";
        ram_buffer(37301) := X"00403021";
        ram_buffer(37302) := X"8FC501EC";
        ram_buffer(37303) := X"8FC401E8";
        ram_buffer(37304) := X"0C02DCA6";
        ram_buffer(37305) := X"00000000";
        ram_buffer(37306) := X"1440007D";
        ram_buffer(37307) := X"00000000";
        ram_buffer(37308) := X"AFC000BC";
        ram_buffer(37309) := X"27D000C4";
        ram_buffer(37310) := X"1000007A";
        ram_buffer(37311) := X"00000000";
        ram_buffer(37312) := X"00000000";
        ram_buffer(37313) := X"10000077";
        ram_buffer(37314) := X"00000000";
        ram_buffer(37315) := X"00000000";
        ram_buffer(37316) := X"10000074";
        ram_buffer(37317) := X"00000000";
        ram_buffer(37318) := X"00000000";
        ram_buffer(37319) := X"10000071";
        ram_buffer(37320) := X"00000000";
        ram_buffer(37321) := X"00000000";
        ram_buffer(37322) := X"1000006E";
        ram_buffer(37323) := X"00000000";
        ram_buffer(37324) := X"00000000";
        ram_buffer(37325) := X"1000006B";
        ram_buffer(37326) := X"00000000";
        ram_buffer(37327) := X"00000000";
        ram_buffer(37328) := X"10000068";
        ram_buffer(37329) := X"00000000";
        ram_buffer(37330) := X"00000000";
        ram_buffer(37331) := X"10000065";
        ram_buffer(37332) := X"00000000";
        ram_buffer(37333) := X"00000000";
        ram_buffer(37334) := X"10000062";
        ram_buffer(37335) := X"00000000";
        ram_buffer(37336) := X"00000000";
        ram_buffer(37337) := X"1000005F";
        ram_buffer(37338) := X"00000000";
        ram_buffer(37339) := X"00000000";
        ram_buffer(37340) := X"1000005C";
        ram_buffer(37341) := X"00000000";
        ram_buffer(37342) := X"00000000";
        ram_buffer(37343) := X"10000059";
        ram_buffer(37344) := X"00000000";
        ram_buffer(37345) := X"00000000";
        ram_buffer(37346) := X"10000056";
        ram_buffer(37347) := X"00000000";
        ram_buffer(37348) := X"00000000";
        ram_buffer(37349) := X"10000053";
        ram_buffer(37350) := X"00000000";
        ram_buffer(37351) := X"00000000";
        ram_buffer(37352) := X"10000050";
        ram_buffer(37353) := X"00000000";
        ram_buffer(37354) := X"00000000";
        ram_buffer(37355) := X"1000004D";
        ram_buffer(37356) := X"00000000";
        ram_buffer(37357) := X"00000000";
        ram_buffer(37358) := X"1000004A";
        ram_buffer(37359) := X"00000000";
        ram_buffer(37360) := X"00000000";
        ram_buffer(37361) := X"10000047";
        ram_buffer(37362) := X"00000000";
        ram_buffer(37363) := X"00000000";
        ram_buffer(37364) := X"10000044";
        ram_buffer(37365) := X"00000000";
        ram_buffer(37366) := X"00000000";
        ram_buffer(37367) := X"10000041";
        ram_buffer(37368) := X"00000000";
        ram_buffer(37369) := X"00000000";
        ram_buffer(37370) := X"1000003E";
        ram_buffer(37371) := X"00000000";
        ram_buffer(37372) := X"00000000";
        ram_buffer(37373) := X"1000003B";
        ram_buffer(37374) := X"00000000";
        ram_buffer(37375) := X"00000000";
        ram_buffer(37376) := X"10000038";
        ram_buffer(37377) := X"00000000";
        ram_buffer(37378) := X"00000000";
        ram_buffer(37379) := X"10000035";
        ram_buffer(37380) := X"00000000";
        ram_buffer(37381) := X"00000000";
        ram_buffer(37382) := X"10000032";
        ram_buffer(37383) := X"00000000";
        ram_buffer(37384) := X"00000000";
        ram_buffer(37385) := X"1000002F";
        ram_buffer(37386) := X"00000000";
        ram_buffer(37387) := X"00000000";
        ram_buffer(37388) := X"1000002C";
        ram_buffer(37389) := X"00000000";
        ram_buffer(37390) := X"00000000";
        ram_buffer(37391) := X"10000029";
        ram_buffer(37392) := X"00000000";
        ram_buffer(37393) := X"00000000";
        ram_buffer(37394) := X"10000026";
        ram_buffer(37395) := X"00000000";
        ram_buffer(37396) := X"00000000";
        ram_buffer(37397) := X"10000023";
        ram_buffer(37398) := X"00000000";
        ram_buffer(37399) := X"00000000";
        ram_buffer(37400) := X"10000020";
        ram_buffer(37401) := X"00000000";
        ram_buffer(37402) := X"00000000";
        ram_buffer(37403) := X"1000001D";
        ram_buffer(37404) := X"00000000";
        ram_buffer(37405) := X"00000000";
        ram_buffer(37406) := X"1000001A";
        ram_buffer(37407) := X"00000000";
        ram_buffer(37408) := X"00000000";
        ram_buffer(37409) := X"10000017";
        ram_buffer(37410) := X"00000000";
        ram_buffer(37411) := X"00000000";
        ram_buffer(37412) := X"10000014";
        ram_buffer(37413) := X"00000000";
        ram_buffer(37414) := X"00000000";
        ram_buffer(37415) := X"10000011";
        ram_buffer(37416) := X"00000000";
        ram_buffer(37417) := X"00000000";
        ram_buffer(37418) := X"1000000E";
        ram_buffer(37419) := X"00000000";
        ram_buffer(37420) := X"00000000";
        ram_buffer(37421) := X"1000000B";
        ram_buffer(37422) := X"00000000";
        ram_buffer(37423) := X"00000000";
        ram_buffer(37424) := X"10000008";
        ram_buffer(37425) := X"00000000";
        ram_buffer(37426) := X"00000000";
        ram_buffer(37427) := X"10000005";
        ram_buffer(37428) := X"00000000";
        ram_buffer(37429) := X"00000000";
        ram_buffer(37430) := X"10000002";
        ram_buffer(37431) := X"00000000";
        ram_buffer(37432) := X"00000000";
        ram_buffer(37433) := X"8FC20074";
        ram_buffer(37434) := X"00000000";
        ram_buffer(37435) := X"10400005";
        ram_buffer(37436) := X"00000000";
        ram_buffer(37437) := X"8FC50074";
        ram_buffer(37438) := X"8FC401E8";
        ram_buffer(37439) := X"0C027301";
        ram_buffer(37440) := X"00000000";
        ram_buffer(37441) := X"8FC201EC";
        ram_buffer(37442) := X"00000000";
        ram_buffer(37443) := X"8442000C";
        ram_buffer(37444) := X"00000000";
        ram_buffer(37445) := X"3042FFFF";
        ram_buffer(37446) := X"30420040";
        ram_buffer(37447) := X"14400004";
        ram_buffer(37448) := X"00000000";
        ram_buffer(37449) := X"8FC20030";
        ram_buffer(37450) := X"10000003";
        ram_buffer(37451) := X"00000000";
        ram_buffer(37452) := X"2402FFFF";
        ram_buffer(37453) := X"00000000";
        ram_buffer(37454) := X"03C0E821";
        ram_buffer(37455) := X"8FBF01E4";
        ram_buffer(37456) := X"8FBE01E0";
        ram_buffer(37457) := X"8FB701DC";
        ram_buffer(37458) := X"8FB601D8";
        ram_buffer(37459) := X"8FB501D4";
        ram_buffer(37460) := X"8FB401D0";
        ram_buffer(37461) := X"8FB301CC";
        ram_buffer(37462) := X"8FB201C8";
        ram_buffer(37463) := X"8FB101C4";
        ram_buffer(37464) := X"8FB001C0";
        ram_buffer(37465) := X"27BD01E8";
        ram_buffer(37466) := X"03E00008";
        ram_buffer(37467) := X"00000000";
        ram_buffer(37468) := X"27BDFFB0";
        ram_buffer(37469) := X"AFBF004C";
        ram_buffer(37470) := X"AFBE0048";
        ram_buffer(37471) := X"03A0F021";
        ram_buffer(37472) := X"AFC40050";
        ram_buffer(37473) := X"AFC7005C";
        ram_buffer(37474) := X"AFC60058";
        ram_buffer(37475) := X"8FC3005C";
        ram_buffer(37476) := X"8FC20058";
        ram_buffer(37477) := X"AFC30044";
        ram_buffer(37478) := X"AFC20040";
        ram_buffer(37479) := X"8FC20040";
        ram_buffer(37480) := X"00000000";
        ram_buffer(37481) := X"0441000D";
        ram_buffer(37482) := X"00000000";
        ram_buffer(37483) := X"8FC30058";
        ram_buffer(37484) := X"3C028000";
        ram_buffer(37485) := X"00621026";
        ram_buffer(37486) := X"AFC20058";
        ram_buffer(37487) := X"8FC2005C";
        ram_buffer(37488) := X"00000000";
        ram_buffer(37489) := X"AFC2005C";
        ram_buffer(37490) := X"8FC20068";
        ram_buffer(37491) := X"2403002D";
        ram_buffer(37492) := X"A0430000";
        ram_buffer(37493) := X"10000004";
        ram_buffer(37494) := X"00000000";
        ram_buffer(37495) := X"8FC20068";
        ram_buffer(37496) := X"00000000";
        ram_buffer(37497) := X"A0400000";
        ram_buffer(37498) := X"8FC30070";
        ram_buffer(37499) := X"24020061";
        ram_buffer(37500) := X"10620005";
        ram_buffer(37501) := X"00000000";
        ram_buffer(37502) := X"8FC30070";
        ram_buffer(37503) := X"24020041";
        ram_buffer(37504) := X"146200B3";
        ram_buffer(37505) := X"00000000";
        ram_buffer(37506) := X"8FC6006C";
        ram_buffer(37507) := X"8FC5005C";
        ram_buffer(37508) := X"8FC40058";
        ram_buffer(37509) := X"0C02CB50";
        ram_buffer(37510) := X"00000000";
        ram_buffer(37511) := X"8F8780AC";
        ram_buffer(37512) := X"8F8680A8";
        ram_buffer(37513) := X"00602821";
        ram_buffer(37514) := X"00402021";
        ram_buffer(37515) := X"0C03144F";
        ram_buffer(37516) := X"00000000";
        ram_buffer(37517) := X"AFC3005C";
        ram_buffer(37518) := X"AFC20058";
        ram_buffer(37519) := X"00003821";
        ram_buffer(37520) := X"00003021";
        ram_buffer(37521) := X"8FC5005C";
        ram_buffer(37522) := X"8FC40058";
        ram_buffer(37523) := X"0C03167F";
        ram_buffer(37524) := X"00000000";
        ram_buffer(37525) := X"14400004";
        ram_buffer(37526) := X"00000000";
        ram_buffer(37527) := X"8FC2006C";
        ram_buffer(37528) := X"24030001";
        ram_buffer(37529) := X"AC430000";
        ram_buffer(37530) := X"8FC30070";
        ram_buffer(37531) := X"24020061";
        ram_buffer(37532) := X"14620005";
        ram_buffer(37533) := X"00000000";
        ram_buffer(37534) := X"3C02100D";
        ram_buffer(37535) := X"2442A088";
        ram_buffer(37536) := X"10000003";
        ram_buffer(37537) := X"00000000";
        ram_buffer(37538) := X"3C02100D";
        ram_buffer(37539) := X"2442A0A4";
        ram_buffer(37540) := X"AFC20030";
        ram_buffer(37541) := X"8FC20078";
        ram_buffer(37542) := X"00000000";
        ram_buffer(37543) := X"AFC2002C";
        ram_buffer(37544) := X"8F8780B4";
        ram_buffer(37545) := X"8F8680B0";
        ram_buffer(37546) := X"8FC5005C";
        ram_buffer(37547) := X"8FC40058";
        ram_buffer(37548) := X"0C03174A";
        ram_buffer(37549) := X"00000000";
        ram_buffer(37550) := X"AFC3005C";
        ram_buffer(37551) := X"AFC20058";
        ram_buffer(37552) := X"8FC5005C";
        ram_buffer(37553) := X"8FC40058";
        ram_buffer(37554) := X"0C031B37";
        ram_buffer(37555) := X"00000000";
        ram_buffer(37556) := X"AFC20028";
        ram_buffer(37557) := X"8FC40028";
        ram_buffer(37558) := X"0C031B7C";
        ram_buffer(37559) := X"00000000";
        ram_buffer(37560) := X"00603821";
        ram_buffer(37561) := X"00403021";
        ram_buffer(37562) := X"8FC5005C";
        ram_buffer(37563) := X"8FC40058";
        ram_buffer(37564) := X"0C0318D3";
        ram_buffer(37565) := X"00000000";
        ram_buffer(37566) := X"AFC3005C";
        ram_buffer(37567) := X"AFC20058";
        ram_buffer(37568) := X"8FC2002C";
        ram_buffer(37569) := X"00000000";
        ram_buffer(37570) := X"24430001";
        ram_buffer(37571) := X"AFC3002C";
        ram_buffer(37572) := X"8FC30028";
        ram_buffer(37573) := X"8FC40030";
        ram_buffer(37574) := X"00000000";
        ram_buffer(37575) := X"00831821";
        ram_buffer(37576) := X"80630000";
        ram_buffer(37577) := X"00000000";
        ram_buffer(37578) := X"A0430000";
        ram_buffer(37579) := X"8FC20060";
        ram_buffer(37580) := X"00000000";
        ram_buffer(37581) := X"2443FFFF";
        ram_buffer(37582) := X"AFC30060";
        ram_buffer(37583) := X"10400009";
        ram_buffer(37584) := X"00000000";
        ram_buffer(37585) := X"00003821";
        ram_buffer(37586) := X"00003021";
        ram_buffer(37587) := X"8FC5005C";
        ram_buffer(37588) := X"8FC40058";
        ram_buffer(37589) := X"0C03167F";
        ram_buffer(37590) := X"00000000";
        ram_buffer(37591) := X"1440FFD0";
        ram_buffer(37592) := X"00000000";
        ram_buffer(37593) := X"8F8780BC";
        ram_buffer(37594) := X"8F8680B8";
        ram_buffer(37595) := X"8FC5005C";
        ram_buffer(37596) := X"8FC40058";
        ram_buffer(37597) := X"0C0316AB";
        ram_buffer(37598) := X"00000000";
        ram_buffer(37599) := X"1C40000E";
        ram_buffer(37600) := X"00000000";
        ram_buffer(37601) := X"8F8780BC";
        ram_buffer(37602) := X"8F8680B8";
        ram_buffer(37603) := X"8FC5005C";
        ram_buffer(37604) := X"8FC40058";
        ram_buffer(37605) := X"0C03167F";
        ram_buffer(37606) := X"00000000";
        ram_buffer(37607) := X"14400034";
        ram_buffer(37608) := X"00000000";
        ram_buffer(37609) := X"8FC20028";
        ram_buffer(37610) := X"00000000";
        ram_buffer(37611) := X"30420001";
        ram_buffer(37612) := X"10400037";
        ram_buffer(37613) := X"00000000";
        ram_buffer(37614) := X"8FC2002C";
        ram_buffer(37615) := X"00000000";
        ram_buffer(37616) := X"AFC20038";
        ram_buffer(37617) := X"10000004";
        ram_buffer(37618) := X"00000000";
        ram_buffer(37619) := X"8FC20038";
        ram_buffer(37620) := X"24030030";
        ram_buffer(37621) := X"A0430000";
        ram_buffer(37622) := X"8FC20038";
        ram_buffer(37623) := X"00000000";
        ram_buffer(37624) := X"2442FFFF";
        ram_buffer(37625) := X"AFC20038";
        ram_buffer(37626) := X"8FC20038";
        ram_buffer(37627) := X"00000000";
        ram_buffer(37628) := X"80430000";
        ram_buffer(37629) := X"8FC20030";
        ram_buffer(37630) := X"00000000";
        ram_buffer(37631) := X"2442000F";
        ram_buffer(37632) := X"80420000";
        ram_buffer(37633) := X"00000000";
        ram_buffer(37634) := X"1062FFF0";
        ram_buffer(37635) := X"00000000";
        ram_buffer(37636) := X"8FC30038";
        ram_buffer(37637) := X"8FC20038";
        ram_buffer(37638) := X"00000000";
        ram_buffer(37639) := X"80440000";
        ram_buffer(37640) := X"24020039";
        ram_buffer(37641) := X"14820006";
        ram_buffer(37642) := X"00000000";
        ram_buffer(37643) := X"8FC20030";
        ram_buffer(37644) := X"00000000";
        ram_buffer(37645) := X"8042000A";
        ram_buffer(37646) := X"1000000A";
        ram_buffer(37647) := X"00000000";
        ram_buffer(37648) := X"8FC20038";
        ram_buffer(37649) := X"00000000";
        ram_buffer(37650) := X"80420000";
        ram_buffer(37651) := X"00000000";
        ram_buffer(37652) := X"304200FF";
        ram_buffer(37653) := X"24420001";
        ram_buffer(37654) := X"304200FF";
        ram_buffer(37655) := X"00021600";
        ram_buffer(37656) := X"00021603";
        ram_buffer(37657) := X"A0620000";
        ram_buffer(37658) := X"1000000F";
        ram_buffer(37659) := X"00000000";
        ram_buffer(37660) := X"10000007";
        ram_buffer(37661) := X"00000000";
        ram_buffer(37662) := X"8FC2002C";
        ram_buffer(37663) := X"00000000";
        ram_buffer(37664) := X"24430001";
        ram_buffer(37665) := X"AFC3002C";
        ram_buffer(37666) := X"24030030";
        ram_buffer(37667) := X"A0430000";
        ram_buffer(37668) := X"8FC20060";
        ram_buffer(37669) := X"00000000";
        ram_buffer(37670) := X"2443FFFF";
        ram_buffer(37671) := X"AFC30060";
        ram_buffer(37672) := X"0441FFF5";
        ram_buffer(37673) := X"00000000";
        ram_buffer(37674) := X"8FC3002C";
        ram_buffer(37675) := X"8FC20078";
        ram_buffer(37676) := X"00000000";
        ram_buffer(37677) := X"00621823";
        ram_buffer(37678) := X"8FC20074";
        ram_buffer(37679) := X"00000000";
        ram_buffer(37680) := X"AC430000";
        ram_buffer(37681) := X"8FC20078";
        ram_buffer(37682) := X"10000089";
        ram_buffer(37683) := X"00000000";
        ram_buffer(37684) := X"8FC30070";
        ram_buffer(37685) := X"24020066";
        ram_buffer(37686) := X"10620005";
        ram_buffer(37687) := X"00000000";
        ram_buffer(37688) := X"8FC30070";
        ram_buffer(37689) := X"24020046";
        ram_buffer(37690) := X"14620005";
        ram_buffer(37691) := X"00000000";
        ram_buffer(37692) := X"24020003";
        ram_buffer(37693) := X"AFC20028";
        ram_buffer(37694) := X"1000000F";
        ram_buffer(37695) := X"00000000";
        ram_buffer(37696) := X"8FC30070";
        ram_buffer(37697) := X"24020065";
        ram_buffer(37698) := X"10620005";
        ram_buffer(37699) := X"00000000";
        ram_buffer(37700) := X"8FC30070";
        ram_buffer(37701) := X"24020045";
        ram_buffer(37702) := X"14620005";
        ram_buffer(37703) := X"00000000";
        ram_buffer(37704) := X"8FC20060";
        ram_buffer(37705) := X"00000000";
        ram_buffer(37706) := X"24420001";
        ram_buffer(37707) := X"AFC20060";
        ram_buffer(37708) := X"24020002";
        ram_buffer(37709) := X"AFC20028";
        ram_buffer(37710) := X"27C20038";
        ram_buffer(37711) := X"AFA20020";
        ram_buffer(37712) := X"27C20034";
        ram_buffer(37713) := X"AFA2001C";
        ram_buffer(37714) := X"8FC2006C";
        ram_buffer(37715) := X"00000000";
        ram_buffer(37716) := X"AFA20018";
        ram_buffer(37717) := X"8FC20060";
        ram_buffer(37718) := X"00000000";
        ram_buffer(37719) := X"AFA20014";
        ram_buffer(37720) := X"8FC20028";
        ram_buffer(37721) := X"00000000";
        ram_buffer(37722) := X"AFA20010";
        ram_buffer(37723) := X"8FC7005C";
        ram_buffer(37724) := X"8FC60058";
        ram_buffer(37725) := X"8FC40050";
        ram_buffer(37726) := X"0C02AFA3";
        ram_buffer(37727) := X"00000000";
        ram_buffer(37728) := X"AFC20030";
        ram_buffer(37729) := X"8FC30070";
        ram_buffer(37730) := X"24020067";
        ram_buffer(37731) := X"10620005";
        ram_buffer(37732) := X"00000000";
        ram_buffer(37733) := X"8FC30070";
        ram_buffer(37734) := X"24020047";
        ram_buffer(37735) := X"14620006";
        ram_buffer(37736) := X"00000000";
        ram_buffer(37737) := X"8FC20064";
        ram_buffer(37738) := X"00000000";
        ram_buffer(37739) := X"30420001";
        ram_buffer(37740) := X"10400045";
        ram_buffer(37741) := X"00000000";
        ram_buffer(37742) := X"8FC20060";
        ram_buffer(37743) := X"8FC30030";
        ram_buffer(37744) := X"00000000";
        ram_buffer(37745) := X"00621021";
        ram_buffer(37746) := X"AFC2002C";
        ram_buffer(37747) := X"8FC30070";
        ram_buffer(37748) := X"24020066";
        ram_buffer(37749) := X"10620005";
        ram_buffer(37750) := X"00000000";
        ram_buffer(37751) := X"8FC30070";
        ram_buffer(37752) := X"24020046";
        ram_buffer(37753) := X"1462001F";
        ram_buffer(37754) := X"00000000";
        ram_buffer(37755) := X"8FC20030";
        ram_buffer(37756) := X"00000000";
        ram_buffer(37757) := X"80430000";
        ram_buffer(37758) := X"24020030";
        ram_buffer(37759) := X"14620010";
        ram_buffer(37760) := X"00000000";
        ram_buffer(37761) := X"00003821";
        ram_buffer(37762) := X"00003021";
        ram_buffer(37763) := X"8FC5005C";
        ram_buffer(37764) := X"8FC40058";
        ram_buffer(37765) := X"0C03167F";
        ram_buffer(37766) := X"00000000";
        ram_buffer(37767) := X"10400008";
        ram_buffer(37768) := X"00000000";
        ram_buffer(37769) := X"24030001";
        ram_buffer(37770) := X"8FC20060";
        ram_buffer(37771) := X"00000000";
        ram_buffer(37772) := X"00621823";
        ram_buffer(37773) := X"8FC2006C";
        ram_buffer(37774) := X"00000000";
        ram_buffer(37775) := X"AC430000";
        ram_buffer(37776) := X"8FC2006C";
        ram_buffer(37777) := X"00000000";
        ram_buffer(37778) := X"8C420000";
        ram_buffer(37779) := X"00000000";
        ram_buffer(37780) := X"00401821";
        ram_buffer(37781) := X"8FC2002C";
        ram_buffer(37782) := X"00000000";
        ram_buffer(37783) := X"00431021";
        ram_buffer(37784) := X"AFC2002C";
        ram_buffer(37785) := X"00003821";
        ram_buffer(37786) := X"00003021";
        ram_buffer(37787) := X"8FC5005C";
        ram_buffer(37788) := X"8FC40058";
        ram_buffer(37789) := X"0C03167F";
        ram_buffer(37790) := X"00000000";
        ram_buffer(37791) := X"14400004";
        ram_buffer(37792) := X"00000000";
        ram_buffer(37793) := X"8FC2002C";
        ram_buffer(37794) := X"00000000";
        ram_buffer(37795) := X"AFC20038";
        ram_buffer(37796) := X"10000007";
        ram_buffer(37797) := X"00000000";
        ram_buffer(37798) := X"8FC20038";
        ram_buffer(37799) := X"00000000";
        ram_buffer(37800) := X"24430001";
        ram_buffer(37801) := X"AFC30038";
        ram_buffer(37802) := X"24030030";
        ram_buffer(37803) := X"A0430000";
        ram_buffer(37804) := X"8FC30038";
        ram_buffer(37805) := X"8FC2002C";
        ram_buffer(37806) := X"00000000";
        ram_buffer(37807) := X"0062102B";
        ram_buffer(37808) := X"1440FFF5";
        ram_buffer(37809) := X"00000000";
        ram_buffer(37810) := X"8FC20038";
        ram_buffer(37811) := X"00000000";
        ram_buffer(37812) := X"00401821";
        ram_buffer(37813) := X"8FC20030";
        ram_buffer(37814) := X"00000000";
        ram_buffer(37815) := X"00621823";
        ram_buffer(37816) := X"8FC20074";
        ram_buffer(37817) := X"00000000";
        ram_buffer(37818) := X"AC430000";
        ram_buffer(37819) := X"8FC20030";
        ram_buffer(37820) := X"03C0E821";
        ram_buffer(37821) := X"8FBF004C";
        ram_buffer(37822) := X"8FBE0048";
        ram_buffer(37823) := X"27BD0050";
        ram_buffer(37824) := X"03E00008";
        ram_buffer(37825) := X"00000000";
        ram_buffer(37826) := X"27BDFFE0";
        ram_buffer(37827) := X"AFBE001C";
        ram_buffer(37828) := X"AFB10018";
        ram_buffer(37829) := X"AFB00014";
        ram_buffer(37830) := X"03A0F021";
        ram_buffer(37831) := X"AFC40020";
        ram_buffer(37832) := X"AFC50024";
        ram_buffer(37833) := X"AFC60028";
        ram_buffer(37834) := X"8FC30028";
        ram_buffer(37835) := X"24020061";
        ram_buffer(37836) := X"10620005";
        ram_buffer(37837) := X"00000000";
        ram_buffer(37838) := X"8FC30028";
        ram_buffer(37839) := X"24020041";
        ram_buffer(37840) := X"14620004";
        ram_buffer(37841) := X"00000000";
        ram_buffer(37842) := X"24020001";
        ram_buffer(37843) := X"10000002";
        ram_buffer(37844) := X"00000000";
        ram_buffer(37845) := X"00001021";
        ram_buffer(37846) := X"AFC20000";
        ram_buffer(37847) := X"8FD10020";
        ram_buffer(37848) := X"00000000";
        ram_buffer(37849) := X"02201821";
        ram_buffer(37850) := X"24710001";
        ram_buffer(37851) := X"8FC20000";
        ram_buffer(37852) := X"00000000";
        ram_buffer(37853) := X"1040000A";
        ram_buffer(37854) := X"00000000";
        ram_buffer(37855) := X"8FC20028";
        ram_buffer(37856) := X"00000000";
        ram_buffer(37857) := X"304200FF";
        ram_buffer(37858) := X"2442000F";
        ram_buffer(37859) := X"304200FF";
        ram_buffer(37860) := X"00021600";
        ram_buffer(37861) := X"00021603";
        ram_buffer(37862) := X"10000005";
        ram_buffer(37863) := X"00000000";
        ram_buffer(37864) := X"8FC20028";
        ram_buffer(37865) := X"00000000";
        ram_buffer(37866) := X"00021600";
        ram_buffer(37867) := X"00021603";
        ram_buffer(37868) := X"A0620000";
        ram_buffer(37869) := X"8FC20024";
        ram_buffer(37870) := X"00000000";
        ram_buffer(37871) := X"0441000B";
        ram_buffer(37872) := X"00000000";
        ram_buffer(37873) := X"8FC20024";
        ram_buffer(37874) := X"00000000";
        ram_buffer(37875) := X"00021023";
        ram_buffer(37876) := X"AFC20024";
        ram_buffer(37877) := X"02201021";
        ram_buffer(37878) := X"24510001";
        ram_buffer(37879) := X"2403002D";
        ram_buffer(37880) := X"A0430000";
        ram_buffer(37881) := X"10000005";
        ram_buffer(37882) := X"00000000";
        ram_buffer(37883) := X"02201021";
        ram_buffer(37884) := X"24510001";
        ram_buffer(37885) := X"2403002B";
        ram_buffer(37886) := X"A0430000";
        ram_buffer(37887) := X"27D00004";
        ram_buffer(37888) := X"26100007";
        ram_buffer(37889) := X"8FC20024";
        ram_buffer(37890) := X"00000000";
        ram_buffer(37891) := X"2842000A";
        ram_buffer(37892) := X"14400034";
        ram_buffer(37893) := X"00000000";
        ram_buffer(37894) := X"2610FFFF";
        ram_buffer(37895) := X"8FC30024";
        ram_buffer(37896) := X"2402000A";
        ram_buffer(37897) := X"14400002";
        ram_buffer(37898) := X"0062001A";
        ram_buffer(37899) := X"0007000D";
        ram_buffer(37900) := X"00001010";
        ram_buffer(37901) := X"304200FF";
        ram_buffer(37902) := X"24420030";
        ram_buffer(37903) := X"304200FF";
        ram_buffer(37904) := X"00021600";
        ram_buffer(37905) := X"00021603";
        ram_buffer(37906) := X"A2020000";
        ram_buffer(37907) := X"8FC30024";
        ram_buffer(37908) := X"2402000A";
        ram_buffer(37909) := X"14400002";
        ram_buffer(37910) := X"0062001A";
        ram_buffer(37911) := X"0007000D";
        ram_buffer(37912) := X"00001010";
        ram_buffer(37913) := X"00001012";
        ram_buffer(37914) := X"AFC20024";
        ram_buffer(37915) := X"8FC20024";
        ram_buffer(37916) := X"00000000";
        ram_buffer(37917) := X"2842000A";
        ram_buffer(37918) := X"1040FFE7";
        ram_buffer(37919) := X"00000000";
        ram_buffer(37920) := X"2610FFFF";
        ram_buffer(37921) := X"8FC20024";
        ram_buffer(37922) := X"00000000";
        ram_buffer(37923) := X"304200FF";
        ram_buffer(37924) := X"24420030";
        ram_buffer(37925) := X"304200FF";
        ram_buffer(37926) := X"00021600";
        ram_buffer(37927) := X"00021603";
        ram_buffer(37928) := X"A2020000";
        ram_buffer(37929) := X"10000008";
        ram_buffer(37930) := X"00000000";
        ram_buffer(37931) := X"02201021";
        ram_buffer(37932) := X"24510001";
        ram_buffer(37933) := X"02001821";
        ram_buffer(37934) := X"24700001";
        ram_buffer(37935) := X"80630000";
        ram_buffer(37936) := X"00000000";
        ram_buffer(37937) := X"A0430000";
        ram_buffer(37938) := X"27C20004";
        ram_buffer(37939) := X"24420007";
        ram_buffer(37940) := X"0202102B";
        ram_buffer(37941) := X"1440FFF5";
        ram_buffer(37942) := X"00000000";
        ram_buffer(37943) := X"10000013";
        ram_buffer(37944) := X"00000000";
        ram_buffer(37945) := X"8FC20000";
        ram_buffer(37946) := X"00000000";
        ram_buffer(37947) := X"14400005";
        ram_buffer(37948) := X"00000000";
        ram_buffer(37949) := X"02201021";
        ram_buffer(37950) := X"24510001";
        ram_buffer(37951) := X"24030030";
        ram_buffer(37952) := X"A0430000";
        ram_buffer(37953) := X"02201021";
        ram_buffer(37954) := X"24510001";
        ram_buffer(37955) := X"8FC30024";
        ram_buffer(37956) := X"00000000";
        ram_buffer(37957) := X"306300FF";
        ram_buffer(37958) := X"24630030";
        ram_buffer(37959) := X"306300FF";
        ram_buffer(37960) := X"00031E00";
        ram_buffer(37961) := X"00031E03";
        ram_buffer(37962) := X"A0430000";
        ram_buffer(37963) := X"02201821";
        ram_buffer(37964) := X"8FC20020";
        ram_buffer(37965) := X"00000000";
        ram_buffer(37966) := X"00621023";
        ram_buffer(37967) := X"03C0E821";
        ram_buffer(37968) := X"8FBE001C";
        ram_buffer(37969) := X"8FB10018";
        ram_buffer(37970) := X"8FB00014";
        ram_buffer(37971) := X"27BD0020";
        ram_buffer(37972) := X"03E00008";
        ram_buffer(37973) := X"00000000";
        ram_buffer(37974) := X"27BDFCC0";
        ram_buffer(37975) := X"AFBF033C";
        ram_buffer(37976) := X"AFBE0338";
        ram_buffer(37977) := X"AFB70334";
        ram_buffer(37978) := X"AFB60330";
        ram_buffer(37979) := X"AFB5032C";
        ram_buffer(37980) := X"AFB40328";
        ram_buffer(37981) := X"AFB30324";
        ram_buffer(37982) := X"AFB20320";
        ram_buffer(37983) := X"AFB1031C";
        ram_buffer(37984) := X"AFB00318";
        ram_buffer(37985) := X"03A0F021";
        ram_buffer(37986) := X"AFC40340";
        ram_buffer(37987) := X"00A08821";
        ram_buffer(37988) := X"AFC60348";
        ram_buffer(37989) := X"AFC7034C";
        ram_buffer(37990) := X"8FD50348";
        ram_buffer(37991) := X"AFC00020";
        ram_buffer(37992) := X"24020001";
        ram_buffer(37993) := X"AFC20064";
        ram_buffer(37994) := X"AFC00028";
        ram_buffer(37995) := X"8622000C";
        ram_buffer(37996) := X"00000000";
        ram_buffer(37997) := X"3042FFFF";
        ram_buffer(37998) := X"30422000";
        ram_buffer(37999) := X"1440000B";
        ram_buffer(38000) := X"00000000";
        ram_buffer(38001) := X"8622000C";
        ram_buffer(38002) := X"00000000";
        ram_buffer(38003) := X"34422000";
        ram_buffer(38004) := X"00021400";
        ram_buffer(38005) := X"00021403";
        ram_buffer(38006) := X"A622000C";
        ram_buffer(38007) := X"8E230064";
        ram_buffer(38008) := X"2402DFFF";
        ram_buffer(38009) := X"00621024";
        ram_buffer(38010) := X"AE220064";
        ram_buffer(38011) := X"AFC00018";
        ram_buffer(38012) := X"AFC0001C";
        ram_buffer(38013) := X"92A20000";
        ram_buffer(38014) := X"00000000";
        ram_buffer(38015) := X"AFC200A4";
        ram_buffer(38016) := X"8FC20064";
        ram_buffer(38017) := X"00000000";
        ram_buffer(38018) := X"02A2A821";
        ram_buffer(38019) := X"8FC200A4";
        ram_buffer(38020) := X"00000000";
        ram_buffer(38021) := X"104007D2";
        ram_buffer(38022) := X"00000000";
        ram_buffer(38023) := X"8FC30064";
        ram_buffer(38024) := X"24020001";
        ram_buffer(38025) := X"14620031";
        ram_buffer(38026) := X"00000000";
        ram_buffer(38027) := X"8F838090";
        ram_buffer(38028) := X"8FC200A4";
        ram_buffer(38029) := X"00000000";
        ram_buffer(38030) := X"24420001";
        ram_buffer(38031) := X"00621021";
        ram_buffer(38032) := X"80420000";
        ram_buffer(38033) := X"00000000";
        ram_buffer(38034) := X"304200FF";
        ram_buffer(38035) := X"30420008";
        ram_buffer(38036) := X"10400026";
        ram_buffer(38037) := X"00000000";
        ram_buffer(38038) := X"8E220004";
        ram_buffer(38039) := X"00000000";
        ram_buffer(38040) := X"1C400007";
        ram_buffer(38041) := X"00000000";
        ram_buffer(38042) := X"02202821";
        ram_buffer(38043) := X"8FC40340";
        ram_buffer(38044) := X"0C02E477";
        ram_buffer(38045) := X"00000000";
        ram_buffer(38046) := X"14400784";
        ram_buffer(38047) := X"00000000";
        ram_buffer(38048) := X"8F838090";
        ram_buffer(38049) := X"8E220000";
        ram_buffer(38050) := X"00000000";
        ram_buffer(38051) := X"90420000";
        ram_buffer(38052) := X"00000000";
        ram_buffer(38053) := X"24420001";
        ram_buffer(38054) := X"00621021";
        ram_buffer(38055) := X"80420000";
        ram_buffer(38056) := X"00000000";
        ram_buffer(38057) := X"304200FF";
        ram_buffer(38058) := X"30420008";
        ram_buffer(38059) := X"10400777";
        ram_buffer(38060) := X"00000000";
        ram_buffer(38061) := X"8FC2001C";
        ram_buffer(38062) := X"00000000";
        ram_buffer(38063) := X"24420001";
        ram_buffer(38064) := X"AFC2001C";
        ram_buffer(38065) := X"8E220004";
        ram_buffer(38066) := X"00000000";
        ram_buffer(38067) := X"2442FFFF";
        ram_buffer(38068) := X"AE220004";
        ram_buffer(38069) := X"8E220000";
        ram_buffer(38070) := X"00000000";
        ram_buffer(38071) := X"24420001";
        ram_buffer(38072) := X"AE220000";
        ram_buffer(38073) := X"1000FFDC";
        ram_buffer(38074) := X"00000000";
        ram_buffer(38075) := X"8FC300A4";
        ram_buffer(38076) := X"24020025";
        ram_buffer(38077) := X"14620013";
        ram_buffer(38078) := X"00000000";
        ram_buffer(38079) := X"00009021";
        ram_buffer(38080) := X"00008021";
        ram_buffer(38081) := X"02A01021";
        ram_buffer(38082) := X"24550001";
        ram_buffer(38083) := X"90420000";
        ram_buffer(38084) := X"00000000";
        ram_buffer(38085) := X"0040A021";
        ram_buffer(38086) := X"2E82007B";
        ram_buffer(38087) := X"1040010C";
        ram_buffer(38088) := X"00000000";
        ram_buffer(38089) := X"00141880";
        ram_buffer(38090) := X"3C02100D";
        ram_buffer(38091) := X"2442A26C";
        ram_buffer(38092) := X"00621021";
        ram_buffer(38093) := X"8C420000";
        ram_buffer(38094) := X"00000000";
        ram_buffer(38095) := X"00400008";
        ram_buffer(38096) := X"00000000";
        ram_buffer(38097) := X"00000000";
        ram_buffer(38098) := X"8FC20064";
        ram_buffer(38099) := X"00000000";
        ram_buffer(38100) := X"00021023";
        ram_buffer(38101) := X"02A21021";
        ram_buffer(38102) := X"AFC2002C";
        ram_buffer(38103) := X"0000A021";
        ram_buffer(38104) := X"10000025";
        ram_buffer(38105) := X"00000000";
        ram_buffer(38106) := X"8E220004";
        ram_buffer(38107) := X"00000000";
        ram_buffer(38108) := X"1C400007";
        ram_buffer(38109) := X"00000000";
        ram_buffer(38110) := X"02202821";
        ram_buffer(38111) := X"8FC40340";
        ram_buffer(38112) := X"0C02E477";
        ram_buffer(38113) := X"00000000";
        ram_buffer(38114) := X"1440074F";
        ram_buffer(38115) := X"00000000";
        ram_buffer(38116) := X"8E220000";
        ram_buffer(38117) := X"00000000";
        ram_buffer(38118) := X"90430000";
        ram_buffer(38119) := X"8FC2002C";
        ram_buffer(38120) := X"00000000";
        ram_buffer(38121) := X"90420000";
        ram_buffer(38122) := X"00000000";
        ram_buffer(38123) := X"1462076F";
        ram_buffer(38124) := X"00000000";
        ram_buffer(38125) := X"8E220004";
        ram_buffer(38126) := X"00000000";
        ram_buffer(38127) := X"2442FFFF";
        ram_buffer(38128) := X"AE220004";
        ram_buffer(38129) := X"8E220000";
        ram_buffer(38130) := X"00000000";
        ram_buffer(38131) := X"24420001";
        ram_buffer(38132) := X"AE220000";
        ram_buffer(38133) := X"8FC2001C";
        ram_buffer(38134) := X"00000000";
        ram_buffer(38135) := X"24420001";
        ram_buffer(38136) := X"AFC2001C";
        ram_buffer(38137) := X"8FC2002C";
        ram_buffer(38138) := X"00000000";
        ram_buffer(38139) := X"24420001";
        ram_buffer(38140) := X"AFC2002C";
        ram_buffer(38141) := X"26940001";
        ram_buffer(38142) := X"8FC20064";
        ram_buffer(38143) := X"00000000";
        ram_buffer(38144) := X"0282102A";
        ram_buffer(38145) := X"1440FFD8";
        ram_buffer(38146) := X"00000000";
        ram_buffer(38147) := X"1000072C";
        ram_buffer(38148) := X"00000000";
        ram_buffer(38149) := X"36100010";
        ram_buffer(38150) := X"1000FFBA";
        ram_buffer(38151) := X"00000000";
        ram_buffer(38152) := X"92A30000";
        ram_buffer(38153) := X"2402006C";
        ram_buffer(38154) := X"14620005";
        ram_buffer(38155) := X"00000000";
        ram_buffer(38156) := X"26B50001";
        ram_buffer(38157) := X"36100002";
        ram_buffer(38158) := X"1000FFB2";
        ram_buffer(38159) := X"00000000";
        ram_buffer(38160) := X"36100001";
        ram_buffer(38161) := X"1000FFAF";
        ram_buffer(38162) := X"00000000";
        ram_buffer(38163) := X"36100002";
        ram_buffer(38164) := X"1000FFAC";
        ram_buffer(38165) := X"00000000";
        ram_buffer(38166) := X"92A30000";
        ram_buffer(38167) := X"24020068";
        ram_buffer(38168) := X"14620005";
        ram_buffer(38169) := X"00000000";
        ram_buffer(38170) := X"26B50001";
        ram_buffer(38171) := X"36100008";
        ram_buffer(38172) := X"1000FFA4";
        ram_buffer(38173) := X"00000000";
        ram_buffer(38174) := X"36100004";
        ram_buffer(38175) := X"1000FFA1";
        ram_buffer(38176) := X"00000000";
        ram_buffer(38177) := X"36100002";
        ram_buffer(38178) := X"1000FF9E";
        ram_buffer(38179) := X"00000000";
        ram_buffer(38180) := X"02401021";
        ram_buffer(38181) := X"00021040";
        ram_buffer(38182) := X"00021880";
        ram_buffer(38183) := X"00431021";
        ram_buffer(38184) := X"02801821";
        ram_buffer(38185) := X"00431021";
        ram_buffer(38186) := X"2452FFD0";
        ram_buffer(38187) := X"1000FF95";
        ram_buffer(38188) := X"00000000";
        ram_buffer(38189) := X"36100001";
        ram_buffer(38190) := X"24140003";
        ram_buffer(38191) := X"3C02100B";
        ram_buffer(38192) := X"24426198";
        ram_buffer(38193) := X"AFC20028";
        ram_buffer(38194) := X"2402000A";
        ram_buffer(38195) := X"AFC20020";
        ram_buffer(38196) := X"100000B2";
        ram_buffer(38197) := X"00000000";
        ram_buffer(38198) := X"24140003";
        ram_buffer(38199) := X"3C02100B";
        ram_buffer(38200) := X"24426198";
        ram_buffer(38201) := X"AFC20028";
        ram_buffer(38202) := X"AFC00020";
        ram_buffer(38203) := X"100000AB";
        ram_buffer(38204) := X"00000000";
        ram_buffer(38205) := X"36100001";
        ram_buffer(38206) := X"24140003";
        ram_buffer(38207) := X"3C02100B";
        ram_buffer(38208) := X"24426A64";
        ram_buffer(38209) := X"AFC20028";
        ram_buffer(38210) := X"24020008";
        ram_buffer(38211) := X"AFC20020";
        ram_buffer(38212) := X"100000A2";
        ram_buffer(38213) := X"00000000";
        ram_buffer(38214) := X"24140003";
        ram_buffer(38215) := X"3C02100B";
        ram_buffer(38216) := X"24426A64";
        ram_buffer(38217) := X"AFC20028";
        ram_buffer(38218) := X"2402000A";
        ram_buffer(38219) := X"AFC20020";
        ram_buffer(38220) := X"1000009A";
        ram_buffer(38221) := X"00000000";
        ram_buffer(38222) := X"36100200";
        ram_buffer(38223) := X"24140003";
        ram_buffer(38224) := X"3C02100B";
        ram_buffer(38225) := X"24426A64";
        ram_buffer(38226) := X"AFC20028";
        ram_buffer(38227) := X"24020010";
        ram_buffer(38228) := X"AFC20020";
        ram_buffer(38229) := X"10000091";
        ram_buffer(38230) := X"00000000";
        ram_buffer(38231) := X"24140004";
        ram_buffer(38232) := X"1000008E";
        ram_buffer(38233) := X"00000000";
        ram_buffer(38234) := X"36100001";
        ram_buffer(38235) := X"24140002";
        ram_buffer(38236) := X"1000008A";
        ram_buffer(38237) := X"00000000";
        ram_buffer(38238) := X"27C200A8";
        ram_buffer(38239) := X"02A02821";
        ram_buffer(38240) := X"00402021";
        ram_buffer(38241) := X"0C02CBBB";
        ram_buffer(38242) := X"00000000";
        ram_buffer(38243) := X"0040A821";
        ram_buffer(38244) := X"36100040";
        ram_buffer(38245) := X"24140001";
        ram_buffer(38246) := X"10000080";
        ram_buffer(38247) := X"00000000";
        ram_buffer(38248) := X"36100001";
        ram_buffer(38249) := X"36100040";
        ram_buffer(38250) := X"0000A021";
        ram_buffer(38251) := X"1000007B";
        ram_buffer(38252) := X"00000000";
        ram_buffer(38253) := X"36100220";
        ram_buffer(38254) := X"24140003";
        ram_buffer(38255) := X"3C02100B";
        ram_buffer(38256) := X"24426A64";
        ram_buffer(38257) := X"AFC20028";
        ram_buffer(38258) := X"24020010";
        ram_buffer(38259) := X"AFC20020";
        ram_buffer(38260) := X"10000072";
        ram_buffer(38261) := X"00000000";
        ram_buffer(38262) := X"32020010";
        ram_buffer(38263) := X"144006AE";
        ram_buffer(38264) := X"00000000";
        ram_buffer(38265) := X"32020008";
        ram_buffer(38266) := X"10400011";
        ram_buffer(38267) := X"00000000";
        ram_buffer(38268) := X"8FC2034C";
        ram_buffer(38269) := X"00000000";
        ram_buffer(38270) := X"24430004";
        ram_buffer(38271) := X"AFC3034C";
        ram_buffer(38272) := X"8C420000";
        ram_buffer(38273) := X"00000000";
        ram_buffer(38274) := X"AFC20068";
        ram_buffer(38275) := X"8FC2001C";
        ram_buffer(38276) := X"00000000";
        ram_buffer(38277) := X"00021E00";
        ram_buffer(38278) := X"00031E03";
        ram_buffer(38279) := X"8FC20068";
        ram_buffer(38280) := X"00000000";
        ram_buffer(38281) := X"A0430000";
        ram_buffer(38282) := X"100006A5";
        ram_buffer(38283) := X"00000000";
        ram_buffer(38284) := X"32020004";
        ram_buffer(38285) := X"10400011";
        ram_buffer(38286) := X"00000000";
        ram_buffer(38287) := X"8FC2034C";
        ram_buffer(38288) := X"00000000";
        ram_buffer(38289) := X"24430004";
        ram_buffer(38290) := X"AFC3034C";
        ram_buffer(38291) := X"8C420000";
        ram_buffer(38292) := X"00000000";
        ram_buffer(38293) := X"AFC2006C";
        ram_buffer(38294) := X"8FC2001C";
        ram_buffer(38295) := X"00000000";
        ram_buffer(38296) := X"00021C00";
        ram_buffer(38297) := X"00031C03";
        ram_buffer(38298) := X"8FC2006C";
        ram_buffer(38299) := X"00000000";
        ram_buffer(38300) := X"A4430000";
        ram_buffer(38301) := X"10000692";
        ram_buffer(38302) := X"00000000";
        ram_buffer(38303) := X"32020001";
        ram_buffer(38304) := X"1040000E";
        ram_buffer(38305) := X"00000000";
        ram_buffer(38306) := X"8FC2034C";
        ram_buffer(38307) := X"00000000";
        ram_buffer(38308) := X"24430004";
        ram_buffer(38309) := X"AFC3034C";
        ram_buffer(38310) := X"8C420000";
        ram_buffer(38311) := X"00000000";
        ram_buffer(38312) := X"AFC20070";
        ram_buffer(38313) := X"8FC20070";
        ram_buffer(38314) := X"8FC3001C";
        ram_buffer(38315) := X"00000000";
        ram_buffer(38316) := X"AC430000";
        ram_buffer(38317) := X"10000682";
        ram_buffer(38318) := X"00000000";
        ram_buffer(38319) := X"32020002";
        ram_buffer(38320) := X"10400013";
        ram_buffer(38321) := X"00000000";
        ram_buffer(38322) := X"8FC2034C";
        ram_buffer(38323) := X"00000000";
        ram_buffer(38324) := X"24430004";
        ram_buffer(38325) := X"AFC3034C";
        ram_buffer(38326) := X"8C420000";
        ram_buffer(38327) := X"00000000";
        ram_buffer(38328) := X"AFC20074";
        ram_buffer(38329) := X"8FC2001C";
        ram_buffer(38330) := X"00000000";
        ram_buffer(38331) := X"0040B821";
        ram_buffer(38332) := X"000217C3";
        ram_buffer(38333) := X"0040B021";
        ram_buffer(38334) := X"8FC20074";
        ram_buffer(38335) := X"00000000";
        ram_buffer(38336) := X"AC570004";
        ram_buffer(38337) := X"AC560000";
        ram_buffer(38338) := X"1000066D";
        ram_buffer(38339) := X"00000000";
        ram_buffer(38340) := X"8FC2034C";
        ram_buffer(38341) := X"00000000";
        ram_buffer(38342) := X"24430004";
        ram_buffer(38343) := X"AFC3034C";
        ram_buffer(38344) := X"8C420000";
        ram_buffer(38345) := X"00000000";
        ram_buffer(38346) := X"AFC20078";
        ram_buffer(38347) := X"8FC20078";
        ram_buffer(38348) := X"8FC3001C";
        ram_buffer(38349) := X"00000000";
        ram_buffer(38350) := X"AC430000";
        ram_buffer(38351) := X"10000660";
        ram_buffer(38352) := X"00000000";
        ram_buffer(38353) := X"2402FFFF";
        ram_buffer(38354) := X"10000690";
        ram_buffer(38355) := X"00000000";
        ram_buffer(38356) := X"8F838090";
        ram_buffer(38357) := X"02801021";
        ram_buffer(38358) := X"24420001";
        ram_buffer(38359) := X"00621021";
        ram_buffer(38360) := X"80420000";
        ram_buffer(38361) := X"00000000";
        ram_buffer(38362) := X"304200FF";
        ram_buffer(38363) := X"30430003";
        ram_buffer(38364) := X"24020001";
        ram_buffer(38365) := X"14620002";
        ram_buffer(38366) := X"00000000";
        ram_buffer(38367) := X"36100001";
        ram_buffer(38368) := X"24140003";
        ram_buffer(38369) := X"3C02100B";
        ram_buffer(38370) := X"24426198";
        ram_buffer(38371) := X"AFC20028";
        ram_buffer(38372) := X"2402000A";
        ram_buffer(38373) := X"AFC20020";
        ram_buffer(38374) := X"00000000";
        ram_buffer(38375) := X"8E220004";
        ram_buffer(38376) := X"00000000";
        ram_buffer(38377) := X"1C400007";
        ram_buffer(38378) := X"00000000";
        ram_buffer(38379) := X"02202821";
        ram_buffer(38380) := X"8FC40340";
        ram_buffer(38381) := X"0C02E477";
        ram_buffer(38382) := X"00000000";
        ram_buffer(38383) := X"14400645";
        ram_buffer(38384) := X"00000000";
        ram_buffer(38385) := X"32020040";
        ram_buffer(38386) := X"14400028";
        ram_buffer(38387) := X"00000000";
        ram_buffer(38388) := X"10000019";
        ram_buffer(38389) := X"00000000";
        ram_buffer(38390) := X"8FC2001C";
        ram_buffer(38391) := X"00000000";
        ram_buffer(38392) := X"24420001";
        ram_buffer(38393) := X"AFC2001C";
        ram_buffer(38394) := X"8E220004";
        ram_buffer(38395) := X"00000000";
        ram_buffer(38396) := X"2442FFFF";
        ram_buffer(38397) := X"AE220004";
        ram_buffer(38398) := X"8E220004";
        ram_buffer(38399) := X"00000000";
        ram_buffer(38400) := X"18400007";
        ram_buffer(38401) := X"00000000";
        ram_buffer(38402) := X"8E220000";
        ram_buffer(38403) := X"00000000";
        ram_buffer(38404) := X"24420001";
        ram_buffer(38405) := X"AE220000";
        ram_buffer(38406) := X"10000007";
        ram_buffer(38407) := X"00000000";
        ram_buffer(38408) := X"02202821";
        ram_buffer(38409) := X"8FC40340";
        ram_buffer(38410) := X"0C02E477";
        ram_buffer(38411) := X"00000000";
        ram_buffer(38412) := X"1440062B";
        ram_buffer(38413) := X"00000000";
        ram_buffer(38414) := X"8F838090";
        ram_buffer(38415) := X"8E220000";
        ram_buffer(38416) := X"00000000";
        ram_buffer(38417) := X"90420000";
        ram_buffer(38418) := X"00000000";
        ram_buffer(38419) := X"24420001";
        ram_buffer(38420) := X"00621021";
        ram_buffer(38421) := X"80420000";
        ram_buffer(38422) := X"00000000";
        ram_buffer(38423) := X"304200FF";
        ram_buffer(38424) := X"30420008";
        ram_buffer(38425) := X"1440FFDC";
        ram_buffer(38426) := X"00000000";
        ram_buffer(38427) := X"2E820005";
        ram_buffer(38428) := X"1040FE60";
        ram_buffer(38429) := X"00000000";
        ram_buffer(38430) := X"00141880";
        ram_buffer(38431) := X"3C02100D";
        ram_buffer(38432) := X"2442A458";
        ram_buffer(38433) := X"00621021";
        ram_buffer(38434) := X"8C420000";
        ram_buffer(38435) := X"00000000";
        ram_buffer(38436) := X"00400008";
        ram_buffer(38437) := X"00000000";
        ram_buffer(38438) := X"16400002";
        ram_buffer(38439) := X"00000000";
        ram_buffer(38440) := X"24120001";
        ram_buffer(38441) := X"32020001";
        ram_buffer(38442) := X"10400074";
        ram_buffer(38443) := X"00000000";
        ram_buffer(38444) := X"27C20308";
        ram_buffer(38445) := X"24060008";
        ram_buffer(38446) := X"00002821";
        ram_buffer(38447) := X"00402021";
        ram_buffer(38448) := X"0C02801D";
        ram_buffer(38449) := X"00000000";
        ram_buffer(38450) := X"32020010";
        ram_buffer(38451) := X"1440000A";
        ram_buffer(38452) := X"00000000";
        ram_buffer(38453) := X"8FC2034C";
        ram_buffer(38454) := X"00000000";
        ram_buffer(38455) := X"24430004";
        ram_buffer(38456) := X"AFC3034C";
        ram_buffer(38457) := X"8C420000";
        ram_buffer(38458) := X"00000000";
        ram_buffer(38459) := X"AFC20024";
        ram_buffer(38460) := X"10000002";
        ram_buffer(38461) := X"00000000";
        ram_buffer(38462) := X"AFC00024";
        ram_buffer(38463) := X"0000A021";
        ram_buffer(38464) := X"10000050";
        ram_buffer(38465) := X"00000000";
        ram_buffer(38466) := X"0C02BB09";
        ram_buffer(38467) := X"00000000";
        ram_buffer(38468) := X"105405F6";
        ram_buffer(38469) := X"00000000";
        ram_buffer(38470) := X"02801021";
        ram_buffer(38471) := X"24540001";
        ram_buffer(38472) := X"8E230000";
        ram_buffer(38473) := X"00000000";
        ram_buffer(38474) := X"90630000";
        ram_buffer(38475) := X"00000000";
        ram_buffer(38476) := X"00031E00";
        ram_buffer(38477) := X"00031E03";
        ram_buffer(38478) := X"27C40018";
        ram_buffer(38479) := X"00821021";
        ram_buffer(38480) := X"A0430190";
        ram_buffer(38481) := X"8E220004";
        ram_buffer(38482) := X"00000000";
        ram_buffer(38483) := X"2442FFFF";
        ram_buffer(38484) := X"AE220004";
        ram_buffer(38485) := X"8E220000";
        ram_buffer(38486) := X"00000000";
        ram_buffer(38487) := X"24420001";
        ram_buffer(38488) := X"AE220000";
        ram_buffer(38489) := X"02802021";
        ram_buffer(38490) := X"27C301A8";
        ram_buffer(38491) := X"27C20308";
        ram_buffer(38492) := X"AFA20010";
        ram_buffer(38493) := X"00803821";
        ram_buffer(38494) := X"00603021";
        ram_buffer(38495) := X"8FC50024";
        ram_buffer(38496) := X"8FC40340";
        ram_buffer(38497) := X"0C02BB73";
        ram_buffer(38498) := X"00000000";
        ram_buffer(38499) := X"AFC2007C";
        ram_buffer(38500) := X"8FC3007C";
        ram_buffer(38501) := X"2402FFFF";
        ram_buffer(38502) := X"106205D7";
        ram_buffer(38503) := X"00000000";
        ram_buffer(38504) := X"8FC2007C";
        ram_buffer(38505) := X"00000000";
        ram_buffer(38506) := X"14400007";
        ram_buffer(38507) := X"00000000";
        ram_buffer(38508) := X"32020010";
        ram_buffer(38509) := X"14400004";
        ram_buffer(38510) := X"00000000";
        ram_buffer(38511) := X"8FC20024";
        ram_buffer(38512) := X"00000000";
        ram_buffer(38513) := X"AC400000";
        ram_buffer(38514) := X"8FC3007C";
        ram_buffer(38515) := X"2402FFFE";
        ram_buffer(38516) := X"1062000E";
        ram_buffer(38517) := X"00000000";
        ram_buffer(38518) := X"8FC2001C";
        ram_buffer(38519) := X"00000000";
        ram_buffer(38520) := X"00541021";
        ram_buffer(38521) := X"AFC2001C";
        ram_buffer(38522) := X"2652FFFF";
        ram_buffer(38523) := X"32020010";
        ram_buffer(38524) := X"14400005";
        ram_buffer(38525) := X"00000000";
        ram_buffer(38526) := X"8FC20024";
        ram_buffer(38527) := X"00000000";
        ram_buffer(38528) := X"24420004";
        ram_buffer(38529) := X"AFC20024";
        ram_buffer(38530) := X"0000A021";
        ram_buffer(38531) := X"8E220004";
        ram_buffer(38532) := X"00000000";
        ram_buffer(38533) := X"1C40000B";
        ram_buffer(38534) := X"00000000";
        ram_buffer(38535) := X"02202821";
        ram_buffer(38536) := X"8FC40340";
        ram_buffer(38537) := X"0C02E477";
        ram_buffer(38538) := X"00000000";
        ram_buffer(38539) := X"10400005";
        ram_buffer(38540) := X"00000000";
        ram_buffer(38541) := X"12800007";
        ram_buffer(38542) := X"00000000";
        ram_buffer(38543) := X"100005B8";
        ram_buffer(38544) := X"00000000";
        ram_buffer(38545) := X"1640FFB0";
        ram_buffer(38546) := X"00000000";
        ram_buffer(38547) := X"10000002";
        ram_buffer(38548) := X"00000000";
        ram_buffer(38549) := X"00000000";
        ram_buffer(38550) := X"32020010";
        ram_buffer(38551) := X"14400591";
        ram_buffer(38552) := X"00000000";
        ram_buffer(38553) := X"8FC20018";
        ram_buffer(38554) := X"00000000";
        ram_buffer(38555) := X"24420001";
        ram_buffer(38556) := X"AFC20018";
        ram_buffer(38557) := X"1000058B";
        ram_buffer(38558) := X"00000000";
        ram_buffer(38559) := X"32020010";
        ram_buffer(38560) := X"10400034";
        ram_buffer(38561) := X"00000000";
        ram_buffer(38562) := X"AFC00030";
        ram_buffer(38563) := X"8E340004";
        ram_buffer(38564) := X"02401021";
        ram_buffer(38565) := X"0282102A";
        ram_buffer(38566) := X"10400018";
        ram_buffer(38567) := X"00000000";
        ram_buffer(38568) := X"02801821";
        ram_buffer(38569) := X"8FC20030";
        ram_buffer(38570) := X"00000000";
        ram_buffer(38571) := X"00431021";
        ram_buffer(38572) := X"AFC20030";
        ram_buffer(38573) := X"02801021";
        ram_buffer(38574) := X"02429023";
        ram_buffer(38575) := X"8E220000";
        ram_buffer(38576) := X"02801821";
        ram_buffer(38577) := X"00431021";
        ram_buffer(38578) := X"AE220000";
        ram_buffer(38579) := X"02202821";
        ram_buffer(38580) := X"8FC40340";
        ram_buffer(38581) := X"0C02E477";
        ram_buffer(38582) := X"00000000";
        ram_buffer(38583) := X"1040FFEB";
        ram_buffer(38584) := X"00000000";
        ram_buffer(38585) := X"8FC20030";
        ram_buffer(38586) := X"00000000";
        ram_buffer(38587) := X"14400011";
        ram_buffer(38588) := X"00000000";
        ram_buffer(38589) := X"1000058A";
        ram_buffer(38590) := X"00000000";
        ram_buffer(38591) := X"8FC20030";
        ram_buffer(38592) := X"00000000";
        ram_buffer(38593) := X"00521021";
        ram_buffer(38594) := X"AFC20030";
        ram_buffer(38595) := X"8E220004";
        ram_buffer(38596) := X"00000000";
        ram_buffer(38597) := X"00521023";
        ram_buffer(38598) := X"AE220004";
        ram_buffer(38599) := X"8E220000";
        ram_buffer(38600) := X"00000000";
        ram_buffer(38601) := X"00521021";
        ram_buffer(38602) := X"AE220000";
        ram_buffer(38603) := X"10000002";
        ram_buffer(38604) := X"00000000";
        ram_buffer(38605) := X"00000000";
        ram_buffer(38606) := X"8FC3001C";
        ram_buffer(38607) := X"8FC20030";
        ram_buffer(38608) := X"00000000";
        ram_buffer(38609) := X"00621021";
        ram_buffer(38610) := X"AFC2001C";
        ram_buffer(38611) := X"10000555";
        ram_buffer(38612) := X"00000000";
        ram_buffer(38613) := X"8FC2034C";
        ram_buffer(38614) := X"00000000";
        ram_buffer(38615) := X"24430004";
        ram_buffer(38616) := X"AFC3034C";
        ram_buffer(38617) := X"8C420000";
        ram_buffer(38618) := X"AFB10010";
        ram_buffer(38619) := X"02403821";
        ram_buffer(38620) := X"24060001";
        ram_buffer(38621) := X"00402821";
        ram_buffer(38622) := X"8FC40340";
        ram_buffer(38623) := X"0C02E4AC";
        ram_buffer(38624) := X"00000000";
        ram_buffer(38625) := X"AFC20080";
        ram_buffer(38626) := X"8FC20080";
        ram_buffer(38627) := X"00000000";
        ram_buffer(38628) := X"1040055C";
        ram_buffer(38629) := X"00000000";
        ram_buffer(38630) := X"8FC3001C";
        ram_buffer(38631) := X"8FC20080";
        ram_buffer(38632) := X"00000000";
        ram_buffer(38633) := X"00621021";
        ram_buffer(38634) := X"AFC2001C";
        ram_buffer(38635) := X"8FC20018";
        ram_buffer(38636) := X"00000000";
        ram_buffer(38637) := X"24420001";
        ram_buffer(38638) := X"AFC20018";
        ram_buffer(38639) := X"10000539";
        ram_buffer(38640) := X"00000000";
        ram_buffer(38641) := X"16400002";
        ram_buffer(38642) := X"00000000";
        ram_buffer(38643) := X"2412FFFF";
        ram_buffer(38644) := X"32020010";
        ram_buffer(38645) := X"10400033";
        ram_buffer(38646) := X"00000000";
        ram_buffer(38647) := X"0000A021";
        ram_buffer(38648) := X"1000001B";
        ram_buffer(38649) := X"00000000";
        ram_buffer(38650) := X"26940001";
        ram_buffer(38651) := X"8E220004";
        ram_buffer(38652) := X"00000000";
        ram_buffer(38653) := X"2442FFFF";
        ram_buffer(38654) := X"AE220004";
        ram_buffer(38655) := X"8E220000";
        ram_buffer(38656) := X"00000000";
        ram_buffer(38657) := X"24420001";
        ram_buffer(38658) := X"AE220000";
        ram_buffer(38659) := X"2652FFFF";
        ram_buffer(38660) := X"1240001C";
        ram_buffer(38661) := X"00000000";
        ram_buffer(38662) := X"8E220004";
        ram_buffer(38663) := X"00000000";
        ram_buffer(38664) := X"1C40000B";
        ram_buffer(38665) := X"00000000";
        ram_buffer(38666) := X"02202821";
        ram_buffer(38667) := X"8FC40340";
        ram_buffer(38668) := X"0C02E477";
        ram_buffer(38669) := X"00000000";
        ram_buffer(38670) := X"10400005";
        ram_buffer(38671) := X"00000000";
        ram_buffer(38672) := X"16800013";
        ram_buffer(38673) := X"00000000";
        ram_buffer(38674) := X"10000535";
        ram_buffer(38675) := X"00000000";
        ram_buffer(38676) := X"8E220000";
        ram_buffer(38677) := X"00000000";
        ram_buffer(38678) := X"90420000";
        ram_buffer(38679) := X"00000000";
        ram_buffer(38680) := X"00401821";
        ram_buffer(38681) := X"27C20018";
        ram_buffer(38682) := X"00431021";
        ram_buffer(38683) := X"80420090";
        ram_buffer(38684) := X"00000000";
        ram_buffer(38685) := X"1440FFDC";
        ram_buffer(38686) := X"00000000";
        ram_buffer(38687) := X"10000005";
        ram_buffer(38688) := X"00000000";
        ram_buffer(38689) := X"00000000";
        ram_buffer(38690) := X"10000002";
        ram_buffer(38691) := X"00000000";
        ram_buffer(38692) := X"00000000";
        ram_buffer(38693) := X"16800047";
        ram_buffer(38694) := X"00000000";
        ram_buffer(38695) := X"1000053A";
        ram_buffer(38696) := X"00000000";
        ram_buffer(38697) := X"8FC2034C";
        ram_buffer(38698) := X"00000000";
        ram_buffer(38699) := X"24430004";
        ram_buffer(38700) := X"AFC3034C";
        ram_buffer(38701) := X"8C530000";
        ram_buffer(38702) := X"00000000";
        ram_buffer(38703) := X"02608021";
        ram_buffer(38704) := X"10000021";
        ram_buffer(38705) := X"00000000";
        ram_buffer(38706) := X"8E220004";
        ram_buffer(38707) := X"00000000";
        ram_buffer(38708) := X"2442FFFF";
        ram_buffer(38709) := X"AE220004";
        ram_buffer(38710) := X"02601821";
        ram_buffer(38711) := X"24730001";
        ram_buffer(38712) := X"8E220000";
        ram_buffer(38713) := X"00000000";
        ram_buffer(38714) := X"24440001";
        ram_buffer(38715) := X"AE240000";
        ram_buffer(38716) := X"90420000";
        ram_buffer(38717) := X"00000000";
        ram_buffer(38718) := X"00021600";
        ram_buffer(38719) := X"00021603";
        ram_buffer(38720) := X"A0620000";
        ram_buffer(38721) := X"2652FFFF";
        ram_buffer(38722) := X"1240001C";
        ram_buffer(38723) := X"00000000";
        ram_buffer(38724) := X"8E220004";
        ram_buffer(38725) := X"00000000";
        ram_buffer(38726) := X"1C40000B";
        ram_buffer(38727) := X"00000000";
        ram_buffer(38728) := X"02202821";
        ram_buffer(38729) := X"8FC40340";
        ram_buffer(38730) := X"0C02E477";
        ram_buffer(38731) := X"00000000";
        ram_buffer(38732) := X"10400005";
        ram_buffer(38733) := X"00000000";
        ram_buffer(38734) := X"16700013";
        ram_buffer(38735) := X"00000000";
        ram_buffer(38736) := X"100004F7";
        ram_buffer(38737) := X"00000000";
        ram_buffer(38738) := X"8E220000";
        ram_buffer(38739) := X"00000000";
        ram_buffer(38740) := X"90420000";
        ram_buffer(38741) := X"00000000";
        ram_buffer(38742) := X"00401821";
        ram_buffer(38743) := X"27C20018";
        ram_buffer(38744) := X"00431021";
        ram_buffer(38745) := X"80420090";
        ram_buffer(38746) := X"00000000";
        ram_buffer(38747) := X"1440FFD6";
        ram_buffer(38748) := X"00000000";
        ram_buffer(38749) := X"10000005";
        ram_buffer(38750) := X"00000000";
        ram_buffer(38751) := X"00000000";
        ram_buffer(38752) := X"10000002";
        ram_buffer(38753) := X"00000000";
        ram_buffer(38754) := X"00000000";
        ram_buffer(38755) := X"02601821";
        ram_buffer(38756) := X"02001021";
        ram_buffer(38757) := X"0062A023";
        ram_buffer(38758) := X"128004F7";
        ram_buffer(38759) := X"00000000";
        ram_buffer(38760) := X"A2600000";
        ram_buffer(38761) := X"8FC20018";
        ram_buffer(38762) := X"00000000";
        ram_buffer(38763) := X"24420001";
        ram_buffer(38764) := X"AFC20018";
        ram_buffer(38765) := X"8FC2001C";
        ram_buffer(38766) := X"00000000";
        ram_buffer(38767) := X"00541021";
        ram_buffer(38768) := X"AFC2001C";
        ram_buffer(38769) := X"100004BE";
        ram_buffer(38770) := X"00000000";
        ram_buffer(38771) := X"16400002";
        ram_buffer(38772) := X"00000000";
        ram_buffer(38773) := X"2412FFFF";
        ram_buffer(38774) := X"32020001";
        ram_buffer(38775) := X"1040009C";
        ram_buffer(38776) := X"00000000";
        ram_buffer(38777) := X"27C20310";
        ram_buffer(38778) := X"24060008";
        ram_buffer(38779) := X"00002821";
        ram_buffer(38780) := X"00402021";
        ram_buffer(38781) := X"0C02801D";
        ram_buffer(38782) := X"00000000";
        ram_buffer(38783) := X"32020010";
        ram_buffer(38784) := X"1440000A";
        ram_buffer(38785) := X"00000000";
        ram_buffer(38786) := X"8FC2034C";
        ram_buffer(38787) := X"00000000";
        ram_buffer(38788) := X"24430004";
        ram_buffer(38789) := X"AFC3034C";
        ram_buffer(38790) := X"8C420000";
        ram_buffer(38791) := X"00000000";
        ram_buffer(38792) := X"AFC20024";
        ram_buffer(38793) := X"10000003";
        ram_buffer(38794) := X"00000000";
        ram_buffer(38795) := X"27C200A4";
        ram_buffer(38796) := X"AFC20024";
        ram_buffer(38797) := X"0000A021";
        ram_buffer(38798) := X"10000067";
        ram_buffer(38799) := X"00000000";
        ram_buffer(38800) := X"0C02BB09";
        ram_buffer(38801) := X"00000000";
        ram_buffer(38802) := X"105404B1";
        ram_buffer(38803) := X"00000000";
        ram_buffer(38804) := X"02801021";
        ram_buffer(38805) := X"24540001";
        ram_buffer(38806) := X"8E230000";
        ram_buffer(38807) := X"00000000";
        ram_buffer(38808) := X"90630000";
        ram_buffer(38809) := X"00000000";
        ram_buffer(38810) := X"00031E00";
        ram_buffer(38811) := X"00031E03";
        ram_buffer(38812) := X"27C40018";
        ram_buffer(38813) := X"00821021";
        ram_buffer(38814) := X"A0430190";
        ram_buffer(38815) := X"8E220004";
        ram_buffer(38816) := X"00000000";
        ram_buffer(38817) := X"2442FFFF";
        ram_buffer(38818) := X"AE220004";
        ram_buffer(38819) := X"8E220000";
        ram_buffer(38820) := X"00000000";
        ram_buffer(38821) := X"24420001";
        ram_buffer(38822) := X"AE220000";
        ram_buffer(38823) := X"02802021";
        ram_buffer(38824) := X"27C301A8";
        ram_buffer(38825) := X"27C20310";
        ram_buffer(38826) := X"AFA20010";
        ram_buffer(38827) := X"00803821";
        ram_buffer(38828) := X"00603021";
        ram_buffer(38829) := X"8FC50024";
        ram_buffer(38830) := X"8FC40340";
        ram_buffer(38831) := X"0C02BB73";
        ram_buffer(38832) := X"00000000";
        ram_buffer(38833) := X"AFC2007C";
        ram_buffer(38834) := X"8FC3007C";
        ram_buffer(38835) := X"2402FFFF";
        ram_buffer(38836) := X"10620492";
        ram_buffer(38837) := X"00000000";
        ram_buffer(38838) := X"8FC2007C";
        ram_buffer(38839) := X"00000000";
        ram_buffer(38840) := X"14400004";
        ram_buffer(38841) := X"00000000";
        ram_buffer(38842) := X"8FC20024";
        ram_buffer(38843) := X"00000000";
        ram_buffer(38844) := X"AC400000";
        ram_buffer(38845) := X"8FC3007C";
        ram_buffer(38846) := X"2402FFFE";
        ram_buffer(38847) := X"10620028";
        ram_buffer(38848) := X"00000000";
        ram_buffer(38849) := X"8FC20024";
        ram_buffer(38850) := X"00000000";
        ram_buffer(38851) := X"8C420000";
        ram_buffer(38852) := X"00000000";
        ram_buffer(38853) := X"00402021";
        ram_buffer(38854) := X"0C02BABA";
        ram_buffer(38855) := X"00000000";
        ram_buffer(38856) := X"10400012";
        ram_buffer(38857) := X"00000000";
        ram_buffer(38858) := X"1000000C";
        ram_buffer(38859) := X"00000000";
        ram_buffer(38860) := X"2694FFFF";
        ram_buffer(38861) := X"27C20018";
        ram_buffer(38862) := X"00541021";
        ram_buffer(38863) := X"80420190";
        ram_buffer(38864) := X"00000000";
        ram_buffer(38865) := X"304200FF";
        ram_buffer(38866) := X"02203021";
        ram_buffer(38867) := X"00402821";
        ram_buffer(38868) := X"8FC40340";
        ram_buffer(38869) := X"0C02E402";
        ram_buffer(38870) := X"00000000";
        ram_buffer(38871) := X"1680FFF4";
        ram_buffer(38872) := X"00000000";
        ram_buffer(38873) := X"1000002E";
        ram_buffer(38874) := X"00000000";
        ram_buffer(38875) := X"8FC2001C";
        ram_buffer(38876) := X"00000000";
        ram_buffer(38877) := X"00541021";
        ram_buffer(38878) := X"AFC2001C";
        ram_buffer(38879) := X"2652FFFF";
        ram_buffer(38880) := X"32020010";
        ram_buffer(38881) := X"14400005";
        ram_buffer(38882) := X"00000000";
        ram_buffer(38883) := X"8FC20024";
        ram_buffer(38884) := X"00000000";
        ram_buffer(38885) := X"24420004";
        ram_buffer(38886) := X"AFC20024";
        ram_buffer(38887) := X"0000A021";
        ram_buffer(38888) := X"8E220004";
        ram_buffer(38889) := X"00000000";
        ram_buffer(38890) := X"1C40000B";
        ram_buffer(38891) := X"00000000";
        ram_buffer(38892) := X"02202821";
        ram_buffer(38893) := X"8FC40340";
        ram_buffer(38894) := X"0C02E477";
        ram_buffer(38895) := X"00000000";
        ram_buffer(38896) := X"10400005";
        ram_buffer(38897) := X"00000000";
        ram_buffer(38898) := X"12800014";
        ram_buffer(38899) := X"00000000";
        ram_buffer(38900) := X"10000453";
        ram_buffer(38901) := X"00000000";
        ram_buffer(38902) := X"8F838090";
        ram_buffer(38903) := X"8E220000";
        ram_buffer(38904) := X"00000000";
        ram_buffer(38905) := X"90420000";
        ram_buffer(38906) := X"00000000";
        ram_buffer(38907) := X"24420001";
        ram_buffer(38908) := X"00621021";
        ram_buffer(38909) := X"80420000";
        ram_buffer(38910) := X"00000000";
        ram_buffer(38911) := X"304200FF";
        ram_buffer(38912) := X"30420008";
        ram_buffer(38913) := X"14400006";
        ram_buffer(38914) := X"00000000";
        ram_buffer(38915) := X"1640FF8C";
        ram_buffer(38916) := X"00000000";
        ram_buffer(38917) := X"10000002";
        ram_buffer(38918) := X"00000000";
        ram_buffer(38919) := X"00000000";
        ram_buffer(38920) := X"32020010";
        ram_buffer(38921) := X"14400422";
        ram_buffer(38922) := X"00000000";
        ram_buffer(38923) := X"8FC20024";
        ram_buffer(38924) := X"00000000";
        ram_buffer(38925) := X"AC400000";
        ram_buffer(38926) := X"8FC20018";
        ram_buffer(38927) := X"00000000";
        ram_buffer(38928) := X"24420001";
        ram_buffer(38929) := X"AFC20018";
        ram_buffer(38930) := X"10000419";
        ram_buffer(38931) := X"00000000";
        ram_buffer(38932) := X"32020010";
        ram_buffer(38933) := X"10400033";
        ram_buffer(38934) := X"00000000";
        ram_buffer(38935) := X"0000A021";
        ram_buffer(38936) := X"10000017";
        ram_buffer(38937) := X"00000000";
        ram_buffer(38938) := X"26940001";
        ram_buffer(38939) := X"8E220004";
        ram_buffer(38940) := X"00000000";
        ram_buffer(38941) := X"2442FFFF";
        ram_buffer(38942) := X"AE220004";
        ram_buffer(38943) := X"8E220000";
        ram_buffer(38944) := X"00000000";
        ram_buffer(38945) := X"24420001";
        ram_buffer(38946) := X"AE220000";
        ram_buffer(38947) := X"2652FFFF";
        ram_buffer(38948) := X"1240001A";
        ram_buffer(38949) := X"00000000";
        ram_buffer(38950) := X"8E220004";
        ram_buffer(38951) := X"00000000";
        ram_buffer(38952) := X"1C400007";
        ram_buffer(38953) := X"00000000";
        ram_buffer(38954) := X"02202821";
        ram_buffer(38955) := X"8FC40340";
        ram_buffer(38956) := X"0C02E477";
        ram_buffer(38957) := X"00000000";
        ram_buffer(38958) := X"14400013";
        ram_buffer(38959) := X"00000000";
        ram_buffer(38960) := X"8F838090";
        ram_buffer(38961) := X"8E220000";
        ram_buffer(38962) := X"00000000";
        ram_buffer(38963) := X"90420000";
        ram_buffer(38964) := X"00000000";
        ram_buffer(38965) := X"24420001";
        ram_buffer(38966) := X"00621021";
        ram_buffer(38967) := X"80420000";
        ram_buffer(38968) := X"00000000";
        ram_buffer(38969) := X"304200FF";
        ram_buffer(38970) := X"30420008";
        ram_buffer(38971) := X"1040FFDE";
        ram_buffer(38972) := X"00000000";
        ram_buffer(38973) := X"10000005";
        ram_buffer(38974) := X"00000000";
        ram_buffer(38975) := X"00000000";
        ram_buffer(38976) := X"10000002";
        ram_buffer(38977) := X"00000000";
        ram_buffer(38978) := X"00000000";
        ram_buffer(38979) := X"8FC2001C";
        ram_buffer(38980) := X"00000000";
        ram_buffer(38981) := X"00541021";
        ram_buffer(38982) := X"AFC2001C";
        ram_buffer(38983) := X"100003E4";
        ram_buffer(38984) := X"00000000";
        ram_buffer(38985) := X"8FC2034C";
        ram_buffer(38986) := X"00000000";
        ram_buffer(38987) := X"24430004";
        ram_buffer(38988) := X"AFC3034C";
        ram_buffer(38989) := X"8C530000";
        ram_buffer(38990) := X"00000000";
        ram_buffer(38991) := X"02608021";
        ram_buffer(38992) := X"1000001D";
        ram_buffer(38993) := X"00000000";
        ram_buffer(38994) := X"8E220004";
        ram_buffer(38995) := X"00000000";
        ram_buffer(38996) := X"2442FFFF";
        ram_buffer(38997) := X"AE220004";
        ram_buffer(38998) := X"02601821";
        ram_buffer(38999) := X"24730001";
        ram_buffer(39000) := X"8E220000";
        ram_buffer(39001) := X"00000000";
        ram_buffer(39002) := X"24440001";
        ram_buffer(39003) := X"AE240000";
        ram_buffer(39004) := X"90420000";
        ram_buffer(39005) := X"00000000";
        ram_buffer(39006) := X"00021600";
        ram_buffer(39007) := X"00021603";
        ram_buffer(39008) := X"A0620000";
        ram_buffer(39009) := X"2652FFFF";
        ram_buffer(39010) := X"1240001A";
        ram_buffer(39011) := X"00000000";
        ram_buffer(39012) := X"8E220004";
        ram_buffer(39013) := X"00000000";
        ram_buffer(39014) := X"1C400007";
        ram_buffer(39015) := X"00000000";
        ram_buffer(39016) := X"02202821";
        ram_buffer(39017) := X"8FC40340";
        ram_buffer(39018) := X"0C02E477";
        ram_buffer(39019) := X"00000000";
        ram_buffer(39020) := X"14400013";
        ram_buffer(39021) := X"00000000";
        ram_buffer(39022) := X"8F838090";
        ram_buffer(39023) := X"8E220000";
        ram_buffer(39024) := X"00000000";
        ram_buffer(39025) := X"90420000";
        ram_buffer(39026) := X"00000000";
        ram_buffer(39027) := X"24420001";
        ram_buffer(39028) := X"00621021";
        ram_buffer(39029) := X"80420000";
        ram_buffer(39030) := X"00000000";
        ram_buffer(39031) := X"304200FF";
        ram_buffer(39032) := X"30420008";
        ram_buffer(39033) := X"1040FFD8";
        ram_buffer(39034) := X"00000000";
        ram_buffer(39035) := X"10000005";
        ram_buffer(39036) := X"00000000";
        ram_buffer(39037) := X"00000000";
        ram_buffer(39038) := X"10000002";
        ram_buffer(39039) := X"00000000";
        ram_buffer(39040) := X"00000000";
        ram_buffer(39041) := X"A2600000";
        ram_buffer(39042) := X"02601821";
        ram_buffer(39043) := X"02001021";
        ram_buffer(39044) := X"00621023";
        ram_buffer(39045) := X"8FC3001C";
        ram_buffer(39046) := X"00000000";
        ram_buffer(39047) := X"00621021";
        ram_buffer(39048) := X"AFC2001C";
        ram_buffer(39049) := X"8FC20018";
        ram_buffer(39050) := X"00000000";
        ram_buffer(39051) := X"24420001";
        ram_buffer(39052) := X"AFC20018";
        ram_buffer(39053) := X"1000039E";
        ram_buffer(39054) := X"00000000";
        ram_buffer(39055) := X"AFC00034";
        ram_buffer(39056) := X"AFC00038";
        ram_buffer(39057) := X"2642FFFF";
        ram_buffer(39058) := X"2C42015D";
        ram_buffer(39059) := X"14400004";
        ram_buffer(39060) := X"00000000";
        ram_buffer(39061) := X"2642FEA3";
        ram_buffer(39062) := X"AFC20034";
        ram_buffer(39063) := X"2412015D";
        ram_buffer(39064) := X"36100D80";
        ram_buffer(39065) := X"27D301A8";
        ram_buffer(39066) := X"10000095";
        ram_buffer(39067) := X"00000000";
        ram_buffer(39068) := X"8E220000";
        ram_buffer(39069) := X"00000000";
        ram_buffer(39070) := X"90420000";
        ram_buffer(39071) := X"00000000";
        ram_buffer(39072) := X"0040A021";
        ram_buffer(39073) := X"2682FFD5";
        ram_buffer(39074) := X"2C43004E";
        ram_buffer(39075) := X"10600090";
        ram_buffer(39076) := X"00000000";
        ram_buffer(39077) := X"00021880";
        ram_buffer(39078) := X"3C02100D";
        ram_buffer(39079) := X"2442A46C";
        ram_buffer(39080) := X"00621021";
        ram_buffer(39081) := X"8C420000";
        ram_buffer(39082) := X"00000000";
        ram_buffer(39083) := X"00400008";
        ram_buffer(39084) := X"00000000";
        ram_buffer(39085) := X"32020800";
        ram_buffer(39086) := X"10400066";
        ram_buffer(39087) := X"00000000";
        ram_buffer(39088) := X"8FC20020";
        ram_buffer(39089) := X"00000000";
        ram_buffer(39090) := X"14400004";
        ram_buffer(39091) := X"00000000";
        ram_buffer(39092) := X"24020008";
        ram_buffer(39093) := X"AFC20020";
        ram_buffer(39094) := X"36100200";
        ram_buffer(39095) := X"32020400";
        ram_buffer(39096) := X"10400005";
        ram_buffer(39097) := X"00000000";
        ram_buffer(39098) := X"2402FA7F";
        ram_buffer(39099) := X"02028024";
        ram_buffer(39100) := X"10000059";
        ram_buffer(39101) := X"00000000";
        ram_buffer(39102) := X"2402FC7F";
        ram_buffer(39103) := X"02028024";
        ram_buffer(39104) := X"8FC20034";
        ram_buffer(39105) := X"00000000";
        ram_buffer(39106) := X"10400006";
        ram_buffer(39107) := X"00000000";
        ram_buffer(39108) := X"8FC20034";
        ram_buffer(39109) := X"00000000";
        ram_buffer(39110) := X"2442FFFF";
        ram_buffer(39111) := X"AFC20034";
        ram_buffer(39112) := X"26520001";
        ram_buffer(39113) := X"8FC20038";
        ram_buffer(39114) := X"00000000";
        ram_buffer(39115) := X"24420001";
        ram_buffer(39116) := X"AFC20038";
        ram_buffer(39117) := X"1000004D";
        ram_buffer(39118) := X"00000000";
        ram_buffer(39119) := X"3C02100D";
        ram_buffer(39120) := X"8FC30020";
        ram_buffer(39121) := X"00000000";
        ram_buffer(39122) := X"00031840";
        ram_buffer(39123) := X"2442A6E0";
        ram_buffer(39124) := X"00621021";
        ram_buffer(39125) := X"84420000";
        ram_buffer(39126) := X"00000000";
        ram_buffer(39127) := X"AFC20020";
        ram_buffer(39128) := X"2402F47F";
        ram_buffer(39129) := X"02028024";
        ram_buffer(39130) := X"1000003B";
        ram_buffer(39131) := X"00000000";
        ram_buffer(39132) := X"3C02100D";
        ram_buffer(39133) := X"8FC30020";
        ram_buffer(39134) := X"00000000";
        ram_buffer(39135) := X"00031840";
        ram_buffer(39136) := X"2442A6E0";
        ram_buffer(39137) := X"00621021";
        ram_buffer(39138) := X"84420000";
        ram_buffer(39139) := X"00000000";
        ram_buffer(39140) := X"AFC20020";
        ram_buffer(39141) := X"8FC20020";
        ram_buffer(39142) := X"00000000";
        ram_buffer(39143) := X"28420009";
        ram_buffer(39144) := X"14400020";
        ram_buffer(39145) := X"00000000";
        ram_buffer(39146) := X"2402F47F";
        ram_buffer(39147) := X"02028024";
        ram_buffer(39148) := X"10000029";
        ram_buffer(39149) := X"00000000";
        ram_buffer(39150) := X"8FC20020";
        ram_buffer(39151) := X"00000000";
        ram_buffer(39152) := X"2842000B";
        ram_buffer(39153) := X"1440001A";
        ram_buffer(39154) := X"00000000";
        ram_buffer(39155) := X"2402F47F";
        ram_buffer(39156) := X"02028024";
        ram_buffer(39157) := X"10000020";
        ram_buffer(39158) := X"00000000";
        ram_buffer(39159) := X"32020080";
        ram_buffer(39160) := X"10400016";
        ram_buffer(39161) := X"00000000";
        ram_buffer(39162) := X"2402FF7F";
        ram_buffer(39163) := X"02028024";
        ram_buffer(39164) := X"10000019";
        ram_buffer(39165) := X"00000000";
        ram_buffer(39166) := X"32030600";
        ram_buffer(39167) := X"24020200";
        ram_buffer(39168) := X"14620011";
        ram_buffer(39169) := X"00000000";
        ram_buffer(39170) := X"24020010";
        ram_buffer(39171) := X"AFC20020";
        ram_buffer(39172) := X"2402FDFF";
        ram_buffer(39173) := X"02028024";
        ram_buffer(39174) := X"36100500";
        ram_buffer(39175) := X"1000000E";
        ram_buffer(39176) := X"00000000";
        ram_buffer(39177) := X"00000000";
        ram_buffer(39178) := X"10000029";
        ram_buffer(39179) := X"00000000";
        ram_buffer(39180) := X"00000000";
        ram_buffer(39181) := X"10000026";
        ram_buffer(39182) := X"00000000";
        ram_buffer(39183) := X"00000000";
        ram_buffer(39184) := X"10000023";
        ram_buffer(39185) := X"00000000";
        ram_buffer(39186) := X"00000000";
        ram_buffer(39187) := X"10000020";
        ram_buffer(39188) := X"00000000";
        ram_buffer(39189) := X"00000000";
        ram_buffer(39190) := X"02601021";
        ram_buffer(39191) := X"24530001";
        ram_buffer(39192) := X"00141E00";
        ram_buffer(39193) := X"00031E03";
        ram_buffer(39194) := X"A0430000";
        ram_buffer(39195) := X"8E220004";
        ram_buffer(39196) := X"00000000";
        ram_buffer(39197) := X"2442FFFF";
        ram_buffer(39198) := X"AE220004";
        ram_buffer(39199) := X"8E220004";
        ram_buffer(39200) := X"00000000";
        ram_buffer(39201) := X"18400007";
        ram_buffer(39202) := X"00000000";
        ram_buffer(39203) := X"8E220000";
        ram_buffer(39204) := X"00000000";
        ram_buffer(39205) := X"24420001";
        ram_buffer(39206) := X"AE220000";
        ram_buffer(39207) := X"10000007";
        ram_buffer(39208) := X"00000000";
        ram_buffer(39209) := X"02202821";
        ram_buffer(39210) := X"8FC40340";
        ram_buffer(39211) := X"0C02E477";
        ram_buffer(39212) := X"00000000";
        ram_buffer(39213) := X"14400009";
        ram_buffer(39214) := X"00000000";
        ram_buffer(39215) := X"2652FFFF";
        ram_buffer(39216) := X"1640FF6B";
        ram_buffer(39217) := X"00000000";
        ram_buffer(39218) := X"10000005";
        ram_buffer(39219) := X"00000000";
        ram_buffer(39220) := X"00000000";
        ram_buffer(39221) := X"10000002";
        ram_buffer(39222) := X"00000000";
        ram_buffer(39223) := X"00000000";
        ram_buffer(39224) := X"32020100";
        ram_buffer(39225) := X"1040000F";
        ram_buffer(39226) := X"00000000";
        ram_buffer(39227) := X"27C201A8";
        ram_buffer(39228) := X"0053102B";
        ram_buffer(39229) := X"10400008";
        ram_buffer(39230) := X"00000000";
        ram_buffer(39231) := X"2673FFFF";
        ram_buffer(39232) := X"82620000";
        ram_buffer(39233) := X"02203021";
        ram_buffer(39234) := X"00402821";
        ram_buffer(39235) := X"8FC40340";
        ram_buffer(39236) := X"0C02E402";
        ram_buffer(39237) := X"00000000";
        ram_buffer(39238) := X"27C201A8";
        ram_buffer(39239) := X"12620319";
        ram_buffer(39240) := X"00000000";
        ram_buffer(39241) := X"32020010";
        ram_buffer(39242) := X"1440008B";
        ram_buffer(39243) := X"00000000";
        ram_buffer(39244) := X"A2600000";
        ram_buffer(39245) := X"27C301A8";
        ram_buffer(39246) := X"8FC20028";
        ram_buffer(39247) := X"8FC70020";
        ram_buffer(39248) := X"00003021";
        ram_buffer(39249) := X"00602821";
        ram_buffer(39250) := X"8FC40340";
        ram_buffer(39251) := X"0040F809";
        ram_buffer(39252) := X"00000000";
        ram_buffer(39253) := X"AFC20084";
        ram_buffer(39254) := X"32020020";
        ram_buffer(39255) := X"1040000E";
        ram_buffer(39256) := X"00000000";
        ram_buffer(39257) := X"8FC2034C";
        ram_buffer(39258) := X"00000000";
        ram_buffer(39259) := X"24430004";
        ram_buffer(39260) := X"AFC3034C";
        ram_buffer(39261) := X"8C420000";
        ram_buffer(39262) := X"00000000";
        ram_buffer(39263) := X"AFC20088";
        ram_buffer(39264) := X"8FC30084";
        ram_buffer(39265) := X"8FC20088";
        ram_buffer(39266) := X"00000000";
        ram_buffer(39267) := X"AC430000";
        ram_buffer(39268) := X"1000006D";
        ram_buffer(39269) := X"00000000";
        ram_buffer(39270) := X"32020008";
        ram_buffer(39271) := X"10400011";
        ram_buffer(39272) := X"00000000";
        ram_buffer(39273) := X"8FC2034C";
        ram_buffer(39274) := X"00000000";
        ram_buffer(39275) := X"24430004";
        ram_buffer(39276) := X"AFC3034C";
        ram_buffer(39277) := X"8C420000";
        ram_buffer(39278) := X"00000000";
        ram_buffer(39279) := X"AFC20068";
        ram_buffer(39280) := X"8FC20084";
        ram_buffer(39281) := X"00000000";
        ram_buffer(39282) := X"00021E00";
        ram_buffer(39283) := X"00031E03";
        ram_buffer(39284) := X"8FC20068";
        ram_buffer(39285) := X"00000000";
        ram_buffer(39286) := X"A0430000";
        ram_buffer(39287) := X"1000005A";
        ram_buffer(39288) := X"00000000";
        ram_buffer(39289) := X"32020004";
        ram_buffer(39290) := X"10400011";
        ram_buffer(39291) := X"00000000";
        ram_buffer(39292) := X"8FC2034C";
        ram_buffer(39293) := X"00000000";
        ram_buffer(39294) := X"24430004";
        ram_buffer(39295) := X"AFC3034C";
        ram_buffer(39296) := X"8C420000";
        ram_buffer(39297) := X"00000000";
        ram_buffer(39298) := X"AFC2006C";
        ram_buffer(39299) := X"8FC20084";
        ram_buffer(39300) := X"00000000";
        ram_buffer(39301) := X"00021C00";
        ram_buffer(39302) := X"00031C03";
        ram_buffer(39303) := X"8FC2006C";
        ram_buffer(39304) := X"00000000";
        ram_buffer(39305) := X"A4430000";
        ram_buffer(39306) := X"10000047";
        ram_buffer(39307) := X"00000000";
        ram_buffer(39308) := X"32020001";
        ram_buffer(39309) := X"1040000E";
        ram_buffer(39310) := X"00000000";
        ram_buffer(39311) := X"8FC2034C";
        ram_buffer(39312) := X"00000000";
        ram_buffer(39313) := X"24430004";
        ram_buffer(39314) := X"AFC3034C";
        ram_buffer(39315) := X"8C420000";
        ram_buffer(39316) := X"00000000";
        ram_buffer(39317) := X"AFC20070";
        ram_buffer(39318) := X"8FC30084";
        ram_buffer(39319) := X"8FC20070";
        ram_buffer(39320) := X"00000000";
        ram_buffer(39321) := X"AC430000";
        ram_buffer(39322) := X"10000037";
        ram_buffer(39323) := X"00000000";
        ram_buffer(39324) := X"32020002";
        ram_buffer(39325) := X"10400029";
        ram_buffer(39326) := X"00000000";
        ram_buffer(39327) := X"8FC30028";
        ram_buffer(39328) := X"3C02100B";
        ram_buffer(39329) := X"24426A64";
        ram_buffer(39330) := X"1462000C";
        ram_buffer(39331) := X"00000000";
        ram_buffer(39332) := X"27C201A8";
        ram_buffer(39333) := X"8FC70020";
        ram_buffer(39334) := X"00003021";
        ram_buffer(39335) := X"00402821";
        ram_buffer(39336) := X"8FC40340";
        ram_buffer(39337) := X"0C02DB85";
        ram_buffer(39338) := X"00000000";
        ram_buffer(39339) := X"AFC30044";
        ram_buffer(39340) := X"AFC20040";
        ram_buffer(39341) := X"1000000A";
        ram_buffer(39342) := X"00000000";
        ram_buffer(39343) := X"27C201A8";
        ram_buffer(39344) := X"8FC70020";
        ram_buffer(39345) := X"00003021";
        ram_buffer(39346) := X"00402821";
        ram_buffer(39347) := X"8FC40340";
        ram_buffer(39348) := X"0C02D961";
        ram_buffer(39349) := X"00000000";
        ram_buffer(39350) := X"AFC30044";
        ram_buffer(39351) := X"AFC20040";
        ram_buffer(39352) := X"8FC2034C";
        ram_buffer(39353) := X"00000000";
        ram_buffer(39354) := X"24430004";
        ram_buffer(39355) := X"AFC3034C";
        ram_buffer(39356) := X"8C420000";
        ram_buffer(39357) := X"00000000";
        ram_buffer(39358) := X"AFC20074";
        ram_buffer(39359) := X"8FC30044";
        ram_buffer(39360) := X"8FC20040";
        ram_buffer(39361) := X"8FC40074";
        ram_buffer(39362) := X"00000000";
        ram_buffer(39363) := X"AC830004";
        ram_buffer(39364) := X"AC820000";
        ram_buffer(39365) := X"1000000C";
        ram_buffer(39366) := X"00000000";
        ram_buffer(39367) := X"8FC2034C";
        ram_buffer(39368) := X"00000000";
        ram_buffer(39369) := X"24430004";
        ram_buffer(39370) := X"AFC3034C";
        ram_buffer(39371) := X"8C420000";
        ram_buffer(39372) := X"00000000";
        ram_buffer(39373) := X"AFC20078";
        ram_buffer(39374) := X"8FC30084";
        ram_buffer(39375) := X"8FC20078";
        ram_buffer(39376) := X"00000000";
        ram_buffer(39377) := X"AC430000";
        ram_buffer(39378) := X"8FC20018";
        ram_buffer(39379) := X"00000000";
        ram_buffer(39380) := X"24420001";
        ram_buffer(39381) := X"AFC20018";
        ram_buffer(39382) := X"02601821";
        ram_buffer(39383) := X"27C201A8";
        ram_buffer(39384) := X"00621823";
        ram_buffer(39385) := X"8FC20038";
        ram_buffer(39386) := X"00000000";
        ram_buffer(39387) := X"00621021";
        ram_buffer(39388) := X"8FC3001C";
        ram_buffer(39389) := X"00000000";
        ram_buffer(39390) := X"00621021";
        ram_buffer(39391) := X"AFC2001C";
        ram_buffer(39392) := X"1000024F";
        ram_buffer(39393) := X"00000000";
        ram_buffer(39394) := X"AFC00048";
        ram_buffer(39395) := X"AFC00054";
        ram_buffer(39396) := X"AFC00058";
        ram_buffer(39397) := X"A3C0005C";
        ram_buffer(39398) := X"A3C0005D";
        ram_buffer(39399) := X"8FC40340";
        ram_buffer(39400) := X"0C02BB25";
        ram_buffer(39401) := X"00000000";
        ram_buffer(39402) := X"8C420000";
        ram_buffer(39403) := X"00000000";
        ram_buffer(39404) := X"AFC2008C";
        ram_buffer(39405) := X"2642FFFF";
        ram_buffer(39406) := X"2C42015D";
        ram_buffer(39407) := X"14400004";
        ram_buffer(39408) := X"00000000";
        ram_buffer(39409) := X"2642FEA3";
        ram_buffer(39410) := X"AFC20058";
        ram_buffer(39411) := X"2412015D";
        ram_buffer(39412) := X"36100780";
        ram_buffer(39413) := X"AFC0004C";
        ram_buffer(39414) := X"AFC00050";
        ram_buffer(39415) := X"27D301A8";
        ram_buffer(39416) := X"1000010E";
        ram_buffer(39417) := X"00000000";
        ram_buffer(39418) := X"8E220000";
        ram_buffer(39419) := X"00000000";
        ram_buffer(39420) := X"90420000";
        ram_buffer(39421) := X"00000000";
        ram_buffer(39422) := X"0040A021";
        ram_buffer(39423) := X"2682FFD5";
        ram_buffer(39424) := X"2C43004F";
        ram_buffer(39425) := X"106000B4";
        ram_buffer(39426) := X"00000000";
        ram_buffer(39427) := X"00021880";
        ram_buffer(39428) := X"3C02100D";
        ram_buffer(39429) := X"2442A5A4";
        ram_buffer(39430) := X"00621021";
        ram_buffer(39431) := X"8C420000";
        ram_buffer(39432) := X"00000000";
        ram_buffer(39433) := X"00400008";
        ram_buffer(39434) := X"00000000";
        ram_buffer(39435) := X"32020100";
        ram_buffer(39436) := X"10400012";
        ram_buffer(39437) := X"00000000";
        ram_buffer(39438) := X"2402FF7F";
        ram_buffer(39439) := X"02028024";
        ram_buffer(39440) := X"8FC2004C";
        ram_buffer(39441) := X"00000000";
        ram_buffer(39442) := X"24420001";
        ram_buffer(39443) := X"AFC2004C";
        ram_buffer(39444) := X"8FC20058";
        ram_buffer(39445) := X"00000000";
        ram_buffer(39446) := X"104000D6";
        ram_buffer(39447) := X"00000000";
        ram_buffer(39448) := X"8FC20058";
        ram_buffer(39449) := X"00000000";
        ram_buffer(39450) := X"2442FFFF";
        ram_buffer(39451) := X"AFC20058";
        ram_buffer(39452) := X"26520001";
        ram_buffer(39453) := X"100000CF";
        ram_buffer(39454) := X"00000000";
        ram_buffer(39455) := X"83C3005C";
        ram_buffer(39456) := X"83C2005D";
        ram_buffer(39457) := X"00000000";
        ram_buffer(39458) := X"00621021";
        ram_buffer(39459) := X"144000A4";
        ram_buffer(39460) := X"00000000";
        ram_buffer(39461) := X"2402FE7F";
        ram_buffer(39462) := X"02028024";
        ram_buffer(39463) := X"100000BE";
        ram_buffer(39464) := X"00000000";
        ram_buffer(39465) := X"32020080";
        ram_buffer(39466) := X"104000A0";
        ram_buffer(39467) := X"00000000";
        ram_buffer(39468) := X"2402FF7F";
        ram_buffer(39469) := X"02028024";
        ram_buffer(39470) := X"100000B7";
        ram_buffer(39471) := X"00000000";
        ram_buffer(39472) := X"83C2005C";
        ram_buffer(39473) := X"00000000";
        ram_buffer(39474) := X"1440000F";
        ram_buffer(39475) := X"00000000";
        ram_buffer(39476) := X"8FC2004C";
        ram_buffer(39477) := X"00000000";
        ram_buffer(39478) := X"1440000B";
        ram_buffer(39479) := X"00000000";
        ram_buffer(39480) := X"32030700";
        ram_buffer(39481) := X"24020700";
        ram_buffer(39482) := X"14620007";
        ram_buffer(39483) := X"00000000";
        ram_buffer(39484) := X"2402F87F";
        ram_buffer(39485) := X"02028024";
        ram_buffer(39486) := X"24020001";
        ram_buffer(39487) := X"A3C2005C";
        ram_buffer(39488) := X"100000A5";
        ram_buffer(39489) := X"00000000";
        ram_buffer(39490) := X"83C3005C";
        ram_buffer(39491) := X"24020002";
        ram_buffer(39492) := X"14620005";
        ram_buffer(39493) := X"00000000";
        ram_buffer(39494) := X"24020003";
        ram_buffer(39495) := X"A3C2005C";
        ram_buffer(39496) := X"1000009D";
        ram_buffer(39497) := X"00000000";
        ram_buffer(39498) := X"83C3005D";
        ram_buffer(39499) := X"24020001";
        ram_buffer(39500) := X"10620005";
        ram_buffer(39501) := X"00000000";
        ram_buffer(39502) := X"83C3005D";
        ram_buffer(39503) := X"24020004";
        ram_buffer(39504) := X"1462007D";
        ram_buffer(39505) := X"00000000";
        ram_buffer(39506) := X"83C2005D";
        ram_buffer(39507) := X"00000000";
        ram_buffer(39508) := X"304200FF";
        ram_buffer(39509) := X"24420001";
        ram_buffer(39510) := X"304200FF";
        ram_buffer(39511) := X"A3C2005D";
        ram_buffer(39512) := X"1000008D";
        ram_buffer(39513) := X"00000000";
        ram_buffer(39514) := X"83C3005C";
        ram_buffer(39515) := X"24020001";
        ram_buffer(39516) := X"14620074";
        ram_buffer(39517) := X"00000000";
        ram_buffer(39518) := X"24020002";
        ram_buffer(39519) := X"A3C2005C";
        ram_buffer(39520) := X"10000085";
        ram_buffer(39521) := X"00000000";
        ram_buffer(39522) := X"83C2005D";
        ram_buffer(39523) := X"00000000";
        ram_buffer(39524) := X"1440000F";
        ram_buffer(39525) := X"00000000";
        ram_buffer(39526) := X"8FC2004C";
        ram_buffer(39527) := X"00000000";
        ram_buffer(39528) := X"1440000B";
        ram_buffer(39529) := X"00000000";
        ram_buffer(39530) := X"32030700";
        ram_buffer(39531) := X"24020700";
        ram_buffer(39532) := X"14620007";
        ram_buffer(39533) := X"00000000";
        ram_buffer(39534) := X"2402F87F";
        ram_buffer(39535) := X"02028024";
        ram_buffer(39536) := X"24020001";
        ram_buffer(39537) := X"A3C2005D";
        ram_buffer(39538) := X"10000073";
        ram_buffer(39539) := X"00000000";
        ram_buffer(39540) := X"83C3005D";
        ram_buffer(39541) := X"24020003";
        ram_buffer(39542) := X"10620005";
        ram_buffer(39543) := X"00000000";
        ram_buffer(39544) := X"83C3005D";
        ram_buffer(39545) := X"24020005";
        ram_buffer(39546) := X"14620059";
        ram_buffer(39547) := X"00000000";
        ram_buffer(39548) := X"83C2005D";
        ram_buffer(39549) := X"00000000";
        ram_buffer(39550) := X"304200FF";
        ram_buffer(39551) := X"24420001";
        ram_buffer(39552) := X"304200FF";
        ram_buffer(39553) := X"A3C2005D";
        ram_buffer(39554) := X"10000063";
        ram_buffer(39555) := X"00000000";
        ram_buffer(39556) := X"83C3005D";
        ram_buffer(39557) := X"24020002";
        ram_buffer(39558) := X"14620050";
        ram_buffer(39559) := X"00000000";
        ram_buffer(39560) := X"24020003";
        ram_buffer(39561) := X"A3C2005D";
        ram_buffer(39562) := X"1000005B";
        ram_buffer(39563) := X"00000000";
        ram_buffer(39564) := X"83C3005D";
        ram_buffer(39565) := X"24020006";
        ram_buffer(39566) := X"1462004B";
        ram_buffer(39567) := X"00000000";
        ram_buffer(39568) := X"24020007";
        ram_buffer(39569) := X"A3C2005D";
        ram_buffer(39570) := X"10000053";
        ram_buffer(39571) := X"00000000";
        ram_buffer(39572) := X"83C3005D";
        ram_buffer(39573) := X"24020007";
        ram_buffer(39574) := X"14620046";
        ram_buffer(39575) := X"00000000";
        ram_buffer(39576) := X"24020008";
        ram_buffer(39577) := X"A3C2005D";
        ram_buffer(39578) := X"1000004B";
        ram_buffer(39579) := X"00000000";
        ram_buffer(39580) := X"32030500";
        ram_buffer(39581) := X"24020400";
        ram_buffer(39582) := X"10620008";
        ram_buffer(39583) := X"00000000";
        ram_buffer(39584) := X"32020400";
        ram_buffer(39585) := X"1040003E";
        ram_buffer(39586) := X"00000000";
        ram_buffer(39587) := X"8FC2004C";
        ram_buffer(39588) := X"00000000";
        ram_buffer(39589) := X"1040003A";
        ram_buffer(39590) := X"00000000";
        ram_buffer(39591) := X"32020200";
        ram_buffer(39592) := X"14400007";
        ram_buffer(39593) := X"00000000";
        ram_buffer(39594) := X"8FC3004C";
        ram_buffer(39595) := X"8FC20048";
        ram_buffer(39596) := X"00000000";
        ram_buffer(39597) := X"00621023";
        ram_buffer(39598) := X"AFC20050";
        ram_buffer(39599) := X"AFD30054";
        ram_buffer(39600) := X"2402F87F";
        ram_buffer(39601) := X"02021024";
        ram_buffer(39602) := X"34500180";
        ram_buffer(39603) := X"AFC0004C";
        ram_buffer(39604) := X"10000031";
        ram_buffer(39605) := X"00000000";
        ram_buffer(39606) := X"328200FF";
        ram_buffer(39607) := X"8FC3008C";
        ram_buffer(39608) := X"00000000";
        ram_buffer(39609) := X"80630000";
        ram_buffer(39610) := X"00000000";
        ram_buffer(39611) := X"306300FF";
        ram_buffer(39612) := X"14430026";
        ram_buffer(39613) := X"00000000";
        ram_buffer(39614) := X"32020200";
        ram_buffer(39615) := X"10400023";
        ram_buffer(39616) := X"00000000";
        ram_buffer(39617) := X"2402FD7F";
        ram_buffer(39618) := X"02028024";
        ram_buffer(39619) := X"8FC2004C";
        ram_buffer(39620) := X"00000000";
        ram_buffer(39621) := X"AFC20048";
        ram_buffer(39622) := X"1000001F";
        ram_buffer(39623) := X"00000000";
        ram_buffer(39624) := X"00000000";
        ram_buffer(39625) := X"10000042";
        ram_buffer(39626) := X"00000000";
        ram_buffer(39627) := X"00000000";
        ram_buffer(39628) := X"1000003F";
        ram_buffer(39629) := X"00000000";
        ram_buffer(39630) := X"00000000";
        ram_buffer(39631) := X"1000003C";
        ram_buffer(39632) := X"00000000";
        ram_buffer(39633) := X"00000000";
        ram_buffer(39634) := X"10000039";
        ram_buffer(39635) := X"00000000";
        ram_buffer(39636) := X"00000000";
        ram_buffer(39637) := X"10000036";
        ram_buffer(39638) := X"00000000";
        ram_buffer(39639) := X"00000000";
        ram_buffer(39640) := X"10000033";
        ram_buffer(39641) := X"00000000";
        ram_buffer(39642) := X"00000000";
        ram_buffer(39643) := X"10000030";
        ram_buffer(39644) := X"00000000";
        ram_buffer(39645) := X"00000000";
        ram_buffer(39646) := X"1000002D";
        ram_buffer(39647) := X"00000000";
        ram_buffer(39648) := X"00000000";
        ram_buffer(39649) := X"1000002A";
        ram_buffer(39650) := X"00000000";
        ram_buffer(39651) := X"00000000";
        ram_buffer(39652) := X"10000027";
        ram_buffer(39653) := X"00000000";
        ram_buffer(39654) := X"02601021";
        ram_buffer(39655) := X"24530001";
        ram_buffer(39656) := X"00141E00";
        ram_buffer(39657) := X"00031E03";
        ram_buffer(39658) := X"A0430000";
        ram_buffer(39659) := X"10000002";
        ram_buffer(39660) := X"00000000";
        ram_buffer(39661) := X"00000000";
        ram_buffer(39662) := X"2652FFFF";
        ram_buffer(39663) := X"8FC2001C";
        ram_buffer(39664) := X"00000000";
        ram_buffer(39665) := X"24420001";
        ram_buffer(39666) := X"AFC2001C";
        ram_buffer(39667) := X"8E220004";
        ram_buffer(39668) := X"00000000";
        ram_buffer(39669) := X"2442FFFF";
        ram_buffer(39670) := X"AE220004";
        ram_buffer(39671) := X"8E220004";
        ram_buffer(39672) := X"00000000";
        ram_buffer(39673) := X"18400007";
        ram_buffer(39674) := X"00000000";
        ram_buffer(39675) := X"8E220000";
        ram_buffer(39676) := X"00000000";
        ram_buffer(39677) := X"24420001";
        ram_buffer(39678) := X"AE220000";
        ram_buffer(39679) := X"10000007";
        ram_buffer(39680) := X"00000000";
        ram_buffer(39681) := X"02202821";
        ram_buffer(39682) := X"8FC40340";
        ram_buffer(39683) := X"0C02E477";
        ram_buffer(39684) := X"00000000";
        ram_buffer(39685) := X"14400005";
        ram_buffer(39686) := X"00000000";
        ram_buffer(39687) := X"1640FEF2";
        ram_buffer(39688) := X"00000000";
        ram_buffer(39689) := X"10000002";
        ram_buffer(39690) := X"00000000";
        ram_buffer(39691) := X"00000000";
        ram_buffer(39692) := X"8FC2004C";
        ram_buffer(39693) := X"00000000";
        ram_buffer(39694) := X"10400003";
        ram_buffer(39695) := X"00000000";
        ram_buffer(39696) := X"2402FEFF";
        ram_buffer(39697) := X"02028024";
        ram_buffer(39698) := X"83C2005C";
        ram_buffer(39699) := X"00000000";
        ram_buffer(39700) := X"2442FFFF";
        ram_buffer(39701) := X"2C420002";
        ram_buffer(39702) := X"10400014";
        ram_buffer(39703) := X"00000000";
        ram_buffer(39704) := X"1000000C";
        ram_buffer(39705) := X"00000000";
        ram_buffer(39706) := X"2673FFFF";
        ram_buffer(39707) := X"82620000";
        ram_buffer(39708) := X"02203021";
        ram_buffer(39709) := X"00402821";
        ram_buffer(39710) := X"8FC40340";
        ram_buffer(39711) := X"0C02E402";
        ram_buffer(39712) := X"00000000";
        ram_buffer(39713) := X"8FC2001C";
        ram_buffer(39714) := X"00000000";
        ram_buffer(39715) := X"2442FFFF";
        ram_buffer(39716) := X"AFC2001C";
        ram_buffer(39717) := X"27C201A8";
        ram_buffer(39718) := X"0053102B";
        ram_buffer(39719) := X"1440FFF2";
        ram_buffer(39720) := X"00000000";
        ram_buffer(39721) := X"10000138";
        ram_buffer(39722) := X"00000000";
        ram_buffer(39723) := X"83C2005D";
        ram_buffer(39724) := X"00000000";
        ram_buffer(39725) := X"2442FFFF";
        ram_buffer(39726) := X"2C420007";
        ram_buffer(39727) := X"1040002F";
        ram_buffer(39728) := X"00000000";
        ram_buffer(39729) := X"83C2005D";
        ram_buffer(39730) := X"00000000";
        ram_buffer(39731) := X"28420003";
        ram_buffer(39732) := X"14400024";
        ram_buffer(39733) := X"00000000";
        ram_buffer(39734) := X"1000000C";
        ram_buffer(39735) := X"00000000";
        ram_buffer(39736) := X"2673FFFF";
        ram_buffer(39737) := X"82620000";
        ram_buffer(39738) := X"02203021";
        ram_buffer(39739) := X"00402821";
        ram_buffer(39740) := X"8FC40340";
        ram_buffer(39741) := X"0C02E402";
        ram_buffer(39742) := X"00000000";
        ram_buffer(39743) := X"8FC2001C";
        ram_buffer(39744) := X"00000000";
        ram_buffer(39745) := X"2442FFFF";
        ram_buffer(39746) := X"AFC2001C";
        ram_buffer(39747) := X"83C2005D";
        ram_buffer(39748) := X"00000000";
        ram_buffer(39749) := X"304300FF";
        ram_buffer(39750) := X"2463FFFF";
        ram_buffer(39751) := X"306300FF";
        ram_buffer(39752) := X"A3C3005D";
        ram_buffer(39753) := X"28420004";
        ram_buffer(39754) := X"1040FFED";
        ram_buffer(39755) := X"00000000";
        ram_buffer(39756) := X"10000012";
        ram_buffer(39757) := X"00000000";
        ram_buffer(39758) := X"2673FFFF";
        ram_buffer(39759) := X"82620000";
        ram_buffer(39760) := X"02203021";
        ram_buffer(39761) := X"00402821";
        ram_buffer(39762) := X"8FC40340";
        ram_buffer(39763) := X"0C02E402";
        ram_buffer(39764) := X"00000000";
        ram_buffer(39765) := X"8FC2001C";
        ram_buffer(39766) := X"00000000";
        ram_buffer(39767) := X"2442FFFF";
        ram_buffer(39768) := X"AFC2001C";
        ram_buffer(39769) := X"27C201A8";
        ram_buffer(39770) := X"0053102B";
        ram_buffer(39771) := X"1440FFF2";
        ram_buffer(39772) := X"00000000";
        ram_buffer(39773) := X"10000104";
        ram_buffer(39774) := X"00000000";
        ram_buffer(39775) := X"32020100";
        ram_buffer(39776) := X"10400037";
        ram_buffer(39777) := X"00000000";
        ram_buffer(39778) := X"32020400";
        ram_buffer(39779) := X"10400014";
        ram_buffer(39780) := X"00000000";
        ram_buffer(39781) := X"1000000C";
        ram_buffer(39782) := X"00000000";
        ram_buffer(39783) := X"2673FFFF";
        ram_buffer(39784) := X"82620000";
        ram_buffer(39785) := X"02203021";
        ram_buffer(39786) := X"00402821";
        ram_buffer(39787) := X"8FC40340";
        ram_buffer(39788) := X"0C02E402";
        ram_buffer(39789) := X"00000000";
        ram_buffer(39790) := X"8FC2001C";
        ram_buffer(39791) := X"00000000";
        ram_buffer(39792) := X"2442FFFF";
        ram_buffer(39793) := X"AFC2001C";
        ram_buffer(39794) := X"27C201A8";
        ram_buffer(39795) := X"0053102B";
        ram_buffer(39796) := X"1440FFF2";
        ram_buffer(39797) := X"00000000";
        ram_buffer(39798) := X"100000EB";
        ram_buffer(39799) := X"00000000";
        ram_buffer(39800) := X"2673FFFF";
        ram_buffer(39801) := X"82620000";
        ram_buffer(39802) := X"00000000";
        ram_buffer(39803) := X"0040A021";
        ram_buffer(39804) := X"8FC2001C";
        ram_buffer(39805) := X"00000000";
        ram_buffer(39806) := X"2442FFFF";
        ram_buffer(39807) := X"AFC2001C";
        ram_buffer(39808) := X"24020065";
        ram_buffer(39809) := X"12820011";
        ram_buffer(39810) := X"00000000";
        ram_buffer(39811) := X"24020045";
        ram_buffer(39812) := X"1282000E";
        ram_buffer(39813) := X"00000000";
        ram_buffer(39814) := X"02203021";
        ram_buffer(39815) := X"02802821";
        ram_buffer(39816) := X"8FC40340";
        ram_buffer(39817) := X"0C02E402";
        ram_buffer(39818) := X"00000000";
        ram_buffer(39819) := X"2673FFFF";
        ram_buffer(39820) := X"82620000";
        ram_buffer(39821) := X"00000000";
        ram_buffer(39822) := X"0040A021";
        ram_buffer(39823) := X"8FC2001C";
        ram_buffer(39824) := X"00000000";
        ram_buffer(39825) := X"2442FFFF";
        ram_buffer(39826) := X"AFC2001C";
        ram_buffer(39827) := X"02203021";
        ram_buffer(39828) := X"02802821";
        ram_buffer(39829) := X"8FC40340";
        ram_buffer(39830) := X"0C02E402";
        ram_buffer(39831) := X"00000000";
        ram_buffer(39832) := X"32020010";
        ram_buffer(39833) := X"14400095";
        ram_buffer(39834) := X"00000000";
        ram_buffer(39835) := X"AFC00094";
        ram_buffer(39836) := X"AFC00090";
        ram_buffer(39837) := X"AFC00060";
        ram_buffer(39838) := X"A2600000";
        ram_buffer(39839) := X"32030600";
        ram_buffer(39840) := X"24020400";
        ram_buffer(39841) := X"1462000D";
        ram_buffer(39842) := X"00000000";
        ram_buffer(39843) := X"8FC3004C";
        ram_buffer(39844) := X"8FC20048";
        ram_buffer(39845) := X"00000000";
        ram_buffer(39846) := X"00621023";
        ram_buffer(39847) := X"AFC20050";
        ram_buffer(39848) := X"8FC20050";
        ram_buffer(39849) := X"00000000";
        ram_buffer(39850) := X"00021023";
        ram_buffer(39851) := X"AFC20060";
        ram_buffer(39852) := X"AFD30054";
        ram_buffer(39853) := X"10000013";
        ram_buffer(39854) := X"00000000";
        ram_buffer(39855) := X"8FC20050";
        ram_buffer(39856) := X"00000000";
        ram_buffer(39857) := X"1040000F";
        ram_buffer(39858) := X"00000000";
        ram_buffer(39859) := X"8FC20054";
        ram_buffer(39860) := X"00000000";
        ram_buffer(39861) := X"24420001";
        ram_buffer(39862) := X"2407000A";
        ram_buffer(39863) := X"00003021";
        ram_buffer(39864) := X"00402821";
        ram_buffer(39865) := X"8FC40340";
        ram_buffer(39866) := X"0C02D866";
        ram_buffer(39867) := X"00000000";
        ram_buffer(39868) := X"00401821";
        ram_buffer(39869) := X"8FC20050";
        ram_buffer(39870) := X"00000000";
        ram_buffer(39871) := X"00621023";
        ram_buffer(39872) := X"AFC20060";
        ram_buffer(39873) := X"8FC20050";
        ram_buffer(39874) := X"00000000";
        ram_buffer(39875) := X"10400011";
        ram_buffer(39876) := X"00000000";
        ram_buffer(39877) := X"27C201A8";
        ram_buffer(39878) := X"24420153";
        ram_buffer(39879) := X"8FC30054";
        ram_buffer(39880) := X"00000000";
        ram_buffer(39881) := X"0062102B";
        ram_buffer(39882) := X"14400004";
        ram_buffer(39883) := X"00000000";
        ram_buffer(39884) := X"27C201A8";
        ram_buffer(39885) := X"24420152";
        ram_buffer(39886) := X"AFC20054";
        ram_buffer(39887) := X"8FC60060";
        ram_buffer(39888) := X"3C02100D";
        ram_buffer(39889) := X"2445A264";
        ram_buffer(39890) := X"8FC40054";
        ram_buffer(39891) := X"0C0283DB";
        ram_buffer(39892) := X"00000000";
        ram_buffer(39893) := X"27C201A8";
        ram_buffer(39894) := X"00003021";
        ram_buffer(39895) := X"00402821";
        ram_buffer(39896) := X"8FC40340";
        ram_buffer(39897) := X"0C02CF1C";
        ram_buffer(39898) := X"00000000";
        ram_buffer(39899) := X"AFC30094";
        ram_buffer(39900) := X"AFC20090";
        ram_buffer(39901) := X"32020001";
        ram_buffer(39902) := X"1040000F";
        ram_buffer(39903) := X"00000000";
        ram_buffer(39904) := X"8FC2034C";
        ram_buffer(39905) := X"00000000";
        ram_buffer(39906) := X"24430004";
        ram_buffer(39907) := X"AFC3034C";
        ram_buffer(39908) := X"8C420000";
        ram_buffer(39909) := X"00000000";
        ram_buffer(39910) := X"AFC20098";
        ram_buffer(39911) := X"8FC40098";
        ram_buffer(39912) := X"8FC30094";
        ram_buffer(39913) := X"8FC20090";
        ram_buffer(39914) := X"AC830004";
        ram_buffer(39915) := X"AC820000";
        ram_buffer(39916) := X"10000030";
        ram_buffer(39917) := X"00000000";
        ram_buffer(39918) := X"32020002";
        ram_buffer(39919) := X"1040000F";
        ram_buffer(39920) := X"00000000";
        ram_buffer(39921) := X"8FC2034C";
        ram_buffer(39922) := X"00000000";
        ram_buffer(39923) := X"24430004";
        ram_buffer(39924) := X"AFC3034C";
        ram_buffer(39925) := X"8C420000";
        ram_buffer(39926) := X"00000000";
        ram_buffer(39927) := X"AFC2009C";
        ram_buffer(39928) := X"8FC4009C";
        ram_buffer(39929) := X"8FC30094";
        ram_buffer(39930) := X"8FC20090";
        ram_buffer(39931) := X"AC830004";
        ram_buffer(39932) := X"AC820000";
        ram_buffer(39933) := X"1000001F";
        ram_buffer(39934) := X"00000000";
        ram_buffer(39935) := X"8FC2034C";
        ram_buffer(39936) := X"00000000";
        ram_buffer(39937) := X"24430004";
        ram_buffer(39938) := X"AFC3034C";
        ram_buffer(39939) := X"8C420000";
        ram_buffer(39940) := X"00000000";
        ram_buffer(39941) := X"AFC200A0";
        ram_buffer(39942) := X"8FC50094";
        ram_buffer(39943) := X"8FC40090";
        ram_buffer(39944) := X"0C02CAED";
        ram_buffer(39945) := X"00000000";
        ram_buffer(39946) := X"1440000A";
        ram_buffer(39947) := X"00000000";
        ram_buffer(39948) := X"00002021";
        ram_buffer(39949) := X"0C02CC22";
        ram_buffer(39950) := X"00000000";
        ram_buffer(39951) := X"00401821";
        ram_buffer(39952) := X"8FC200A0";
        ram_buffer(39953) := X"00000000";
        ram_buffer(39954) := X"AC430000";
        ram_buffer(39955) := X"10000009";
        ram_buffer(39956) := X"00000000";
        ram_buffer(39957) := X"8FC50094";
        ram_buffer(39958) := X"8FC40090";
        ram_buffer(39959) := X"0C031C96";
        ram_buffer(39960) := X"00000000";
        ram_buffer(39961) := X"00401821";
        ram_buffer(39962) := X"8FC200A0";
        ram_buffer(39963) := X"00000000";
        ram_buffer(39964) := X"AC430000";
        ram_buffer(39965) := X"8FC20018";
        ram_buffer(39966) := X"00000000";
        ram_buffer(39967) := X"24420001";
        ram_buffer(39968) := X"AFC20018";
        ram_buffer(39969) := X"1000000D";
        ram_buffer(39970) := X"00000000";
        ram_buffer(39971) := X"00000000";
        ram_buffer(39972) := X"1000F858";
        ram_buffer(39973) := X"00000000";
        ram_buffer(39974) := X"00000000";
        ram_buffer(39975) := X"1000F855";
        ram_buffer(39976) := X"00000000";
        ram_buffer(39977) := X"00000000";
        ram_buffer(39978) := X"1000F852";
        ram_buffer(39979) := X"00000000";
        ram_buffer(39980) := X"00000000";
        ram_buffer(39981) := X"1000F84F";
        ram_buffer(39982) := X"00000000";
        ram_buffer(39983) := X"00000000";
        ram_buffer(39984) := X"1000F84C";
        ram_buffer(39985) := X"00000000";
        ram_buffer(39986) := X"00000000";
        ram_buffer(39987) := X"10000014";
        ram_buffer(39988) := X"00000000";
        ram_buffer(39989) := X"00000000";
        ram_buffer(39990) := X"10000011";
        ram_buffer(39991) := X"00000000";
        ram_buffer(39992) := X"00000000";
        ram_buffer(39993) := X"1000000E";
        ram_buffer(39994) := X"00000000";
        ram_buffer(39995) := X"00000000";
        ram_buffer(39996) := X"1000000B";
        ram_buffer(39997) := X"00000000";
        ram_buffer(39998) := X"00000000";
        ram_buffer(39999) := X"10000008";
        ram_buffer(40000) := X"00000000";
        ram_buffer(40001) := X"00000000";
        ram_buffer(40002) := X"10000005";
        ram_buffer(40003) := X"00000000";
        ram_buffer(40004) := X"00000000";
        ram_buffer(40005) := X"10000002";
        ram_buffer(40006) := X"00000000";
        ram_buffer(40007) := X"00000000";
        ram_buffer(40008) := X"8FC20018";
        ram_buffer(40009) := X"00000000";
        ram_buffer(40010) := X"1040000A";
        ram_buffer(40011) := X"00000000";
        ram_buffer(40012) := X"8622000C";
        ram_buffer(40013) := X"00000000";
        ram_buffer(40014) := X"3042FFFF";
        ram_buffer(40015) := X"30420040";
        ram_buffer(40016) := X"14400004";
        ram_buffer(40017) := X"00000000";
        ram_buffer(40018) := X"8FC20018";
        ram_buffer(40019) := X"1000000F";
        ram_buffer(40020) := X"00000000";
        ram_buffer(40021) := X"2402FFFF";
        ram_buffer(40022) := X"1000000C";
        ram_buffer(40023) := X"00000000";
        ram_buffer(40024) := X"00000000";
        ram_buffer(40025) := X"10000008";
        ram_buffer(40026) := X"00000000";
        ram_buffer(40027) := X"00000000";
        ram_buffer(40028) := X"10000005";
        ram_buffer(40029) := X"00000000";
        ram_buffer(40030) := X"00000000";
        ram_buffer(40031) := X"10000002";
        ram_buffer(40032) := X"00000000";
        ram_buffer(40033) := X"00000000";
        ram_buffer(40034) := X"8FC20018";
        ram_buffer(40035) := X"03C0E821";
        ram_buffer(40036) := X"8FBF033C";
        ram_buffer(40037) := X"8FBE0338";
        ram_buffer(40038) := X"8FB70334";
        ram_buffer(40039) := X"8FB60330";
        ram_buffer(40040) := X"8FB5032C";
        ram_buffer(40041) := X"8FB40328";
        ram_buffer(40042) := X"8FB30324";
        ram_buffer(40043) := X"8FB20320";
        ram_buffer(40044) := X"8FB1031C";
        ram_buffer(40045) := X"8FB00318";
        ram_buffer(40046) := X"27BD0340";
        ram_buffer(40047) := X"03E00008";
        ram_buffer(40048) := X"00000000";
        ram_buffer(40049) := X"27BDFFD8";
        ram_buffer(40050) := X"AFBF0024";
        ram_buffer(40051) := X"AFBE0020";
        ram_buffer(40052) := X"AFB2001C";
        ram_buffer(40053) := X"AFB10018";
        ram_buffer(40054) := X"AFB00014";
        ram_buffer(40055) := X"03A0F021";
        ram_buffer(40056) := X"AFC40028";
        ram_buffer(40057) := X"00A08021";
        ram_buffer(40058) := X"8E030030";
        ram_buffer(40059) := X"26020040";
        ram_buffer(40060) := X"1462001F";
        ram_buffer(40061) := X"00000000";
        ram_buffer(40062) := X"24050400";
        ram_buffer(40063) := X"8FC40028";
        ram_buffer(40064) := X"0C027B8F";
        ram_buffer(40065) := X"00000000";
        ram_buffer(40066) := X"00408821";
        ram_buffer(40067) := X"16200004";
        ram_buffer(40068) := X"00000000";
        ram_buffer(40069) := X"2402FFFF";
        ram_buffer(40070) := X"10000032";
        ram_buffer(40071) := X"00000000";
        ram_buffer(40072) := X"AE110030";
        ram_buffer(40073) := X"24020400";
        ram_buffer(40074) := X"AE020034";
        ram_buffer(40075) := X"263103FD";
        ram_buffer(40076) := X"24120003";
        ram_buffer(40077) := X"10000007";
        ram_buffer(40078) := X"00000000";
        ram_buffer(40079) := X"02401021";
        ram_buffer(40080) := X"02221021";
        ram_buffer(40081) := X"02121821";
        ram_buffer(40082) := X"90630040";
        ram_buffer(40083) := X"00000000";
        ram_buffer(40084) := X"A0430000";
        ram_buffer(40085) := X"2652FFFF";
        ram_buffer(40086) := X"0641FFF8";
        ram_buffer(40087) := X"00000000";
        ram_buffer(40088) := X"AE110000";
        ram_buffer(40089) := X"00001021";
        ram_buffer(40090) := X"1000001E";
        ram_buffer(40091) := X"00000000";
        ram_buffer(40092) := X"8E120034";
        ram_buffer(40093) := X"8E020030";
        ram_buffer(40094) := X"00121840";
        ram_buffer(40095) := X"00603021";
        ram_buffer(40096) := X"00402821";
        ram_buffer(40097) := X"8FC40028";
        ram_buffer(40098) := X"0C02C6A7";
        ram_buffer(40099) := X"00000000";
        ram_buffer(40100) := X"00408821";
        ram_buffer(40101) := X"16200004";
        ram_buffer(40102) := X"00000000";
        ram_buffer(40103) := X"2402FFFF";
        ram_buffer(40104) := X"10000010";
        ram_buffer(40105) := X"00000000";
        ram_buffer(40106) := X"02401021";
        ram_buffer(40107) := X"02221021";
        ram_buffer(40108) := X"02401821";
        ram_buffer(40109) := X"00603021";
        ram_buffer(40110) := X"02202821";
        ram_buffer(40111) := X"00402021";
        ram_buffer(40112) := X"0C027F93";
        ram_buffer(40113) := X"00000000";
        ram_buffer(40114) := X"02401021";
        ram_buffer(40115) := X"02221021";
        ram_buffer(40116) := X"AE020000";
        ram_buffer(40117) := X"AE110030";
        ram_buffer(40118) := X"00121040";
        ram_buffer(40119) := X"AE020034";
        ram_buffer(40120) := X"00001021";
        ram_buffer(40121) := X"03C0E821";
        ram_buffer(40122) := X"8FBF0024";
        ram_buffer(40123) := X"8FBE0020";
        ram_buffer(40124) := X"8FB2001C";
        ram_buffer(40125) := X"8FB10018";
        ram_buffer(40126) := X"8FB00014";
        ram_buffer(40127) := X"27BD0028";
        ram_buffer(40128) := X"03E00008";
        ram_buffer(40129) := X"00000000";
        ram_buffer(40130) := X"27BDFFD8";
        ram_buffer(40131) := X"AFBF0024";
        ram_buffer(40132) := X"AFBE0020";
        ram_buffer(40133) := X"AFB0001C";
        ram_buffer(40134) := X"03A0F021";
        ram_buffer(40135) := X"AFC40028";
        ram_buffer(40136) := X"AFC5002C";
        ram_buffer(40137) := X"00C08021";
        ram_buffer(40138) := X"8FC3002C";
        ram_buffer(40139) := X"2402FFFF";
        ram_buffer(40140) := X"14620004";
        ram_buffer(40141) := X"00000000";
        ram_buffer(40142) := X"2402FFFF";
        ram_buffer(40143) := X"100000AC";
        ram_buffer(40144) := X"00000000";
        ram_buffer(40145) := X"8FC20028";
        ram_buffer(40146) := X"00000000";
        ram_buffer(40147) := X"AFC20010";
        ram_buffer(40148) := X"8FC20010";
        ram_buffer(40149) := X"00000000";
        ram_buffer(40150) := X"1040000A";
        ram_buffer(40151) := X"00000000";
        ram_buffer(40152) := X"8FC20010";
        ram_buffer(40153) := X"00000000";
        ram_buffer(40154) := X"8C420038";
        ram_buffer(40155) := X"00000000";
        ram_buffer(40156) := X"14400004";
        ram_buffer(40157) := X"00000000";
        ram_buffer(40158) := X"8FC40010";
        ram_buffer(40159) := X"0C027069";
        ram_buffer(40160) := X"00000000";
        ram_buffer(40161) := X"8602000C";
        ram_buffer(40162) := X"00000000";
        ram_buffer(40163) := X"3042FFFF";
        ram_buffer(40164) := X"30422000";
        ram_buffer(40165) := X"1440000B";
        ram_buffer(40166) := X"00000000";
        ram_buffer(40167) := X"8602000C";
        ram_buffer(40168) := X"00000000";
        ram_buffer(40169) := X"34422000";
        ram_buffer(40170) := X"00021400";
        ram_buffer(40171) := X"00021403";
        ram_buffer(40172) := X"A602000C";
        ram_buffer(40173) := X"8E030064";
        ram_buffer(40174) := X"2402DFFF";
        ram_buffer(40175) := X"00621024";
        ram_buffer(40176) := X"AE020064";
        ram_buffer(40177) := X"8603000C";
        ram_buffer(40178) := X"2402FFDF";
        ram_buffer(40179) := X"00621024";
        ram_buffer(40180) := X"00021400";
        ram_buffer(40181) := X"00021403";
        ram_buffer(40182) := X"A602000C";
        ram_buffer(40183) := X"8602000C";
        ram_buffer(40184) := X"00000000";
        ram_buffer(40185) := X"3042FFFF";
        ram_buffer(40186) := X"30420004";
        ram_buffer(40187) := X"14400027";
        ram_buffer(40188) := X"00000000";
        ram_buffer(40189) := X"8602000C";
        ram_buffer(40190) := X"00000000";
        ram_buffer(40191) := X"3042FFFF";
        ram_buffer(40192) := X"30420010";
        ram_buffer(40193) := X"14400004";
        ram_buffer(40194) := X"00000000";
        ram_buffer(40195) := X"2402FFFF";
        ram_buffer(40196) := X"10000077";
        ram_buffer(40197) := X"00000000";
        ram_buffer(40198) := X"8602000C";
        ram_buffer(40199) := X"00000000";
        ram_buffer(40200) := X"3042FFFF";
        ram_buffer(40201) := X"30420008";
        ram_buffer(40202) := X"10400012";
        ram_buffer(40203) := X"00000000";
        ram_buffer(40204) := X"02002821";
        ram_buffer(40205) := X"8FC40028";
        ram_buffer(40206) := X"0C026EE1";
        ram_buffer(40207) := X"00000000";
        ram_buffer(40208) := X"10400004";
        ram_buffer(40209) := X"00000000";
        ram_buffer(40210) := X"2402FFFF";
        ram_buffer(40211) := X"10000068";
        ram_buffer(40212) := X"00000000";
        ram_buffer(40213) := X"8603000C";
        ram_buffer(40214) := X"2402FFF7";
        ram_buffer(40215) := X"00621024";
        ram_buffer(40216) := X"00021400";
        ram_buffer(40217) := X"00021403";
        ram_buffer(40218) := X"A602000C";
        ram_buffer(40219) := X"AE000008";
        ram_buffer(40220) := X"AE000018";
        ram_buffer(40221) := X"8602000C";
        ram_buffer(40222) := X"00000000";
        ram_buffer(40223) := X"34420004";
        ram_buffer(40224) := X"00021400";
        ram_buffer(40225) := X"00021403";
        ram_buffer(40226) := X"A602000C";
        ram_buffer(40227) := X"8FC2002C";
        ram_buffer(40228) := X"00000000";
        ram_buffer(40229) := X"304200FF";
        ram_buffer(40230) := X"AFC2002C";
        ram_buffer(40231) := X"8E020030";
        ram_buffer(40232) := X"00000000";
        ram_buffer(40233) := X"10400020";
        ram_buffer(40234) := X"00000000";
        ram_buffer(40235) := X"8E030004";
        ram_buffer(40236) := X"8E020034";
        ram_buffer(40237) := X"00000000";
        ram_buffer(40238) := X"0062102A";
        ram_buffer(40239) := X"1440000A";
        ram_buffer(40240) := X"00000000";
        ram_buffer(40241) := X"02002821";
        ram_buffer(40242) := X"8FC40028";
        ram_buffer(40243) := X"0C029C71";
        ram_buffer(40244) := X"00000000";
        ram_buffer(40245) := X"10400004";
        ram_buffer(40246) := X"00000000";
        ram_buffer(40247) := X"2402FFFF";
        ram_buffer(40248) := X"10000043";
        ram_buffer(40249) := X"00000000";
        ram_buffer(40250) := X"8E020000";
        ram_buffer(40251) := X"00000000";
        ram_buffer(40252) := X"2442FFFF";
        ram_buffer(40253) := X"AE020000";
        ram_buffer(40254) := X"8E020000";
        ram_buffer(40255) := X"8FC3002C";
        ram_buffer(40256) := X"00000000";
        ram_buffer(40257) := X"306300FF";
        ram_buffer(40258) := X"A0430000";
        ram_buffer(40259) := X"8E020004";
        ram_buffer(40260) := X"00000000";
        ram_buffer(40261) := X"24420001";
        ram_buffer(40262) := X"AE020004";
        ram_buffer(40263) := X"8FC2002C";
        ram_buffer(40264) := X"10000033";
        ram_buffer(40265) := X"00000000";
        ram_buffer(40266) := X"8E020010";
        ram_buffer(40267) := X"00000000";
        ram_buffer(40268) := X"1040001C";
        ram_buffer(40269) := X"00000000";
        ram_buffer(40270) := X"8E030000";
        ram_buffer(40271) := X"8E020010";
        ram_buffer(40272) := X"00000000";
        ram_buffer(40273) := X"0043102B";
        ram_buffer(40274) := X"10400016";
        ram_buffer(40275) := X"00000000";
        ram_buffer(40276) := X"8E020000";
        ram_buffer(40277) := X"00000000";
        ram_buffer(40278) := X"2442FFFF";
        ram_buffer(40279) := X"90420000";
        ram_buffer(40280) := X"00000000";
        ram_buffer(40281) := X"00401821";
        ram_buffer(40282) := X"8FC2002C";
        ram_buffer(40283) := X"00000000";
        ram_buffer(40284) := X"1462000C";
        ram_buffer(40285) := X"00000000";
        ram_buffer(40286) := X"8E020000";
        ram_buffer(40287) := X"00000000";
        ram_buffer(40288) := X"2442FFFF";
        ram_buffer(40289) := X"AE020000";
        ram_buffer(40290) := X"8E020004";
        ram_buffer(40291) := X"00000000";
        ram_buffer(40292) := X"24420001";
        ram_buffer(40293) := X"AE020004";
        ram_buffer(40294) := X"8FC2002C";
        ram_buffer(40295) := X"10000014";
        ram_buffer(40296) := X"00000000";
        ram_buffer(40297) := X"8E020004";
        ram_buffer(40298) := X"00000000";
        ram_buffer(40299) := X"AE02003C";
        ram_buffer(40300) := X"8E020000";
        ram_buffer(40301) := X"00000000";
        ram_buffer(40302) := X"AE020038";
        ram_buffer(40303) := X"26020040";
        ram_buffer(40304) := X"AE020030";
        ram_buffer(40305) := X"24020003";
        ram_buffer(40306) := X"AE020034";
        ram_buffer(40307) := X"8FC2002C";
        ram_buffer(40308) := X"00000000";
        ram_buffer(40309) := X"304200FF";
        ram_buffer(40310) := X"A2020042";
        ram_buffer(40311) := X"26020042";
        ram_buffer(40312) := X"AE020000";
        ram_buffer(40313) := X"24020001";
        ram_buffer(40314) := X"AE020004";
        ram_buffer(40315) := X"8FC2002C";
        ram_buffer(40316) := X"03C0E821";
        ram_buffer(40317) := X"8FBF0024";
        ram_buffer(40318) := X"8FBE0020";
        ram_buffer(40319) := X"8FB0001C";
        ram_buffer(40320) := X"27BD0028";
        ram_buffer(40321) := X"03E00008";
        ram_buffer(40322) := X"00000000";
        ram_buffer(40323) := X"27BDFFE8";
        ram_buffer(40324) := X"AFBF0014";
        ram_buffer(40325) := X"AFBE0010";
        ram_buffer(40326) := X"03A0F021";
        ram_buffer(40327) := X"AFC40018";
        ram_buffer(40328) := X"00A01821";
        ram_buffer(40329) := X"8F828098";
        ram_buffer(40330) := X"00603021";
        ram_buffer(40331) := X"8FC50018";
        ram_buffer(40332) := X"00402021";
        ram_buffer(40333) := X"0C029CC2";
        ram_buffer(40334) := X"00000000";
        ram_buffer(40335) := X"03C0E821";
        ram_buffer(40336) := X"8FBF0014";
        ram_buffer(40337) := X"8FBE0010";
        ram_buffer(40338) := X"27BD0018";
        ram_buffer(40339) := X"03E00008";
        ram_buffer(40340) := X"00000000";
        ram_buffer(40341) := X"27BDFB70";
        ram_buffer(40342) := X"AFBF048C";
        ram_buffer(40343) := X"AFBE0488";
        ram_buffer(40344) := X"AFB00484";
        ram_buffer(40345) := X"03A0F021";
        ram_buffer(40346) := X"AFC40490";
        ram_buffer(40347) := X"00A08021";
        ram_buffer(40348) := X"AFC60498";
        ram_buffer(40349) := X"AFC7049C";
        ram_buffer(40350) := X"8603000C";
        ram_buffer(40351) := X"2402FFFD";
        ram_buffer(40352) := X"00621024";
        ram_buffer(40353) := X"00021400";
        ram_buffer(40354) := X"00021403";
        ram_buffer(40355) := X"A7C20020";
        ram_buffer(40356) := X"8E020064";
        ram_buffer(40357) := X"00000000";
        ram_buffer(40358) := X"AFC20078";
        ram_buffer(40359) := X"8602000E";
        ram_buffer(40360) := X"00000000";
        ram_buffer(40361) := X"A7C20022";
        ram_buffer(40362) := X"8E02001C";
        ram_buffer(40363) := X"00000000";
        ram_buffer(40364) := X"AFC20030";
        ram_buffer(40365) := X"8E020024";
        ram_buffer(40366) := X"00000000";
        ram_buffer(40367) := X"AFC20038";
        ram_buffer(40368) := X"27C2007C";
        ram_buffer(40369) := X"AFC20014";
        ram_buffer(40370) := X"8FC20014";
        ram_buffer(40371) := X"00000000";
        ram_buffer(40372) := X"AFC20024";
        ram_buffer(40373) := X"24020400";
        ram_buffer(40374) := X"AFC2001C";
        ram_buffer(40375) := X"8FC2001C";
        ram_buffer(40376) := X"00000000";
        ram_buffer(40377) := X"AFC20028";
        ram_buffer(40378) := X"AFC0002C";
        ram_buffer(40379) := X"27C20014";
        ram_buffer(40380) := X"8FC7049C";
        ram_buffer(40381) := X"8FC60498";
        ram_buffer(40382) := X"00402821";
        ram_buffer(40383) := X"8FC40490";
        ram_buffer(40384) := X"0C029DFA";
        ram_buffer(40385) := X"00000000";
        ram_buffer(40386) := X"AFC20010";
        ram_buffer(40387) := X"8FC20010";
        ram_buffer(40388) := X"00000000";
        ram_buffer(40389) := X"0440000A";
        ram_buffer(40390) := X"00000000";
        ram_buffer(40391) := X"27C20014";
        ram_buffer(40392) := X"00402821";
        ram_buffer(40393) := X"8FC40490";
        ram_buffer(40394) := X"0C026EE1";
        ram_buffer(40395) := X"00000000";
        ram_buffer(40396) := X"10400003";
        ram_buffer(40397) := X"00000000";
        ram_buffer(40398) := X"2402FFFF";
        ram_buffer(40399) := X"AFC20010";
        ram_buffer(40400) := X"87C20020";
        ram_buffer(40401) := X"00000000";
        ram_buffer(40402) := X"3042FFFF";
        ram_buffer(40403) := X"30420040";
        ram_buffer(40404) := X"10400007";
        ram_buffer(40405) := X"00000000";
        ram_buffer(40406) := X"8602000C";
        ram_buffer(40407) := X"00000000";
        ram_buffer(40408) := X"34420040";
        ram_buffer(40409) := X"00021400";
        ram_buffer(40410) := X"00021403";
        ram_buffer(40411) := X"A602000C";
        ram_buffer(40412) := X"8FC20010";
        ram_buffer(40413) := X"03C0E821";
        ram_buffer(40414) := X"8FBF048C";
        ram_buffer(40415) := X"8FBE0488";
        ram_buffer(40416) := X"8FB00484";
        ram_buffer(40417) := X"27BD0490";
        ram_buffer(40418) := X"03E00008";
        ram_buffer(40419) := X"00000000";
        ram_buffer(40420) := X"27BDFFE0";
        ram_buffer(40421) := X"AFBF001C";
        ram_buffer(40422) := X"AFBE0018";
        ram_buffer(40423) := X"03A0F021";
        ram_buffer(40424) := X"AFC40020";
        ram_buffer(40425) := X"AFC50024";
        ram_buffer(40426) := X"AFC60028";
        ram_buffer(40427) := X"8F828098";
        ram_buffer(40428) := X"8FC70028";
        ram_buffer(40429) := X"8FC60024";
        ram_buffer(40430) := X"8FC50020";
        ram_buffer(40431) := X"00402021";
        ram_buffer(40432) := X"0C029DFA";
        ram_buffer(40433) := X"00000000";
        ram_buffer(40434) := X"AFC20010";
        ram_buffer(40435) := X"8FC20010";
        ram_buffer(40436) := X"03C0E821";
        ram_buffer(40437) := X"8FBF001C";
        ram_buffer(40438) := X"8FBE0018";
        ram_buffer(40439) := X"27BD0020";
        ram_buffer(40440) := X"03E00008";
        ram_buffer(40441) := X"00000000";
        ram_buffer(40442) := X"27BDFE18";
        ram_buffer(40443) := X"AFBF01E4";
        ram_buffer(40444) := X"AFBE01E0";
        ram_buffer(40445) := X"AFB701DC";
        ram_buffer(40446) := X"AFB601D8";
        ram_buffer(40447) := X"AFB501D4";
        ram_buffer(40448) := X"AFB401D0";
        ram_buffer(40449) := X"AFB301CC";
        ram_buffer(40450) := X"AFB201C8";
        ram_buffer(40451) := X"AFB101C4";
        ram_buffer(40452) := X"AFB001C0";
        ram_buffer(40453) := X"03A0F021";
        ram_buffer(40454) := X"AFC401E8";
        ram_buffer(40455) := X"AFC501EC";
        ram_buffer(40456) := X"AFC601F0";
        ram_buffer(40457) := X"AFC701F4";
        ram_buffer(40458) := X"AFC0003C";
        ram_buffer(40459) := X"AFC00040";
        ram_buffer(40460) := X"AFC00044";
        ram_buffer(40461) := X"8FC401E8";
        ram_buffer(40462) := X"0C02BB25";
        ram_buffer(40463) := X"00000000";
        ram_buffer(40464) := X"8C420000";
        ram_buffer(40465) := X"00000000";
        ram_buffer(40466) := X"AFC20084";
        ram_buffer(40467) := X"8FC40084";
        ram_buffer(40468) := X"0C02851E";
        ram_buffer(40469) := X"00000000";
        ram_buffer(40470) := X"AFC20088";
        ram_buffer(40471) := X"00001821";
        ram_buffer(40472) := X"00001021";
        ram_buffer(40473) := X"AFC300A4";
        ram_buffer(40474) := X"AFC200A0";
        ram_buffer(40475) := X"AFC00048";
        ram_buffer(40476) := X"AFC000B4";
        ram_buffer(40477) := X"AFC00070";
        ram_buffer(40478) := X"AFC00074";
        ram_buffer(40479) := X"8FC201E8";
        ram_buffer(40480) := X"00000000";
        ram_buffer(40481) := X"AFC2008C";
        ram_buffer(40482) := X"8FC2008C";
        ram_buffer(40483) := X"00000000";
        ram_buffer(40484) := X"1040000A";
        ram_buffer(40485) := X"00000000";
        ram_buffer(40486) := X"8FC2008C";
        ram_buffer(40487) := X"00000000";
        ram_buffer(40488) := X"8C420038";
        ram_buffer(40489) := X"00000000";
        ram_buffer(40490) := X"14400004";
        ram_buffer(40491) := X"00000000";
        ram_buffer(40492) := X"8FC4008C";
        ram_buffer(40493) := X"0C027069";
        ram_buffer(40494) := X"00000000";
        ram_buffer(40495) := X"8FC201EC";
        ram_buffer(40496) := X"00000000";
        ram_buffer(40497) := X"8442000C";
        ram_buffer(40498) := X"00000000";
        ram_buffer(40499) := X"3042FFFF";
        ram_buffer(40500) := X"30422000";
        ram_buffer(40501) := X"14400013";
        ram_buffer(40502) := X"00000000";
        ram_buffer(40503) := X"8FC201EC";
        ram_buffer(40504) := X"00000000";
        ram_buffer(40505) := X"8442000C";
        ram_buffer(40506) := X"00000000";
        ram_buffer(40507) := X"34422000";
        ram_buffer(40508) := X"00021C00";
        ram_buffer(40509) := X"00031C03";
        ram_buffer(40510) := X"8FC201EC";
        ram_buffer(40511) := X"00000000";
        ram_buffer(40512) := X"A443000C";
        ram_buffer(40513) := X"8FC201EC";
        ram_buffer(40514) := X"00000000";
        ram_buffer(40515) := X"8C430064";
        ram_buffer(40516) := X"2402DFFF";
        ram_buffer(40517) := X"00621824";
        ram_buffer(40518) := X"8FC201EC";
        ram_buffer(40519) := X"00000000";
        ram_buffer(40520) := X"AC430064";
        ram_buffer(40521) := X"8FC201EC";
        ram_buffer(40522) := X"00000000";
        ram_buffer(40523) := X"8442000C";
        ram_buffer(40524) := X"00000000";
        ram_buffer(40525) := X"3042FFFF";
        ram_buffer(40526) := X"30420008";
        ram_buffer(40527) := X"10400007";
        ram_buffer(40528) := X"00000000";
        ram_buffer(40529) := X"8FC201EC";
        ram_buffer(40530) := X"00000000";
        ram_buffer(40531) := X"8C420010";
        ram_buffer(40532) := X"00000000";
        ram_buffer(40533) := X"1440000A";
        ram_buffer(40534) := X"00000000";
        ram_buffer(40535) := X"8FC501EC";
        ram_buffer(40536) := X"8FC401E8";
        ram_buffer(40537) := X"0C02ACF1";
        ram_buffer(40538) := X"00000000";
        ram_buffer(40539) := X"10400004";
        ram_buffer(40540) := X"00000000";
        ram_buffer(40541) := X"2402FFFF";
        ram_buffer(40542) := X"10000C68";
        ram_buffer(40543) := X"00000000";
        ram_buffer(40544) := X"8FC201EC";
        ram_buffer(40545) := X"00000000";
        ram_buffer(40546) := X"8442000C";
        ram_buffer(40547) := X"00000000";
        ram_buffer(40548) := X"3042FFFF";
        ram_buffer(40549) := X"3043001A";
        ram_buffer(40550) := X"2402000A";
        ram_buffer(40551) := X"1462000F";
        ram_buffer(40552) := X"00000000";
        ram_buffer(40553) := X"8FC201EC";
        ram_buffer(40554) := X"00000000";
        ram_buffer(40555) := X"8442000E";
        ram_buffer(40556) := X"00000000";
        ram_buffer(40557) := X"04400009";
        ram_buffer(40558) := X"00000000";
        ram_buffer(40559) := X"8FC701F4";
        ram_buffer(40560) := X"8FC601F0";
        ram_buffer(40561) := X"8FC501EC";
        ram_buffer(40562) := X"8FC401E8";
        ram_buffer(40563) := X"0C029D95";
        ram_buffer(40564) := X"00000000";
        ram_buffer(40565) := X"10000C51";
        ram_buffer(40566) := X"00000000";
        ram_buffer(40567) := X"8FD501F0";
        ram_buffer(40568) := X"27D000C4";
        ram_buffer(40569) := X"AFD000B8";
        ram_buffer(40570) := X"AFC000C0";
        ram_buffer(40571) := X"AFC000BC";
        ram_buffer(40572) := X"AFC00030";
        ram_buffer(40573) := X"02A09821";
        ram_buffer(40574) := X"10000002";
        ram_buffer(40575) := X"00000000";
        ram_buffer(40576) := X"26B50001";
        ram_buffer(40577) := X"82A20000";
        ram_buffer(40578) := X"00000000";
        ram_buffer(40579) := X"10400005";
        ram_buffer(40580) := X"00000000";
        ram_buffer(40581) := X"82A30000";
        ram_buffer(40582) := X"24020025";
        ram_buffer(40583) := X"1462FFF8";
        ram_buffer(40584) := X"00000000";
        ram_buffer(40585) := X"02A01821";
        ram_buffer(40586) := X"02601021";
        ram_buffer(40587) := X"00628823";
        ram_buffer(40588) := X"1220001F";
        ram_buffer(40589) := X"00000000";
        ram_buffer(40590) := X"AE130000";
        ram_buffer(40591) := X"02201021";
        ram_buffer(40592) := X"AE020004";
        ram_buffer(40593) := X"8FC300C0";
        ram_buffer(40594) := X"02201021";
        ram_buffer(40595) := X"00621021";
        ram_buffer(40596) := X"AFC200C0";
        ram_buffer(40597) := X"26100008";
        ram_buffer(40598) := X"8FC200BC";
        ram_buffer(40599) := X"00000000";
        ram_buffer(40600) := X"24420001";
        ram_buffer(40601) := X"AFC200BC";
        ram_buffer(40602) := X"8FC200BC";
        ram_buffer(40603) := X"00000000";
        ram_buffer(40604) := X"28420008";
        ram_buffer(40605) := X"1440000A";
        ram_buffer(40606) := X"00000000";
        ram_buffer(40607) := X"27C200B8";
        ram_buffer(40608) := X"00403021";
        ram_buffer(40609) := X"8FC501EC";
        ram_buffer(40610) := X"8FC401E8";
        ram_buffer(40611) := X"0C02EAF5";
        ram_buffer(40612) := X"00000000";
        ram_buffer(40613) := X"14400B93";
        ram_buffer(40614) := X"00000000";
        ram_buffer(40615) := X"27D000C4";
        ram_buffer(40616) := X"8FC20030";
        ram_buffer(40617) := X"00000000";
        ram_buffer(40618) := X"00511021";
        ram_buffer(40619) := X"AFC20030";
        ram_buffer(40620) := X"82A20000";
        ram_buffer(40621) := X"00000000";
        ram_buffer(40622) := X"10400B76";
        ram_buffer(40623) := X"00000000";
        ram_buffer(40624) := X"AFD50090";
        ram_buffer(40625) := X"26B50001";
        ram_buffer(40626) := X"00009021";
        ram_buffer(40627) := X"AFC00064";
        ram_buffer(40628) := X"AFC00034";
        ram_buffer(40629) := X"2402FFFF";
        ram_buffer(40630) := X"AFC20038";
        ram_buffer(40631) := X"A3C0009C";
        ram_buffer(40632) := X"AFC0004C";
        ram_buffer(40633) := X"AFC00054";
        ram_buffer(40634) := X"8FC20054";
        ram_buffer(40635) := X"00000000";
        ram_buffer(40636) := X"AFC20050";
        ram_buffer(40637) := X"02A01021";
        ram_buffer(40638) := X"24550001";
        ram_buffer(40639) := X"80420000";
        ram_buffer(40640) := X"00000000";
        ram_buffer(40641) := X"0040A021";
        ram_buffer(40642) := X"2683FFE0";
        ram_buffer(40643) := X"2C62005B";
        ram_buffer(40644) := X"1040055B";
        ram_buffer(40645) := X"00000000";
        ram_buffer(40646) := X"00031880";
        ram_buffer(40647) := X"3C02100D";
        ram_buffer(40648) := X"2442A764";
        ram_buffer(40649) := X"00621021";
        ram_buffer(40650) := X"8C420000";
        ram_buffer(40651) := X"00000000";
        ram_buffer(40652) := X"00400008";
        ram_buffer(40653) := X"00000000";
        ram_buffer(40654) := X"8FC401E8";
        ram_buffer(40655) := X"0C02BB25";
        ram_buffer(40656) := X"00000000";
        ram_buffer(40657) := X"8C420004";
        ram_buffer(40658) := X"00000000";
        ram_buffer(40659) := X"AFC2003C";
        ram_buffer(40660) := X"8FC4003C";
        ram_buffer(40661) := X"0C02851E";
        ram_buffer(40662) := X"00000000";
        ram_buffer(40663) := X"AFC20040";
        ram_buffer(40664) := X"8FC401E8";
        ram_buffer(40665) := X"0C02BB25";
        ram_buffer(40666) := X"00000000";
        ram_buffer(40667) := X"8C420008";
        ram_buffer(40668) := X"00000000";
        ram_buffer(40669) := X"AFC20044";
        ram_buffer(40670) := X"8FC20040";
        ram_buffer(40671) := X"00000000";
        ram_buffer(40672) := X"1040FFDC";
        ram_buffer(40673) := X"00000000";
        ram_buffer(40674) := X"8FC20044";
        ram_buffer(40675) := X"00000000";
        ram_buffer(40676) := X"1040FFD8";
        ram_buffer(40677) := X"00000000";
        ram_buffer(40678) := X"8FC20044";
        ram_buffer(40679) := X"00000000";
        ram_buffer(40680) := X"80420000";
        ram_buffer(40681) := X"00000000";
        ram_buffer(40682) := X"1040FFD2";
        ram_buffer(40683) := X"00000000";
        ram_buffer(40684) := X"36520400";
        ram_buffer(40685) := X"1000FFCF";
        ram_buffer(40686) := X"00000000";
        ram_buffer(40687) := X"83C2009C";
        ram_buffer(40688) := X"00000000";
        ram_buffer(40689) := X"1440FFCB";
        ram_buffer(40690) := X"00000000";
        ram_buffer(40691) := X"24020020";
        ram_buffer(40692) := X"A3C2009C";
        ram_buffer(40693) := X"1000FFC7";
        ram_buffer(40694) := X"00000000";
        ram_buffer(40695) := X"36520001";
        ram_buffer(40696) := X"1000FFC4";
        ram_buffer(40697) := X"00000000";
        ram_buffer(40698) := X"8FC301F4";
        ram_buffer(40699) := X"00000000";
        ram_buffer(40700) := X"24620004";
        ram_buffer(40701) := X"AFC201F4";
        ram_buffer(40702) := X"8C620000";
        ram_buffer(40703) := X"00000000";
        ram_buffer(40704) := X"AFC20034";
        ram_buffer(40705) := X"8FC20034";
        ram_buffer(40706) := X"00000000";
        ram_buffer(40707) := X"04400003";
        ram_buffer(40708) := X"00000000";
        ram_buffer(40709) := X"1000FFB7";
        ram_buffer(40710) := X"00000000";
        ram_buffer(40711) := X"8FC20034";
        ram_buffer(40712) := X"00000000";
        ram_buffer(40713) := X"00021023";
        ram_buffer(40714) := X"AFC20034";
        ram_buffer(40715) := X"36520004";
        ram_buffer(40716) := X"1000FFB0";
        ram_buffer(40717) := X"00000000";
        ram_buffer(40718) := X"2402002B";
        ram_buffer(40719) := X"A3C2009C";
        ram_buffer(40720) := X"1000FFAC";
        ram_buffer(40721) := X"00000000";
        ram_buffer(40722) := X"02A01021";
        ram_buffer(40723) := X"24550001";
        ram_buffer(40724) := X"80420000";
        ram_buffer(40725) := X"00000000";
        ram_buffer(40726) := X"0040A021";
        ram_buffer(40727) := X"2402002A";
        ram_buffer(40728) := X"16820010";
        ram_buffer(40729) := X"00000000";
        ram_buffer(40730) := X"8FC301F4";
        ram_buffer(40731) := X"00000000";
        ram_buffer(40732) := X"24620004";
        ram_buffer(40733) := X"AFC201F4";
        ram_buffer(40734) := X"8C620000";
        ram_buffer(40735) := X"00000000";
        ram_buffer(40736) := X"AFC20038";
        ram_buffer(40737) := X"8FC20038";
        ram_buffer(40738) := X"00000000";
        ram_buffer(40739) := X"0441FF99";
        ram_buffer(40740) := X"00000000";
        ram_buffer(40741) := X"2402FFFF";
        ram_buffer(40742) := X"AFC20038";
        ram_buffer(40743) := X"1000FF95";
        ram_buffer(40744) := X"00000000";
        ram_buffer(40745) := X"00008821";
        ram_buffer(40746) := X"1000000D";
        ram_buffer(40747) := X"00000000";
        ram_buffer(40748) := X"02201821";
        ram_buffer(40749) := X"00031040";
        ram_buffer(40750) := X"00401821";
        ram_buffer(40751) := X"00031080";
        ram_buffer(40752) := X"00621821";
        ram_buffer(40753) := X"2682FFD0";
        ram_buffer(40754) := X"00628821";
        ram_buffer(40755) := X"02A01021";
        ram_buffer(40756) := X"24550001";
        ram_buffer(40757) := X"80420000";
        ram_buffer(40758) := X"00000000";
        ram_buffer(40759) := X"0040A021";
        ram_buffer(40760) := X"2682FFD0";
        ram_buffer(40761) := X"2C42000A";
        ram_buffer(40762) := X"1440FFF1";
        ram_buffer(40763) := X"00000000";
        ram_buffer(40764) := X"02201021";
        ram_buffer(40765) := X"04410002";
        ram_buffer(40766) := X"00000000";
        ram_buffer(40767) := X"2402FFFF";
        ram_buffer(40768) := X"AFC20038";
        ram_buffer(40769) := X"1000FF80";
        ram_buffer(40770) := X"00000000";
        ram_buffer(40771) := X"36520080";
        ram_buffer(40772) := X"1000FF78";
        ram_buffer(40773) := X"00000000";
        ram_buffer(40774) := X"00008821";
        ram_buffer(40775) := X"02201821";
        ram_buffer(40776) := X"00031040";
        ram_buffer(40777) := X"00401821";
        ram_buffer(40778) := X"00031080";
        ram_buffer(40779) := X"00621821";
        ram_buffer(40780) := X"2682FFD0";
        ram_buffer(40781) := X"00628821";
        ram_buffer(40782) := X"02A01021";
        ram_buffer(40783) := X"24550001";
        ram_buffer(40784) := X"80420000";
        ram_buffer(40785) := X"00000000";
        ram_buffer(40786) := X"0040A021";
        ram_buffer(40787) := X"2682FFD0";
        ram_buffer(40788) := X"2C42000A";
        ram_buffer(40789) := X"1440FFF1";
        ram_buffer(40790) := X"00000000";
        ram_buffer(40791) := X"AFD10034";
        ram_buffer(40792) := X"1000FF69";
        ram_buffer(40793) := X"00000000";
        ram_buffer(40794) := X"36520008";
        ram_buffer(40795) := X"1000FF61";
        ram_buffer(40796) := X"00000000";
        ram_buffer(40797) := X"82A30000";
        ram_buffer(40798) := X"24020068";
        ram_buffer(40799) := X"14620005";
        ram_buffer(40800) := X"00000000";
        ram_buffer(40801) := X"26B50001";
        ram_buffer(40802) := X"36520200";
        ram_buffer(40803) := X"1000FF59";
        ram_buffer(40804) := X"00000000";
        ram_buffer(40805) := X"36520040";
        ram_buffer(40806) := X"1000FF56";
        ram_buffer(40807) := X"00000000";
        ram_buffer(40808) := X"82A30000";
        ram_buffer(40809) := X"2402006C";
        ram_buffer(40810) := X"14620005";
        ram_buffer(40811) := X"00000000";
        ram_buffer(40812) := X"26B50001";
        ram_buffer(40813) := X"36520020";
        ram_buffer(40814) := X"1000FF4E";
        ram_buffer(40815) := X"00000000";
        ram_buffer(40816) := X"36520010";
        ram_buffer(40817) := X"1000FF4B";
        ram_buffer(40818) := X"00000000";
        ram_buffer(40819) := X"36520020";
        ram_buffer(40820) := X"1000FF48";
        ram_buffer(40821) := X"00000000";
        ram_buffer(40822) := X"36520020";
        ram_buffer(40823) := X"1000FF45";
        ram_buffer(40824) := X"00000000";
        ram_buffer(40825) := X"27D30104";
        ram_buffer(40826) := X"8FC301F4";
        ram_buffer(40827) := X"00000000";
        ram_buffer(40828) := X"24620004";
        ram_buffer(40829) := X"AFC201F4";
        ram_buffer(40830) := X"8C620000";
        ram_buffer(40831) := X"00000000";
        ram_buffer(40832) := X"00021600";
        ram_buffer(40833) := X"00021603";
        ram_buffer(40834) := X"A2620000";
        ram_buffer(40835) := X"24020001";
        ram_buffer(40836) := X"AFC2006C";
        ram_buffer(40837) := X"A3C0009C";
        ram_buffer(40838) := X"100004A5";
        ram_buffer(40839) := X"00000000";
        ram_buffer(40840) := X"36520010";
        ram_buffer(40841) := X"32420020";
        ram_buffer(40842) := X"1040000E";
        ram_buffer(40843) := X"00000000";
        ram_buffer(40844) := X"8FC201F4";
        ram_buffer(40845) := X"00000000";
        ram_buffer(40846) := X"24430007";
        ram_buffer(40847) := X"2402FFF8";
        ram_buffer(40848) := X"00621024";
        ram_buffer(40849) := X"24430008";
        ram_buffer(40850) := X"AFC301F4";
        ram_buffer(40851) := X"8C430004";
        ram_buffer(40852) := X"8C420000";
        ram_buffer(40853) := X"AFC30174";
        ram_buffer(40854) := X"AFC20170";
        ram_buffer(40855) := X"10000038";
        ram_buffer(40856) := X"00000000";
        ram_buffer(40857) := X"32420010";
        ram_buffer(40858) := X"1040000C";
        ram_buffer(40859) := X"00000000";
        ram_buffer(40860) := X"8FC301F4";
        ram_buffer(40861) := X"00000000";
        ram_buffer(40862) := X"24620004";
        ram_buffer(40863) := X"AFC201F4";
        ram_buffer(40864) := X"8C620000";
        ram_buffer(40865) := X"00000000";
        ram_buffer(40866) := X"AFC20174";
        ram_buffer(40867) := X"000217C3";
        ram_buffer(40868) := X"AFC20170";
        ram_buffer(40869) := X"1000002A";
        ram_buffer(40870) := X"00000000";
        ram_buffer(40871) := X"32420040";
        ram_buffer(40872) := X"1040000E";
        ram_buffer(40873) := X"00000000";
        ram_buffer(40874) := X"8FC301F4";
        ram_buffer(40875) := X"00000000";
        ram_buffer(40876) := X"24620004";
        ram_buffer(40877) := X"AFC201F4";
        ram_buffer(40878) := X"8C620000";
        ram_buffer(40879) := X"00000000";
        ram_buffer(40880) := X"00021400";
        ram_buffer(40881) := X"00021403";
        ram_buffer(40882) := X"AFC20174";
        ram_buffer(40883) := X"000217C3";
        ram_buffer(40884) := X"AFC20170";
        ram_buffer(40885) := X"1000001A";
        ram_buffer(40886) := X"00000000";
        ram_buffer(40887) := X"32420200";
        ram_buffer(40888) := X"1040000E";
        ram_buffer(40889) := X"00000000";
        ram_buffer(40890) := X"8FC301F4";
        ram_buffer(40891) := X"00000000";
        ram_buffer(40892) := X"24620004";
        ram_buffer(40893) := X"AFC201F4";
        ram_buffer(40894) := X"8C620000";
        ram_buffer(40895) := X"00000000";
        ram_buffer(40896) := X"00021600";
        ram_buffer(40897) := X"00021603";
        ram_buffer(40898) := X"AFC20174";
        ram_buffer(40899) := X"000217C3";
        ram_buffer(40900) := X"AFC20170";
        ram_buffer(40901) := X"1000000A";
        ram_buffer(40902) := X"00000000";
        ram_buffer(40903) := X"8FC301F4";
        ram_buffer(40904) := X"00000000";
        ram_buffer(40905) := X"24620004";
        ram_buffer(40906) := X"AFC201F4";
        ram_buffer(40907) := X"8C620000";
        ram_buffer(40908) := X"00000000";
        ram_buffer(40909) := X"AFC20174";
        ram_buffer(40910) := X"000217C3";
        ram_buffer(40911) := X"AFC20170";
        ram_buffer(40912) := X"8FC30174";
        ram_buffer(40913) := X"8FC20170";
        ram_buffer(40914) := X"AFC3005C";
        ram_buffer(40915) := X"AFC20058";
        ram_buffer(40916) := X"8FC3005C";
        ram_buffer(40917) := X"8FC20058";
        ram_buffer(40918) := X"00000000";
        ram_buffer(40919) := X"0441000E";
        ram_buffer(40920) := X"00000000";
        ram_buffer(40921) := X"00001821";
        ram_buffer(40922) := X"00001021";
        ram_buffer(40923) := X"8FC5005C";
        ram_buffer(40924) := X"8FC40058";
        ram_buffer(40925) := X"00653823";
        ram_buffer(40926) := X"0067402B";
        ram_buffer(40927) := X"00443023";
        ram_buffer(40928) := X"00C81023";
        ram_buffer(40929) := X"00403021";
        ram_buffer(40930) := X"AFC7005C";
        ram_buffer(40931) := X"AFC60058";
        ram_buffer(40932) := X"2402002D";
        ram_buffer(40933) := X"A3C2009C";
        ram_buffer(40934) := X"24020001";
        ram_buffer(40935) := X"A3C20060";
        ram_buffer(40936) := X"10000344";
        ram_buffer(40937) := X"00000000";
        ram_buffer(40938) := X"32420008";
        ram_buffer(40939) := X"1040000F";
        ram_buffer(40940) := X"00000000";
        ram_buffer(40941) := X"8FC201F4";
        ram_buffer(40942) := X"00000000";
        ram_buffer(40943) := X"24430007";
        ram_buffer(40944) := X"2402FFF8";
        ram_buffer(40945) := X"00621824";
        ram_buffer(40946) := X"24620008";
        ram_buffer(40947) := X"AFC201F4";
        ram_buffer(40948) := X"8C620000";
        ram_buffer(40949) := X"8C630004";
        ram_buffer(40950) := X"00000000";
        ram_buffer(40951) := X"AFC300A4";
        ram_buffer(40952) := X"AFC200A0";
        ram_buffer(40953) := X"1000000D";
        ram_buffer(40954) := X"00000000";
        ram_buffer(40955) := X"8FC201F4";
        ram_buffer(40956) := X"00000000";
        ram_buffer(40957) := X"24430007";
        ram_buffer(40958) := X"2402FFF8";
        ram_buffer(40959) := X"00621824";
        ram_buffer(40960) := X"24620008";
        ram_buffer(40961) := X"AFC201F4";
        ram_buffer(40962) := X"8C620000";
        ram_buffer(40963) := X"8C630004";
        ram_buffer(40964) := X"00000000";
        ram_buffer(40965) := X"AFC300A4";
        ram_buffer(40966) := X"AFC200A0";
        ram_buffer(40967) := X"8FC300A4";
        ram_buffer(40968) := X"8FC200A0";
        ram_buffer(40969) := X"00602821";
        ram_buffer(40970) := X"00402021";
        ram_buffer(40971) := X"0C02CAED";
        ram_buffer(40972) := X"00000000";
        ram_buffer(40973) := X"00401821";
        ram_buffer(40974) := X"24020001";
        ram_buffer(40975) := X"1462001C";
        ram_buffer(40976) := X"00000000";
        ram_buffer(40977) := X"8FC300A4";
        ram_buffer(40978) := X"8FC200A0";
        ram_buffer(40979) := X"00003821";
        ram_buffer(40980) := X"00003021";
        ram_buffer(40981) := X"00602821";
        ram_buffer(40982) := X"00402021";
        ram_buffer(40983) := X"0C0316F7";
        ram_buffer(40984) := X"00000000";
        ram_buffer(40985) := X"04410003";
        ram_buffer(40986) := X"00000000";
        ram_buffer(40987) := X"2402002D";
        ram_buffer(40988) := X"A3C2009C";
        ram_buffer(40989) := X"2A820048";
        ram_buffer(40990) := X"10400005";
        ram_buffer(40991) := X"00000000";
        ram_buffer(40992) := X"3C02100D";
        ram_buffer(40993) := X"2453A704";
        ram_buffer(40994) := X"10000003";
        ram_buffer(40995) := X"00000000";
        ram_buffer(40996) := X"3C02100D";
        ram_buffer(40997) := X"2453A708";
        ram_buffer(40998) := X"24020003";
        ram_buffer(40999) := X"AFC2006C";
        ram_buffer(41000) := X"2402FF7F";
        ram_buffer(41001) := X"02429024";
        ram_buffer(41002) := X"10000401";
        ram_buffer(41003) := X"00000000";
        ram_buffer(41004) := X"8FC300A4";
        ram_buffer(41005) := X"8FC200A0";
        ram_buffer(41006) := X"00602821";
        ram_buffer(41007) := X"00402021";
        ram_buffer(41008) := X"0C02CAED";
        ram_buffer(41009) := X"00000000";
        ram_buffer(41010) := X"14400010";
        ram_buffer(41011) := X"00000000";
        ram_buffer(41012) := X"2A820048";
        ram_buffer(41013) := X"10400005";
        ram_buffer(41014) := X"00000000";
        ram_buffer(41015) := X"3C02100D";
        ram_buffer(41016) := X"2453A70C";
        ram_buffer(41017) := X"10000003";
        ram_buffer(41018) := X"00000000";
        ram_buffer(41019) := X"3C02100D";
        ram_buffer(41020) := X"2453A710";
        ram_buffer(41021) := X"24020003";
        ram_buffer(41022) := X"AFC2006C";
        ram_buffer(41023) := X"2402FF7F";
        ram_buffer(41024) := X"02429024";
        ram_buffer(41025) := X"100003EA";
        ram_buffer(41026) := X"00000000";
        ram_buffer(41027) := X"24020061";
        ram_buffer(41028) := X"12820004";
        ram_buffer(41029) := X"00000000";
        ram_buffer(41030) := X"24020041";
        ram_buffer(41031) := X"1682002F";
        ram_buffer(41032) := X"00000000";
        ram_buffer(41033) := X"24020030";
        ram_buffer(41034) := X"A3C20168";
        ram_buffer(41035) := X"24020061";
        ram_buffer(41036) := X"16820004";
        ram_buffer(41037) := X"00000000";
        ram_buffer(41038) := X"24020078";
        ram_buffer(41039) := X"10000002";
        ram_buffer(41040) := X"00000000";
        ram_buffer(41041) := X"24020058";
        ram_buffer(41042) := X"A3C20169";
        ram_buffer(41043) := X"36520002";
        ram_buffer(41044) := X"8FC20038";
        ram_buffer(41045) := X"00000000";
        ram_buffer(41046) := X"28420064";
        ram_buffer(41047) := X"1440001C";
        ram_buffer(41048) := X"00000000";
        ram_buffer(41049) := X"8FC20038";
        ram_buffer(41050) := X"00000000";
        ram_buffer(41051) := X"24420001";
        ram_buffer(41052) := X"00402821";
        ram_buffer(41053) := X"8FC401E8";
        ram_buffer(41054) := X"0C027B8F";
        ram_buffer(41055) := X"00000000";
        ram_buffer(41056) := X"AFC20074";
        ram_buffer(41057) := X"8FC20074";
        ram_buffer(41058) := X"00000000";
        ram_buffer(41059) := X"1440000D";
        ram_buffer(41060) := X"00000000";
        ram_buffer(41061) := X"8FC201EC";
        ram_buffer(41062) := X"00000000";
        ram_buffer(41063) := X"8442000C";
        ram_buffer(41064) := X"00000000";
        ram_buffer(41065) := X"34420040";
        ram_buffer(41066) := X"00021C00";
        ram_buffer(41067) := X"00031C03";
        ram_buffer(41068) := X"8FC201EC";
        ram_buffer(41069) := X"00000000";
        ram_buffer(41070) := X"A443000C";
        ram_buffer(41071) := X"10000A42";
        ram_buffer(41072) := X"00000000";
        ram_buffer(41073) := X"8FD30074";
        ram_buffer(41074) := X"10000018";
        ram_buffer(41075) := X"00000000";
        ram_buffer(41076) := X"27D30104";
        ram_buffer(41077) := X"10000015";
        ram_buffer(41078) := X"00000000";
        ram_buffer(41079) := X"8FC30038";
        ram_buffer(41080) := X"2402FFFF";
        ram_buffer(41081) := X"14620005";
        ram_buffer(41082) := X"00000000";
        ram_buffer(41083) := X"24020006";
        ram_buffer(41084) := X"AFC20038";
        ram_buffer(41085) := X"1000000D";
        ram_buffer(41086) := X"00000000";
        ram_buffer(41087) := X"24020067";
        ram_buffer(41088) := X"12820004";
        ram_buffer(41089) := X"00000000";
        ram_buffer(41090) := X"24020047";
        ram_buffer(41091) := X"16820007";
        ram_buffer(41092) := X"00000000";
        ram_buffer(41093) := X"8FC20038";
        ram_buffer(41094) := X"00000000";
        ram_buffer(41095) := X"14400003";
        ram_buffer(41096) := X"00000000";
        ram_buffer(41097) := X"24020001";
        ram_buffer(41098) := X"AFC20038";
        ram_buffer(41099) := X"36520100";
        ram_buffer(41100) := X"8FC500A4";
        ram_buffer(41101) := X"8FC400A0";
        ram_buffer(41102) := X"AFB30028";
        ram_buffer(41103) := X"27C200B4";
        ram_buffer(41104) := X"AFA20024";
        ram_buffer(41105) := X"AFB40020";
        ram_buffer(41106) := X"27C200A8";
        ram_buffer(41107) := X"AFA2001C";
        ram_buffer(41108) := X"27C2009D";
        ram_buffer(41109) := X"AFA20018";
        ram_buffer(41110) := X"AFB20014";
        ram_buffer(41111) := X"8FC20038";
        ram_buffer(41112) := X"00000000";
        ram_buffer(41113) := X"AFA20010";
        ram_buffer(41114) := X"00A03821";
        ram_buffer(41115) := X"00803021";
        ram_buffer(41116) := X"8FC401E8";
        ram_buffer(41117) := X"0C02AAD5";
        ram_buffer(41118) := X"00000000";
        ram_buffer(41119) := X"00409821";
        ram_buffer(41120) := X"24020067";
        ram_buffer(41121) := X"12820004";
        ram_buffer(41122) := X"00000000";
        ram_buffer(41123) := X"24020047";
        ram_buffer(41124) := X"16820012";
        ram_buffer(41125) := X"00000000";
        ram_buffer(41126) := X"8FC200A8";
        ram_buffer(41127) := X"00000000";
        ram_buffer(41128) := X"2842FFFD";
        ram_buffer(41129) := X"14400007";
        ram_buffer(41130) := X"00000000";
        ram_buffer(41131) := X"8FC300A8";
        ram_buffer(41132) := X"8FC20038";
        ram_buffer(41133) := X"00000000";
        ram_buffer(41134) := X"0043102A";
        ram_buffer(41135) := X"10400004";
        ram_buffer(41136) := X"00000000";
        ram_buffer(41137) := X"2694FFFE";
        ram_buffer(41138) := X"10000008";
        ram_buffer(41139) := X"00000000";
        ram_buffer(41140) := X"24140067";
        ram_buffer(41141) := X"10000005";
        ram_buffer(41142) := X"00000000";
        ram_buffer(41143) := X"24020046";
        ram_buffer(41144) := X"16820002";
        ram_buffer(41145) := X"00000000";
        ram_buffer(41146) := X"24140066";
        ram_buffer(41147) := X"2A820066";
        ram_buffer(41148) := X"10400022";
        ram_buffer(41149) := X"00000000";
        ram_buffer(41150) := X"8FC200A8";
        ram_buffer(41151) := X"00000000";
        ram_buffer(41152) := X"2442FFFF";
        ram_buffer(41153) := X"AFC200A8";
        ram_buffer(41154) := X"8FC300A8";
        ram_buffer(41155) := X"27C200AC";
        ram_buffer(41156) := X"02803021";
        ram_buffer(41157) := X"00602821";
        ram_buffer(41158) := X"00402021";
        ram_buffer(41159) := X"0C02AC3B";
        ram_buffer(41160) := X"00000000";
        ram_buffer(41161) := X"AFC20048";
        ram_buffer(41162) := X"8FC300B4";
        ram_buffer(41163) := X"8FC20048";
        ram_buffer(41164) := X"00000000";
        ram_buffer(41165) := X"00431021";
        ram_buffer(41166) := X"AFC2006C";
        ram_buffer(41167) := X"8FC200B4";
        ram_buffer(41168) := X"00000000";
        ram_buffer(41169) := X"28420002";
        ram_buffer(41170) := X"10400004";
        ram_buffer(41171) := X"00000000";
        ram_buffer(41172) := X"32420001";
        ram_buffer(41173) := X"10400005";
        ram_buffer(41174) := X"00000000";
        ram_buffer(41175) := X"8FC2006C";
        ram_buffer(41176) := X"00000000";
        ram_buffer(41177) := X"24420001";
        ram_buffer(41178) := X"AFC2006C";
        ram_buffer(41179) := X"2402FBFF";
        ram_buffer(41180) := X"02429024";
        ram_buffer(41181) := X"1000009D";
        ram_buffer(41182) := X"00000000";
        ram_buffer(41183) := X"24020066";
        ram_buffer(41184) := X"16820028";
        ram_buffer(41185) := X"00000000";
        ram_buffer(41186) := X"8FC200A8";
        ram_buffer(41187) := X"00000000";
        ram_buffer(41188) := X"18400014";
        ram_buffer(41189) := X"00000000";
        ram_buffer(41190) := X"8FC200A8";
        ram_buffer(41191) := X"00000000";
        ram_buffer(41192) := X"AFC2006C";
        ram_buffer(41193) := X"8FC20038";
        ram_buffer(41194) := X"00000000";
        ram_buffer(41195) := X"14400004";
        ram_buffer(41196) := X"00000000";
        ram_buffer(41197) := X"32420001";
        ram_buffer(41198) := X"1040003A";
        ram_buffer(41199) := X"00000000";
        ram_buffer(41200) := X"8FC20038";
        ram_buffer(41201) := X"00000000";
        ram_buffer(41202) := X"24430001";
        ram_buffer(41203) := X"8FC2006C";
        ram_buffer(41204) := X"00000000";
        ram_buffer(41205) := X"00431021";
        ram_buffer(41206) := X"AFC2006C";
        ram_buffer(41207) := X"10000031";
        ram_buffer(41208) := X"00000000";
        ram_buffer(41209) := X"8FC20038";
        ram_buffer(41210) := X"00000000";
        ram_buffer(41211) := X"14400004";
        ram_buffer(41212) := X"00000000";
        ram_buffer(41213) := X"32420001";
        ram_buffer(41214) := X"10400006";
        ram_buffer(41215) := X"00000000";
        ram_buffer(41216) := X"8FC20038";
        ram_buffer(41217) := X"00000000";
        ram_buffer(41218) := X"24420002";
        ram_buffer(41219) := X"10000002";
        ram_buffer(41220) := X"00000000";
        ram_buffer(41221) := X"24020001";
        ram_buffer(41222) := X"AFC2006C";
        ram_buffer(41223) := X"10000021";
        ram_buffer(41224) := X"00000000";
        ram_buffer(41225) := X"8FC300A8";
        ram_buffer(41226) := X"8FC200B4";
        ram_buffer(41227) := X"00000000";
        ram_buffer(41228) := X"0062102A";
        ram_buffer(41229) := X"1440000D";
        ram_buffer(41230) := X"00000000";
        ram_buffer(41231) := X"8FC200A8";
        ram_buffer(41232) := X"00000000";
        ram_buffer(41233) := X"AFC2006C";
        ram_buffer(41234) := X"32420001";
        ram_buffer(41235) := X"10400015";
        ram_buffer(41236) := X"00000000";
        ram_buffer(41237) := X"8FC2006C";
        ram_buffer(41238) := X"00000000";
        ram_buffer(41239) := X"24420001";
        ram_buffer(41240) := X"AFC2006C";
        ram_buffer(41241) := X"1000000F";
        ram_buffer(41242) := X"00000000";
        ram_buffer(41243) := X"8FC200A8";
        ram_buffer(41244) := X"00000000";
        ram_buffer(41245) := X"1C400006";
        ram_buffer(41246) := X"00000000";
        ram_buffer(41247) := X"8FC300A8";
        ram_buffer(41248) := X"24020002";
        ram_buffer(41249) := X"00431823";
        ram_buffer(41250) := X"10000002";
        ram_buffer(41251) := X"00000000";
        ram_buffer(41252) := X"24030001";
        ram_buffer(41253) := X"8FC200B4";
        ram_buffer(41254) := X"00000000";
        ram_buffer(41255) := X"00621021";
        ram_buffer(41256) := X"AFC2006C";
        ram_buffer(41257) := X"32420400";
        ram_buffer(41258) := X"1040004D";
        ram_buffer(41259) := X"00000000";
        ram_buffer(41260) := X"8FC200A8";
        ram_buffer(41261) := X"00000000";
        ram_buffer(41262) := X"18400049";
        ram_buffer(41263) := X"00000000";
        ram_buffer(41264) := X"AFC00054";
        ram_buffer(41265) := X"8FC20054";
        ram_buffer(41266) := X"00000000";
        ram_buffer(41267) := X"AFC20050";
        ram_buffer(41268) := X"8FC200A8";
        ram_buffer(41269) := X"00000000";
        ram_buffer(41270) := X"AFC2004C";
        ram_buffer(41271) := X"10000029";
        ram_buffer(41272) := X"00000000";
        ram_buffer(41273) := X"8FC20044";
        ram_buffer(41274) := X"00000000";
        ram_buffer(41275) := X"80420000";
        ram_buffer(41276) := X"00000000";
        ram_buffer(41277) := X"00401821";
        ram_buffer(41278) := X"8FC2004C";
        ram_buffer(41279) := X"00000000";
        ram_buffer(41280) := X"0062102A";
        ram_buffer(41281) := X"10400027";
        ram_buffer(41282) := X"00000000";
        ram_buffer(41283) := X"8FC20044";
        ram_buffer(41284) := X"00000000";
        ram_buffer(41285) := X"80420000";
        ram_buffer(41286) := X"00000000";
        ram_buffer(41287) := X"00401821";
        ram_buffer(41288) := X"8FC2004C";
        ram_buffer(41289) := X"00000000";
        ram_buffer(41290) := X"00431023";
        ram_buffer(41291) := X"AFC2004C";
        ram_buffer(41292) := X"8FC20044";
        ram_buffer(41293) := X"00000000";
        ram_buffer(41294) := X"24420001";
        ram_buffer(41295) := X"80420000";
        ram_buffer(41296) := X"00000000";
        ram_buffer(41297) := X"1040000B";
        ram_buffer(41298) := X"00000000";
        ram_buffer(41299) := X"8FC20050";
        ram_buffer(41300) := X"00000000";
        ram_buffer(41301) := X"24420001";
        ram_buffer(41302) := X"AFC20050";
        ram_buffer(41303) := X"8FC20044";
        ram_buffer(41304) := X"00000000";
        ram_buffer(41305) := X"24420001";
        ram_buffer(41306) := X"AFC20044";
        ram_buffer(41307) := X"10000005";
        ram_buffer(41308) := X"00000000";
        ram_buffer(41309) := X"8FC20054";
        ram_buffer(41310) := X"00000000";
        ram_buffer(41311) := X"24420001";
        ram_buffer(41312) := X"AFC20054";
        ram_buffer(41313) := X"8FC20044";
        ram_buffer(41314) := X"00000000";
        ram_buffer(41315) := X"80430000";
        ram_buffer(41316) := X"2402007F";
        ram_buffer(41317) := X"1462FFD3";
        ram_buffer(41318) := X"00000000";
        ram_buffer(41319) := X"10000002";
        ram_buffer(41320) := X"00000000";
        ram_buffer(41321) := X"00000000";
        ram_buffer(41322) := X"8FC30050";
        ram_buffer(41323) := X"8FC20054";
        ram_buffer(41324) := X"00000000";
        ram_buffer(41325) := X"00621021";
        ram_buffer(41326) := X"00401821";
        ram_buffer(41327) := X"8FC20040";
        ram_buffer(41328) := X"00000000";
        ram_buffer(41329) := X"00620018";
        ram_buffer(41330) := X"8FC2006C";
        ram_buffer(41331) := X"00001812";
        ram_buffer(41332) := X"00621021";
        ram_buffer(41333) := X"AFC2006C";
        ram_buffer(41334) := X"10000004";
        ram_buffer(41335) := X"00000000";
        ram_buffer(41336) := X"8FC200A8";
        ram_buffer(41337) := X"00000000";
        ram_buffer(41338) := X"AFC2004C";
        ram_buffer(41339) := X"83C2009D";
        ram_buffer(41340) := X"00000000";
        ram_buffer(41341) := X"104002AD";
        ram_buffer(41342) := X"00000000";
        ram_buffer(41343) := X"2402002D";
        ram_buffer(41344) := X"A3C2009C";
        ram_buffer(41345) := X"100002A9";
        ram_buffer(41346) := X"00000000";
        ram_buffer(41347) := X"32420020";
        ram_buffer(41348) := X"10400011";
        ram_buffer(41349) := X"00000000";
        ram_buffer(41350) := X"8FC201F4";
        ram_buffer(41351) := X"00000000";
        ram_buffer(41352) := X"24430004";
        ram_buffer(41353) := X"AFC301F4";
        ram_buffer(41354) := X"8C430000";
        ram_buffer(41355) := X"8FC20030";
        ram_buffer(41356) := X"00000000";
        ram_buffer(41357) := X"AFC2018C";
        ram_buffer(41358) := X"000217C3";
        ram_buffer(41359) := X"AFC20188";
        ram_buffer(41360) := X"8FC5018C";
        ram_buffer(41361) := X"8FC40188";
        ram_buffer(41362) := X"AC650004";
        ram_buffer(41363) := X"AC640000";
        ram_buffer(41364) := X"1000088E";
        ram_buffer(41365) := X"00000000";
        ram_buffer(41366) := X"32420010";
        ram_buffer(41367) := X"1040000B";
        ram_buffer(41368) := X"00000000";
        ram_buffer(41369) := X"8FC201F4";
        ram_buffer(41370) := X"00000000";
        ram_buffer(41371) := X"24430004";
        ram_buffer(41372) := X"AFC301F4";
        ram_buffer(41373) := X"8C420000";
        ram_buffer(41374) := X"8FC30030";
        ram_buffer(41375) := X"00000000";
        ram_buffer(41376) := X"AC430000";
        ram_buffer(41377) := X"10000881";
        ram_buffer(41378) := X"00000000";
        ram_buffer(41379) := X"32420040";
        ram_buffer(41380) := X"1040000D";
        ram_buffer(41381) := X"00000000";
        ram_buffer(41382) := X"8FC201F4";
        ram_buffer(41383) := X"00000000";
        ram_buffer(41384) := X"24430004";
        ram_buffer(41385) := X"AFC301F4";
        ram_buffer(41386) := X"8C420000";
        ram_buffer(41387) := X"8FC30030";
        ram_buffer(41388) := X"00000000";
        ram_buffer(41389) := X"00031C00";
        ram_buffer(41390) := X"00031C03";
        ram_buffer(41391) := X"A4430000";
        ram_buffer(41392) := X"10000872";
        ram_buffer(41393) := X"00000000";
        ram_buffer(41394) := X"32420200";
        ram_buffer(41395) := X"1040000D";
        ram_buffer(41396) := X"00000000";
        ram_buffer(41397) := X"8FC201F4";
        ram_buffer(41398) := X"00000000";
        ram_buffer(41399) := X"24430004";
        ram_buffer(41400) := X"AFC301F4";
        ram_buffer(41401) := X"8C420000";
        ram_buffer(41402) := X"8FC30030";
        ram_buffer(41403) := X"00000000";
        ram_buffer(41404) := X"00031E00";
        ram_buffer(41405) := X"00031E03";
        ram_buffer(41406) := X"A0430000";
        ram_buffer(41407) := X"10000863";
        ram_buffer(41408) := X"00000000";
        ram_buffer(41409) := X"8FC201F4";
        ram_buffer(41410) := X"00000000";
        ram_buffer(41411) := X"24430004";
        ram_buffer(41412) := X"AFC301F4";
        ram_buffer(41413) := X"8C420000";
        ram_buffer(41414) := X"8FC30030";
        ram_buffer(41415) := X"00000000";
        ram_buffer(41416) := X"AC430000";
        ram_buffer(41417) := X"10000859";
        ram_buffer(41418) := X"00000000";
        ram_buffer(41419) := X"36520010";
        ram_buffer(41420) := X"32420020";
        ram_buffer(41421) := X"1040000C";
        ram_buffer(41422) := X"00000000";
        ram_buffer(41423) := X"8FC201F4";
        ram_buffer(41424) := X"00000000";
        ram_buffer(41425) := X"24430007";
        ram_buffer(41426) := X"2402FFF8";
        ram_buffer(41427) := X"00621024";
        ram_buffer(41428) := X"24430008";
        ram_buffer(41429) := X"AFC301F4";
        ram_buffer(41430) := X"8C570004";
        ram_buffer(41431) := X"8C560000";
        ram_buffer(41432) := X"1000003C";
        ram_buffer(41433) := X"00000000";
        ram_buffer(41434) := X"32420010";
        ram_buffer(41435) := X"1040000B";
        ram_buffer(41436) := X"00000000";
        ram_buffer(41437) := X"8FC301F4";
        ram_buffer(41438) := X"00000000";
        ram_buffer(41439) := X"24620004";
        ram_buffer(41440) := X"AFC201F4";
        ram_buffer(41441) := X"8C620000";
        ram_buffer(41442) := X"00000000";
        ram_buffer(41443) := X"0040B821";
        ram_buffer(41444) := X"0000B021";
        ram_buffer(41445) := X"1000002F";
        ram_buffer(41446) := X"00000000";
        ram_buffer(41447) := X"32420040";
        ram_buffer(41448) := X"10400011";
        ram_buffer(41449) := X"00000000";
        ram_buffer(41450) := X"8FC301F4";
        ram_buffer(41451) := X"00000000";
        ram_buffer(41452) := X"24620004";
        ram_buffer(41453) := X"AFC201F4";
        ram_buffer(41454) := X"8C620000";
        ram_buffer(41455) := X"00000000";
        ram_buffer(41456) := X"AFC20194";
        ram_buffer(41457) := X"AFC00190";
        ram_buffer(41458) := X"8FC30194";
        ram_buffer(41459) := X"8FC20190";
        ram_buffer(41460) := X"00000000";
        ram_buffer(41461) := X"00402021";
        ram_buffer(41462) := X"30960000";
        ram_buffer(41463) := X"3077FFFF";
        ram_buffer(41464) := X"1000001C";
        ram_buffer(41465) := X"00000000";
        ram_buffer(41466) := X"32420200";
        ram_buffer(41467) := X"10400011";
        ram_buffer(41468) := X"00000000";
        ram_buffer(41469) := X"8FC301F4";
        ram_buffer(41470) := X"00000000";
        ram_buffer(41471) := X"24620004";
        ram_buffer(41472) := X"AFC201F4";
        ram_buffer(41473) := X"8C620000";
        ram_buffer(41474) := X"00000000";
        ram_buffer(41475) := X"AFC2019C";
        ram_buffer(41476) := X"AFC00198";
        ram_buffer(41477) := X"8FC3019C";
        ram_buffer(41478) := X"8FC20198";
        ram_buffer(41479) := X"00000000";
        ram_buffer(41480) := X"00402021";
        ram_buffer(41481) := X"30960000";
        ram_buffer(41482) := X"307700FF";
        ram_buffer(41483) := X"10000009";
        ram_buffer(41484) := X"00000000";
        ram_buffer(41485) := X"8FC301F4";
        ram_buffer(41486) := X"00000000";
        ram_buffer(41487) := X"24620004";
        ram_buffer(41488) := X"AFC201F4";
        ram_buffer(41489) := X"8C620000";
        ram_buffer(41490) := X"00000000";
        ram_buffer(41491) := X"0040B821";
        ram_buffer(41492) := X"0000B021";
        ram_buffer(41493) := X"AFD7005C";
        ram_buffer(41494) := X"AFD60058";
        ram_buffer(41495) := X"A3C00060";
        ram_buffer(41496) := X"2402FBFF";
        ram_buffer(41497) := X"02429024";
        ram_buffer(41498) := X"10000111";
        ram_buffer(41499) := X"00000000";
        ram_buffer(41500) := X"8FC201F4";
        ram_buffer(41501) := X"00000000";
        ram_buffer(41502) := X"24430004";
        ram_buffer(41503) := X"AFC301F4";
        ram_buffer(41504) := X"8C420000";
        ram_buffer(41505) := X"00000000";
        ram_buffer(41506) := X"AFC2005C";
        ram_buffer(41507) := X"AFC00058";
        ram_buffer(41508) := X"24020002";
        ram_buffer(41509) := X"A3C20060";
        ram_buffer(41510) := X"3C02100D";
        ram_buffer(41511) := X"2442A714";
        ram_buffer(41512) := X"AFC20070";
        ram_buffer(41513) := X"36520002";
        ram_buffer(41514) := X"24020030";
        ram_buffer(41515) := X"A3C20168";
        ram_buffer(41516) := X"24140078";
        ram_buffer(41517) := X"24020078";
        ram_buffer(41518) := X"A3C20169";
        ram_buffer(41519) := X"100000FC";
        ram_buffer(41520) := X"00000000";
        ram_buffer(41521) := X"8FC301F4";
        ram_buffer(41522) := X"00000000";
        ram_buffer(41523) := X"24620004";
        ram_buffer(41524) := X"AFC201F4";
        ram_buffer(41525) := X"8C730000";
        ram_buffer(41526) := X"A3C0009C";
        ram_buffer(41527) := X"1660000D";
        ram_buffer(41528) := X"00000000";
        ram_buffer(41529) := X"3C02100D";
        ram_buffer(41530) := X"2453A728";
        ram_buffer(41531) := X"8FC20038";
        ram_buffer(41532) := X"00000000";
        ram_buffer(41533) := X"00401821";
        ram_buffer(41534) := X"2C620007";
        ram_buffer(41535) := X"14400002";
        ram_buffer(41536) := X"00000000";
        ram_buffer(41537) := X"24030006";
        ram_buffer(41538) := X"AFC3006C";
        ram_buffer(41539) := X"100001E8";
        ram_buffer(41540) := X"00000000";
        ram_buffer(41541) := X"8FC20038";
        ram_buffer(41542) := X"00000000";
        ram_buffer(41543) := X"04400018";
        ram_buffer(41544) := X"00000000";
        ram_buffer(41545) := X"8FC20038";
        ram_buffer(41546) := X"00000000";
        ram_buffer(41547) := X"00403021";
        ram_buffer(41548) := X"00002821";
        ram_buffer(41549) := X"02602021";
        ram_buffer(41550) := X"0C02BC51";
        ram_buffer(41551) := X"00000000";
        ram_buffer(41552) := X"AFC20094";
        ram_buffer(41553) := X"8FC20094";
        ram_buffer(41554) := X"00000000";
        ram_buffer(41555) := X"10400007";
        ram_buffer(41556) := X"00000000";
        ram_buffer(41557) := X"8FC30094";
        ram_buffer(41558) := X"02601021";
        ram_buffer(41559) := X"00621023";
        ram_buffer(41560) := X"AFC2006C";
        ram_buffer(41561) := X"100001D2";
        ram_buffer(41562) := X"00000000";
        ram_buffer(41563) := X"8FC20038";
        ram_buffer(41564) := X"00000000";
        ram_buffer(41565) := X"AFC2006C";
        ram_buffer(41566) := X"100001CD";
        ram_buffer(41567) := X"00000000";
        ram_buffer(41568) := X"02602021";
        ram_buffer(41569) := X"0C02851E";
        ram_buffer(41570) := X"00000000";
        ram_buffer(41571) := X"AFC2006C";
        ram_buffer(41572) := X"100001C7";
        ram_buffer(41573) := X"00000000";
        ram_buffer(41574) := X"36520010";
        ram_buffer(41575) := X"32420020";
        ram_buffer(41576) := X"1040000E";
        ram_buffer(41577) := X"00000000";
        ram_buffer(41578) := X"8FC201F4";
        ram_buffer(41579) := X"00000000";
        ram_buffer(41580) := X"24430007";
        ram_buffer(41581) := X"2402FFF8";
        ram_buffer(41582) := X"00621024";
        ram_buffer(41583) := X"24430008";
        ram_buffer(41584) := X"AFC301F4";
        ram_buffer(41585) := X"8C430004";
        ram_buffer(41586) := X"8C420000";
        ram_buffer(41587) := X"AFC3017C";
        ram_buffer(41588) := X"AFC20178";
        ram_buffer(41589) := X"10000040";
        ram_buffer(41590) := X"00000000";
        ram_buffer(41591) := X"32420010";
        ram_buffer(41592) := X"1040000B";
        ram_buffer(41593) := X"00000000";
        ram_buffer(41594) := X"8FC301F4";
        ram_buffer(41595) := X"00000000";
        ram_buffer(41596) := X"24620004";
        ram_buffer(41597) := X"AFC201F4";
        ram_buffer(41598) := X"8C620000";
        ram_buffer(41599) := X"00000000";
        ram_buffer(41600) := X"AFC2017C";
        ram_buffer(41601) := X"AFC00178";
        ram_buffer(41602) := X"10000033";
        ram_buffer(41603) := X"00000000";
        ram_buffer(41604) := X"32420040";
        ram_buffer(41605) := X"10400013";
        ram_buffer(41606) := X"00000000";
        ram_buffer(41607) := X"8FC301F4";
        ram_buffer(41608) := X"00000000";
        ram_buffer(41609) := X"24620004";
        ram_buffer(41610) := X"AFC201F4";
        ram_buffer(41611) := X"8C620000";
        ram_buffer(41612) := X"00000000";
        ram_buffer(41613) := X"AFC201A4";
        ram_buffer(41614) := X"AFC001A0";
        ram_buffer(41615) := X"8FC301A4";
        ram_buffer(41616) := X"8FC201A0";
        ram_buffer(41617) := X"00000000";
        ram_buffer(41618) := X"00402021";
        ram_buffer(41619) := X"30840000";
        ram_buffer(41620) := X"AFC40178";
        ram_buffer(41621) := X"3062FFFF";
        ram_buffer(41622) := X"AFC2017C";
        ram_buffer(41623) := X"1000001E";
        ram_buffer(41624) := X"00000000";
        ram_buffer(41625) := X"32420200";
        ram_buffer(41626) := X"10400013";
        ram_buffer(41627) := X"00000000";
        ram_buffer(41628) := X"8FC301F4";
        ram_buffer(41629) := X"00000000";
        ram_buffer(41630) := X"24620004";
        ram_buffer(41631) := X"AFC201F4";
        ram_buffer(41632) := X"8C620000";
        ram_buffer(41633) := X"00000000";
        ram_buffer(41634) := X"AFC201AC";
        ram_buffer(41635) := X"AFC001A8";
        ram_buffer(41636) := X"8FC301AC";
        ram_buffer(41637) := X"8FC201A8";
        ram_buffer(41638) := X"00000000";
        ram_buffer(41639) := X"00402021";
        ram_buffer(41640) := X"30840000";
        ram_buffer(41641) := X"AFC40178";
        ram_buffer(41642) := X"306200FF";
        ram_buffer(41643) := X"AFC2017C";
        ram_buffer(41644) := X"10000009";
        ram_buffer(41645) := X"00000000";
        ram_buffer(41646) := X"8FC301F4";
        ram_buffer(41647) := X"00000000";
        ram_buffer(41648) := X"24620004";
        ram_buffer(41649) := X"AFC201F4";
        ram_buffer(41650) := X"8C620000";
        ram_buffer(41651) := X"00000000";
        ram_buffer(41652) := X"AFC2017C";
        ram_buffer(41653) := X"AFC00178";
        ram_buffer(41654) := X"8FC3017C";
        ram_buffer(41655) := X"8FC20178";
        ram_buffer(41656) := X"AFC3005C";
        ram_buffer(41657) := X"AFC20058";
        ram_buffer(41658) := X"24020001";
        ram_buffer(41659) := X"A3C20060";
        ram_buffer(41660) := X"1000006F";
        ram_buffer(41661) := X"00000000";
        ram_buffer(41662) := X"3C02100D";
        ram_buffer(41663) := X"2442A730";
        ram_buffer(41664) := X"AFC20070";
        ram_buffer(41665) := X"10000004";
        ram_buffer(41666) := X"00000000";
        ram_buffer(41667) := X"3C02100D";
        ram_buffer(41668) := X"2442A714";
        ram_buffer(41669) := X"AFC20070";
        ram_buffer(41670) := X"32420020";
        ram_buffer(41671) := X"1040000E";
        ram_buffer(41672) := X"00000000";
        ram_buffer(41673) := X"8FC201F4";
        ram_buffer(41674) := X"00000000";
        ram_buffer(41675) := X"24430007";
        ram_buffer(41676) := X"2402FFF8";
        ram_buffer(41677) := X"00621024";
        ram_buffer(41678) := X"24430008";
        ram_buffer(41679) := X"AFC301F4";
        ram_buffer(41680) := X"8C430004";
        ram_buffer(41681) := X"8C420000";
        ram_buffer(41682) := X"AFC30184";
        ram_buffer(41683) := X"AFC20180";
        ram_buffer(41684) := X"10000040";
        ram_buffer(41685) := X"00000000";
        ram_buffer(41686) := X"32420010";
        ram_buffer(41687) := X"1040000B";
        ram_buffer(41688) := X"00000000";
        ram_buffer(41689) := X"8FC301F4";
        ram_buffer(41690) := X"00000000";
        ram_buffer(41691) := X"24620004";
        ram_buffer(41692) := X"AFC201F4";
        ram_buffer(41693) := X"8C620000";
        ram_buffer(41694) := X"00000000";
        ram_buffer(41695) := X"AFC20184";
        ram_buffer(41696) := X"AFC00180";
        ram_buffer(41697) := X"10000033";
        ram_buffer(41698) := X"00000000";
        ram_buffer(41699) := X"32420040";
        ram_buffer(41700) := X"10400013";
        ram_buffer(41701) := X"00000000";
        ram_buffer(41702) := X"8FC301F4";
        ram_buffer(41703) := X"00000000";
        ram_buffer(41704) := X"24620004";
        ram_buffer(41705) := X"AFC201F4";
        ram_buffer(41706) := X"8C620000";
        ram_buffer(41707) := X"00000000";
        ram_buffer(41708) := X"AFC201B4";
        ram_buffer(41709) := X"AFC001B0";
        ram_buffer(41710) := X"8FC301B4";
        ram_buffer(41711) := X"8FC201B0";
        ram_buffer(41712) := X"00000000";
        ram_buffer(41713) := X"00402021";
        ram_buffer(41714) := X"30840000";
        ram_buffer(41715) := X"AFC40180";
        ram_buffer(41716) := X"3062FFFF";
        ram_buffer(41717) := X"AFC20184";
        ram_buffer(41718) := X"1000001E";
        ram_buffer(41719) := X"00000000";
        ram_buffer(41720) := X"32420200";
        ram_buffer(41721) := X"10400013";
        ram_buffer(41722) := X"00000000";
        ram_buffer(41723) := X"8FC301F4";
        ram_buffer(41724) := X"00000000";
        ram_buffer(41725) := X"24620004";
        ram_buffer(41726) := X"AFC201F4";
        ram_buffer(41727) := X"8C620000";
        ram_buffer(41728) := X"00000000";
        ram_buffer(41729) := X"AFC201BC";
        ram_buffer(41730) := X"AFC001B8";
        ram_buffer(41731) := X"8FC301BC";
        ram_buffer(41732) := X"8FC201B8";
        ram_buffer(41733) := X"00000000";
        ram_buffer(41734) := X"00402021";
        ram_buffer(41735) := X"30840000";
        ram_buffer(41736) := X"AFC40180";
        ram_buffer(41737) := X"306200FF";
        ram_buffer(41738) := X"AFC20184";
        ram_buffer(41739) := X"10000009";
        ram_buffer(41740) := X"00000000";
        ram_buffer(41741) := X"8FC301F4";
        ram_buffer(41742) := X"00000000";
        ram_buffer(41743) := X"24620004";
        ram_buffer(41744) := X"AFC201F4";
        ram_buffer(41745) := X"8C620000";
        ram_buffer(41746) := X"00000000";
        ram_buffer(41747) := X"AFC20184";
        ram_buffer(41748) := X"AFC00180";
        ram_buffer(41749) := X"8FC30184";
        ram_buffer(41750) := X"8FC20180";
        ram_buffer(41751) := X"AFC3005C";
        ram_buffer(41752) := X"AFC20058";
        ram_buffer(41753) := X"24020002";
        ram_buffer(41754) := X"A3C20060";
        ram_buffer(41755) := X"32420001";
        ram_buffer(41756) := X"1040000D";
        ram_buffer(41757) := X"00000000";
        ram_buffer(41758) := X"8FC20058";
        ram_buffer(41759) := X"8FC3005C";
        ram_buffer(41760) := X"00000000";
        ram_buffer(41761) := X"00431025";
        ram_buffer(41762) := X"10400007";
        ram_buffer(41763) := X"00000000";
        ram_buffer(41764) := X"24020030";
        ram_buffer(41765) := X"A3C20168";
        ram_buffer(41766) := X"00141600";
        ram_buffer(41767) := X"00021603";
        ram_buffer(41768) := X"A3C20169";
        ram_buffer(41769) := X"36520002";
        ram_buffer(41770) := X"2402FBFF";
        ram_buffer(41771) := X"02429024";
        ram_buffer(41772) := X"A3C0009C";
        ram_buffer(41773) := X"8FC20038";
        ram_buffer(41774) := X"00000000";
        ram_buffer(41775) := X"AFC20064";
        ram_buffer(41776) := X"8FC20064";
        ram_buffer(41777) := X"00000000";
        ram_buffer(41778) := X"04400003";
        ram_buffer(41779) := X"00000000";
        ram_buffer(41780) := X"2402FF7F";
        ram_buffer(41781) := X"02429024";
        ram_buffer(41782) := X"27D30104";
        ram_buffer(41783) := X"26730064";
        ram_buffer(41784) := X"8FC30058";
        ram_buffer(41785) := X"8FC2005C";
        ram_buffer(41786) := X"00000000";
        ram_buffer(41787) := X"00621825";
        ram_buffer(41788) := X"14600005";
        ram_buffer(41789) := X"00000000";
        ram_buffer(41790) := X"8FC20038";
        ram_buffer(41791) := X"00000000";
        ram_buffer(41792) := X"104000CD";
        ram_buffer(41793) := X"00000000";
        ram_buffer(41794) := X"93C30060";
        ram_buffer(41795) := X"24020001";
        ram_buffer(41796) := X"1062002E";
        ram_buffer(41797) := X"00000000";
        ram_buffer(41798) := X"24020002";
        ram_buffer(41799) := X"1062009C";
        ram_buffer(41800) := X"00000000";
        ram_buffer(41801) := X"146000B8";
        ram_buffer(41802) := X"00000000";
        ram_buffer(41803) := X"2673FFFF";
        ram_buffer(41804) := X"93C2005F";
        ram_buffer(41805) := X"00000000";
        ram_buffer(41806) := X"30420007";
        ram_buffer(41807) := X"304200FF";
        ram_buffer(41808) := X"24420030";
        ram_buffer(41809) := X"304200FF";
        ram_buffer(41810) := X"00021600";
        ram_buffer(41811) := X"00021603";
        ram_buffer(41812) := X"A2620000";
        ram_buffer(41813) := X"8FC20058";
        ram_buffer(41814) := X"00000000";
        ram_buffer(41815) := X"00021F40";
        ram_buffer(41816) := X"8FC2005C";
        ram_buffer(41817) := X"00000000";
        ram_buffer(41818) := X"000210C2";
        ram_buffer(41819) := X"00431025";
        ram_buffer(41820) := X"AFC2005C";
        ram_buffer(41821) := X"8FC20058";
        ram_buffer(41822) := X"00000000";
        ram_buffer(41823) := X"000210C2";
        ram_buffer(41824) := X"AFC20058";
        ram_buffer(41825) := X"8FC30058";
        ram_buffer(41826) := X"8FC2005C";
        ram_buffer(41827) := X"00000000";
        ram_buffer(41828) := X"00621825";
        ram_buffer(41829) := X"1460FFE5";
        ram_buffer(41830) := X"00000000";
        ram_buffer(41831) := X"32420001";
        ram_buffer(41832) := X"104000A2";
        ram_buffer(41833) := X"00000000";
        ram_buffer(41834) := X"82630000";
        ram_buffer(41835) := X"24020030";
        ram_buffer(41836) := X"1062009E";
        ram_buffer(41837) := X"00000000";
        ram_buffer(41838) := X"2673FFFF";
        ram_buffer(41839) := X"24020030";
        ram_buffer(41840) := X"A2620000";
        ram_buffer(41841) := X"10000099";
        ram_buffer(41842) := X"00000000";
        ram_buffer(41843) := X"8FC20058";
        ram_buffer(41844) := X"00000000";
        ram_buffer(41845) := X"14400014";
        ram_buffer(41846) := X"00000000";
        ram_buffer(41847) := X"8FC20058";
        ram_buffer(41848) := X"00000000";
        ram_buffer(41849) := X"14400006";
        ram_buffer(41850) := X"00000000";
        ram_buffer(41851) := X"8FC2005C";
        ram_buffer(41852) := X"00000000";
        ram_buffer(41853) := X"2C42000A";
        ram_buffer(41854) := X"1040000B";
        ram_buffer(41855) := X"00000000";
        ram_buffer(41856) := X"2673FFFF";
        ram_buffer(41857) := X"93C2005F";
        ram_buffer(41858) := X"00000000";
        ram_buffer(41859) := X"24420030";
        ram_buffer(41860) := X"304200FF";
        ram_buffer(41861) := X"00021600";
        ram_buffer(41862) := X"00021603";
        ram_buffer(41863) := X"A2620000";
        ram_buffer(41864) := X"10000083";
        ram_buffer(41865) := X"00000000";
        ram_buffer(41866) := X"AFC000B4";
        ram_buffer(41867) := X"2673FFFF";
        ram_buffer(41868) := X"8FC3005C";
        ram_buffer(41869) := X"8FC20058";
        ram_buffer(41870) := X"2407000A";
        ram_buffer(41871) := X"00003021";
        ram_buffer(41872) := X"00602821";
        ram_buffer(41873) := X"00402021";
        ram_buffer(41874) := X"0C030BFE";
        ram_buffer(41875) := X"00000000";
        ram_buffer(41876) := X"306200FF";
        ram_buffer(41877) := X"24420030";
        ram_buffer(41878) := X"304200FF";
        ram_buffer(41879) := X"00021600";
        ram_buffer(41880) := X"00021603";
        ram_buffer(41881) := X"A2620000";
        ram_buffer(41882) := X"8FC200B4";
        ram_buffer(41883) := X"00000000";
        ram_buffer(41884) := X"24420001";
        ram_buffer(41885) := X"AFC200B4";
        ram_buffer(41886) := X"32420400";
        ram_buffer(41887) := X"10400032";
        ram_buffer(41888) := X"00000000";
        ram_buffer(41889) := X"8FC20044";
        ram_buffer(41890) := X"00000000";
        ram_buffer(41891) := X"80420000";
        ram_buffer(41892) := X"00000000";
        ram_buffer(41893) := X"00401821";
        ram_buffer(41894) := X"8FC200B4";
        ram_buffer(41895) := X"00000000";
        ram_buffer(41896) := X"14620029";
        ram_buffer(41897) := X"00000000";
        ram_buffer(41898) := X"8FC20044";
        ram_buffer(41899) := X"00000000";
        ram_buffer(41900) := X"80430000";
        ram_buffer(41901) := X"2402007F";
        ram_buffer(41902) := X"10620023";
        ram_buffer(41903) := X"00000000";
        ram_buffer(41904) := X"8FC20058";
        ram_buffer(41905) := X"00000000";
        ram_buffer(41906) := X"1440000A";
        ram_buffer(41907) := X"00000000";
        ram_buffer(41908) := X"8FC20058";
        ram_buffer(41909) := X"00000000";
        ram_buffer(41910) := X"1440001B";
        ram_buffer(41911) := X"00000000";
        ram_buffer(41912) := X"8FC2005C";
        ram_buffer(41913) := X"00000000";
        ram_buffer(41914) := X"2C42000A";
        ram_buffer(41915) := X"14400016";
        ram_buffer(41916) := X"00000000";
        ram_buffer(41917) := X"8FC20040";
        ram_buffer(41918) := X"00000000";
        ram_buffer(41919) := X"00021023";
        ram_buffer(41920) := X"02629821";
        ram_buffer(41921) := X"8FC60040";
        ram_buffer(41922) := X"8FC5003C";
        ram_buffer(41923) := X"02602021";
        ram_buffer(41924) := X"0C02CCBF";
        ram_buffer(41925) := X"00000000";
        ram_buffer(41926) := X"AFC000B4";
        ram_buffer(41927) := X"8FC20044";
        ram_buffer(41928) := X"00000000";
        ram_buffer(41929) := X"24420001";
        ram_buffer(41930) := X"80420000";
        ram_buffer(41931) := X"00000000";
        ram_buffer(41932) := X"10400005";
        ram_buffer(41933) := X"00000000";
        ram_buffer(41934) := X"8FC20044";
        ram_buffer(41935) := X"00000000";
        ram_buffer(41936) := X"24420001";
        ram_buffer(41937) := X"AFC20044";
        ram_buffer(41938) := X"8FC3005C";
        ram_buffer(41939) := X"8FC20058";
        ram_buffer(41940) := X"2407000A";
        ram_buffer(41941) := X"00003021";
        ram_buffer(41942) := X"00602821";
        ram_buffer(41943) := X"00402021";
        ram_buffer(41944) := X"0C030A67";
        ram_buffer(41945) := X"00000000";
        ram_buffer(41946) := X"AFC3005C";
        ram_buffer(41947) := X"AFC20058";
        ram_buffer(41948) := X"8FC30058";
        ram_buffer(41949) := X"8FC2005C";
        ram_buffer(41950) := X"00000000";
        ram_buffer(41951) := X"00621825";
        ram_buffer(41952) := X"1460FFAA";
        ram_buffer(41953) := X"00000000";
        ram_buffer(41954) := X"10000029";
        ram_buffer(41955) := X"00000000";
        ram_buffer(41956) := X"2673FFFF";
        ram_buffer(41957) := X"8FC2005C";
        ram_buffer(41958) := X"00000000";
        ram_buffer(41959) := X"3043000F";
        ram_buffer(41960) := X"8FC20070";
        ram_buffer(41961) := X"00000000";
        ram_buffer(41962) := X"00431021";
        ram_buffer(41963) := X"80420000";
        ram_buffer(41964) := X"00000000";
        ram_buffer(41965) := X"A2620000";
        ram_buffer(41966) := X"8FC20058";
        ram_buffer(41967) := X"00000000";
        ram_buffer(41968) := X"00021F00";
        ram_buffer(41969) := X"8FC2005C";
        ram_buffer(41970) := X"00000000";
        ram_buffer(41971) := X"00021102";
        ram_buffer(41972) := X"00431025";
        ram_buffer(41973) := X"AFC2005C";
        ram_buffer(41974) := X"8FC20058";
        ram_buffer(41975) := X"00000000";
        ram_buffer(41976) := X"00021102";
        ram_buffer(41977) := X"AFC20058";
        ram_buffer(41978) := X"8FC30058";
        ram_buffer(41979) := X"8FC2005C";
        ram_buffer(41980) := X"00000000";
        ram_buffer(41981) := X"00621825";
        ram_buffer(41982) := X"1460FFE5";
        ram_buffer(41983) := X"00000000";
        ram_buffer(41984) := X"1000000B";
        ram_buffer(41985) := X"00000000";
        ram_buffer(41986) := X"3C02100D";
        ram_buffer(41987) := X"2453A744";
        ram_buffer(41988) := X"02602021";
        ram_buffer(41989) := X"0C02851E";
        ram_buffer(41990) := X"00000000";
        ram_buffer(41991) := X"AFC2006C";
        ram_buffer(41992) := X"00000000";
        ram_buffer(41993) := X"10000022";
        ram_buffer(41994) := X"00000000";
        ram_buffer(41995) := X"00000000";
        ram_buffer(41996) := X"1000000B";
        ram_buffer(41997) := X"00000000";
        ram_buffer(41998) := X"93C20060";
        ram_buffer(41999) := X"00000000";
        ram_buffer(42000) := X"14400007";
        ram_buffer(42001) := X"00000000";
        ram_buffer(42002) := X"32420001";
        ram_buffer(42003) := X"10400004";
        ram_buffer(42004) := X"00000000";
        ram_buffer(42005) := X"2673FFFF";
        ram_buffer(42006) := X"24020030";
        ram_buffer(42007) := X"A2620000";
        ram_buffer(42008) := X"27C20104";
        ram_buffer(42009) := X"24420064";
        ram_buffer(42010) := X"00401821";
        ram_buffer(42011) := X"02601021";
        ram_buffer(42012) := X"00621023";
        ram_buffer(42013) := X"AFC2006C";
        ram_buffer(42014) := X"1000000D";
        ram_buffer(42015) := X"00000000";
        ram_buffer(42016) := X"12800607";
        ram_buffer(42017) := X"00000000";
        ram_buffer(42018) := X"27D30104";
        ram_buffer(42019) := X"00141600";
        ram_buffer(42020) := X"00021603";
        ram_buffer(42021) := X"A2620000";
        ram_buffer(42022) := X"24020001";
        ram_buffer(42023) := X"AFC2006C";
        ram_buffer(42024) := X"A3C0009C";
        ram_buffer(42025) := X"10000002";
        ram_buffer(42026) := X"00000000";
        ram_buffer(42027) := X"00000000";
        ram_buffer(42028) := X"8FC40064";
        ram_buffer(42029) := X"8FC3006C";
        ram_buffer(42030) := X"00000000";
        ram_buffer(42031) := X"0064102A";
        ram_buffer(42032) := X"10400002";
        ram_buffer(42033) := X"00000000";
        ram_buffer(42034) := X"00801821";
        ram_buffer(42035) := X"AFC30068";
        ram_buffer(42036) := X"83C2009C";
        ram_buffer(42037) := X"00000000";
        ram_buffer(42038) := X"10400005";
        ram_buffer(42039) := X"00000000";
        ram_buffer(42040) := X"8FC20068";
        ram_buffer(42041) := X"00000000";
        ram_buffer(42042) := X"24420001";
        ram_buffer(42043) := X"AFC20068";
        ram_buffer(42044) := X"32420002";
        ram_buffer(42045) := X"10400005";
        ram_buffer(42046) := X"00000000";
        ram_buffer(42047) := X"8FC20068";
        ram_buffer(42048) := X"00000000";
        ram_buffer(42049) := X"24420002";
        ram_buffer(42050) := X"AFC20068";
        ram_buffer(42051) := X"32420084";
        ram_buffer(42052) := X"14400045";
        ram_buffer(42053) := X"00000000";
        ram_buffer(42054) := X"8FC30034";
        ram_buffer(42055) := X"8FC20068";
        ram_buffer(42056) := X"00000000";
        ram_buffer(42057) := X"00628823";
        ram_buffer(42058) := X"1A20003F";
        ram_buffer(42059) := X"00000000";
        ram_buffer(42060) := X"1000001E";
        ram_buffer(42061) := X"00000000";
        ram_buffer(42062) := X"3C02100D";
        ram_buffer(42063) := X"2442A8D0";
        ram_buffer(42064) := X"AE020000";
        ram_buffer(42065) := X"24020010";
        ram_buffer(42066) := X"AE020004";
        ram_buffer(42067) := X"8FC200C0";
        ram_buffer(42068) := X"00000000";
        ram_buffer(42069) := X"24420010";
        ram_buffer(42070) := X"AFC200C0";
        ram_buffer(42071) := X"26100008";
        ram_buffer(42072) := X"8FC200BC";
        ram_buffer(42073) := X"00000000";
        ram_buffer(42074) := X"24420001";
        ram_buffer(42075) := X"AFC200BC";
        ram_buffer(42076) := X"8FC200BC";
        ram_buffer(42077) := X"00000000";
        ram_buffer(42078) := X"28420008";
        ram_buffer(42079) := X"1440000A";
        ram_buffer(42080) := X"00000000";
        ram_buffer(42081) := X"27C200B8";
        ram_buffer(42082) := X"00403021";
        ram_buffer(42083) := X"8FC501EC";
        ram_buffer(42084) := X"8FC401E8";
        ram_buffer(42085) := X"0C02EAF5";
        ram_buffer(42086) := X"00000000";
        ram_buffer(42087) := X"144005D4";
        ram_buffer(42088) := X"00000000";
        ram_buffer(42089) := X"27D000C4";
        ram_buffer(42090) := X"2631FFF0";
        ram_buffer(42091) := X"2A220011";
        ram_buffer(42092) := X"1040FFE1";
        ram_buffer(42093) := X"00000000";
        ram_buffer(42094) := X"3C02100D";
        ram_buffer(42095) := X"2442A8D0";
        ram_buffer(42096) := X"AE020000";
        ram_buffer(42097) := X"02201021";
        ram_buffer(42098) := X"AE020004";
        ram_buffer(42099) := X"8FC300C0";
        ram_buffer(42100) := X"02201021";
        ram_buffer(42101) := X"00621021";
        ram_buffer(42102) := X"AFC200C0";
        ram_buffer(42103) := X"26100008";
        ram_buffer(42104) := X"8FC200BC";
        ram_buffer(42105) := X"00000000";
        ram_buffer(42106) := X"24420001";
        ram_buffer(42107) := X"AFC200BC";
        ram_buffer(42108) := X"8FC200BC";
        ram_buffer(42109) := X"00000000";
        ram_buffer(42110) := X"28420008";
        ram_buffer(42111) := X"1440000A";
        ram_buffer(42112) := X"00000000";
        ram_buffer(42113) := X"27C200B8";
        ram_buffer(42114) := X"00403021";
        ram_buffer(42115) := X"8FC501EC";
        ram_buffer(42116) := X"8FC401E8";
        ram_buffer(42117) := X"0C02EAF5";
        ram_buffer(42118) := X"00000000";
        ram_buffer(42119) := X"144005B7";
        ram_buffer(42120) := X"00000000";
        ram_buffer(42121) := X"27D000C4";
        ram_buffer(42122) := X"83C2009C";
        ram_buffer(42123) := X"00000000";
        ram_buffer(42124) := X"1040001C";
        ram_buffer(42125) := X"00000000";
        ram_buffer(42126) := X"27C2009C";
        ram_buffer(42127) := X"AE020000";
        ram_buffer(42128) := X"24020001";
        ram_buffer(42129) := X"AE020004";
        ram_buffer(42130) := X"8FC200C0";
        ram_buffer(42131) := X"00000000";
        ram_buffer(42132) := X"24420001";
        ram_buffer(42133) := X"AFC200C0";
        ram_buffer(42134) := X"26100008";
        ram_buffer(42135) := X"8FC200BC";
        ram_buffer(42136) := X"00000000";
        ram_buffer(42137) := X"24420001";
        ram_buffer(42138) := X"AFC200BC";
        ram_buffer(42139) := X"8FC200BC";
        ram_buffer(42140) := X"00000000";
        ram_buffer(42141) := X"28420008";
        ram_buffer(42142) := X"1440000A";
        ram_buffer(42143) := X"00000000";
        ram_buffer(42144) := X"27C200B8";
        ram_buffer(42145) := X"00403021";
        ram_buffer(42146) := X"8FC501EC";
        ram_buffer(42147) := X"8FC401E8";
        ram_buffer(42148) := X"0C02EAF5";
        ram_buffer(42149) := X"00000000";
        ram_buffer(42150) := X"1440059B";
        ram_buffer(42151) := X"00000000";
        ram_buffer(42152) := X"27D000C4";
        ram_buffer(42153) := X"32420002";
        ram_buffer(42154) := X"1040001C";
        ram_buffer(42155) := X"00000000";
        ram_buffer(42156) := X"27C20168";
        ram_buffer(42157) := X"AE020000";
        ram_buffer(42158) := X"24020002";
        ram_buffer(42159) := X"AE020004";
        ram_buffer(42160) := X"8FC200C0";
        ram_buffer(42161) := X"00000000";
        ram_buffer(42162) := X"24420002";
        ram_buffer(42163) := X"AFC200C0";
        ram_buffer(42164) := X"26100008";
        ram_buffer(42165) := X"8FC200BC";
        ram_buffer(42166) := X"00000000";
        ram_buffer(42167) := X"24420001";
        ram_buffer(42168) := X"AFC200BC";
        ram_buffer(42169) := X"8FC200BC";
        ram_buffer(42170) := X"00000000";
        ram_buffer(42171) := X"28420008";
        ram_buffer(42172) := X"1440000A";
        ram_buffer(42173) := X"00000000";
        ram_buffer(42174) := X"27C200B8";
        ram_buffer(42175) := X"00403021";
        ram_buffer(42176) := X"8FC501EC";
        ram_buffer(42177) := X"8FC401E8";
        ram_buffer(42178) := X"0C02EAF5";
        ram_buffer(42179) := X"00000000";
        ram_buffer(42180) := X"14400580";
        ram_buffer(42181) := X"00000000";
        ram_buffer(42182) := X"27D000C4";
        ram_buffer(42183) := X"32430084";
        ram_buffer(42184) := X"24020080";
        ram_buffer(42185) := X"14620045";
        ram_buffer(42186) := X"00000000";
        ram_buffer(42187) := X"8FC30034";
        ram_buffer(42188) := X"8FC20068";
        ram_buffer(42189) := X"00000000";
        ram_buffer(42190) := X"00628823";
        ram_buffer(42191) := X"1A20003F";
        ram_buffer(42192) := X"00000000";
        ram_buffer(42193) := X"1000001E";
        ram_buffer(42194) := X"00000000";
        ram_buffer(42195) := X"3C02100D";
        ram_buffer(42196) := X"2442A8E0";
        ram_buffer(42197) := X"AE020000";
        ram_buffer(42198) := X"24020010";
        ram_buffer(42199) := X"AE020004";
        ram_buffer(42200) := X"8FC200C0";
        ram_buffer(42201) := X"00000000";
        ram_buffer(42202) := X"24420010";
        ram_buffer(42203) := X"AFC200C0";
        ram_buffer(42204) := X"26100008";
        ram_buffer(42205) := X"8FC200BC";
        ram_buffer(42206) := X"00000000";
        ram_buffer(42207) := X"24420001";
        ram_buffer(42208) := X"AFC200BC";
        ram_buffer(42209) := X"8FC200BC";
        ram_buffer(42210) := X"00000000";
        ram_buffer(42211) := X"28420008";
        ram_buffer(42212) := X"1440000A";
        ram_buffer(42213) := X"00000000";
        ram_buffer(42214) := X"27C200B8";
        ram_buffer(42215) := X"00403021";
        ram_buffer(42216) := X"8FC501EC";
        ram_buffer(42217) := X"8FC401E8";
        ram_buffer(42218) := X"0C02EAF5";
        ram_buffer(42219) := X"00000000";
        ram_buffer(42220) := X"1440055B";
        ram_buffer(42221) := X"00000000";
        ram_buffer(42222) := X"27D000C4";
        ram_buffer(42223) := X"2631FFF0";
        ram_buffer(42224) := X"2A220011";
        ram_buffer(42225) := X"1040FFE1";
        ram_buffer(42226) := X"00000000";
        ram_buffer(42227) := X"3C02100D";
        ram_buffer(42228) := X"2442A8E0";
        ram_buffer(42229) := X"AE020000";
        ram_buffer(42230) := X"02201021";
        ram_buffer(42231) := X"AE020004";
        ram_buffer(42232) := X"8FC300C0";
        ram_buffer(42233) := X"02201021";
        ram_buffer(42234) := X"00621021";
        ram_buffer(42235) := X"AFC200C0";
        ram_buffer(42236) := X"26100008";
        ram_buffer(42237) := X"8FC200BC";
        ram_buffer(42238) := X"00000000";
        ram_buffer(42239) := X"24420001";
        ram_buffer(42240) := X"AFC200BC";
        ram_buffer(42241) := X"8FC200BC";
        ram_buffer(42242) := X"00000000";
        ram_buffer(42243) := X"28420008";
        ram_buffer(42244) := X"1440000A";
        ram_buffer(42245) := X"00000000";
        ram_buffer(42246) := X"27C200B8";
        ram_buffer(42247) := X"00403021";
        ram_buffer(42248) := X"8FC501EC";
        ram_buffer(42249) := X"8FC401E8";
        ram_buffer(42250) := X"0C02EAF5";
        ram_buffer(42251) := X"00000000";
        ram_buffer(42252) := X"1440053E";
        ram_buffer(42253) := X"00000000";
        ram_buffer(42254) := X"27D000C4";
        ram_buffer(42255) := X"8FC30064";
        ram_buffer(42256) := X"8FC2006C";
        ram_buffer(42257) := X"00000000";
        ram_buffer(42258) := X"00628823";
        ram_buffer(42259) := X"1A20003F";
        ram_buffer(42260) := X"00000000";
        ram_buffer(42261) := X"1000001E";
        ram_buffer(42262) := X"00000000";
        ram_buffer(42263) := X"3C02100D";
        ram_buffer(42264) := X"2442A8E0";
        ram_buffer(42265) := X"AE020000";
        ram_buffer(42266) := X"24020010";
        ram_buffer(42267) := X"AE020004";
        ram_buffer(42268) := X"8FC200C0";
        ram_buffer(42269) := X"00000000";
        ram_buffer(42270) := X"24420010";
        ram_buffer(42271) := X"AFC200C0";
        ram_buffer(42272) := X"26100008";
        ram_buffer(42273) := X"8FC200BC";
        ram_buffer(42274) := X"00000000";
        ram_buffer(42275) := X"24420001";
        ram_buffer(42276) := X"AFC200BC";
        ram_buffer(42277) := X"8FC200BC";
        ram_buffer(42278) := X"00000000";
        ram_buffer(42279) := X"28420008";
        ram_buffer(42280) := X"1440000A";
        ram_buffer(42281) := X"00000000";
        ram_buffer(42282) := X"27C200B8";
        ram_buffer(42283) := X"00403021";
        ram_buffer(42284) := X"8FC501EC";
        ram_buffer(42285) := X"8FC401E8";
        ram_buffer(42286) := X"0C02EAF5";
        ram_buffer(42287) := X"00000000";
        ram_buffer(42288) := X"1440051D";
        ram_buffer(42289) := X"00000000";
        ram_buffer(42290) := X"27D000C4";
        ram_buffer(42291) := X"2631FFF0";
        ram_buffer(42292) := X"2A220011";
        ram_buffer(42293) := X"1040FFE1";
        ram_buffer(42294) := X"00000000";
        ram_buffer(42295) := X"3C02100D";
        ram_buffer(42296) := X"2442A8E0";
        ram_buffer(42297) := X"AE020000";
        ram_buffer(42298) := X"02201021";
        ram_buffer(42299) := X"AE020004";
        ram_buffer(42300) := X"8FC300C0";
        ram_buffer(42301) := X"02201021";
        ram_buffer(42302) := X"00621021";
        ram_buffer(42303) := X"AFC200C0";
        ram_buffer(42304) := X"26100008";
        ram_buffer(42305) := X"8FC200BC";
        ram_buffer(42306) := X"00000000";
        ram_buffer(42307) := X"24420001";
        ram_buffer(42308) := X"AFC200BC";
        ram_buffer(42309) := X"8FC200BC";
        ram_buffer(42310) := X"00000000";
        ram_buffer(42311) := X"28420008";
        ram_buffer(42312) := X"1440000A";
        ram_buffer(42313) := X"00000000";
        ram_buffer(42314) := X"27C200B8";
        ram_buffer(42315) := X"00403021";
        ram_buffer(42316) := X"8FC501EC";
        ram_buffer(42317) := X"8FC401E8";
        ram_buffer(42318) := X"0C02EAF5";
        ram_buffer(42319) := X"00000000";
        ram_buffer(42320) := X"14400500";
        ram_buffer(42321) := X"00000000";
        ram_buffer(42322) := X"27D000C4";
        ram_buffer(42323) := X"32420100";
        ram_buffer(42324) := X"1440001F";
        ram_buffer(42325) := X"00000000";
        ram_buffer(42326) := X"AE130000";
        ram_buffer(42327) := X"8FC2006C";
        ram_buffer(42328) := X"00000000";
        ram_buffer(42329) := X"AE020004";
        ram_buffer(42330) := X"8FC300C0";
        ram_buffer(42331) := X"8FC2006C";
        ram_buffer(42332) := X"00000000";
        ram_buffer(42333) := X"00621021";
        ram_buffer(42334) := X"AFC200C0";
        ram_buffer(42335) := X"26100008";
        ram_buffer(42336) := X"8FC200BC";
        ram_buffer(42337) := X"00000000";
        ram_buffer(42338) := X"24420001";
        ram_buffer(42339) := X"AFC200BC";
        ram_buffer(42340) := X"8FC200BC";
        ram_buffer(42341) := X"00000000";
        ram_buffer(42342) := X"28420008";
        ram_buffer(42343) := X"14400452";
        ram_buffer(42344) := X"00000000";
        ram_buffer(42345) := X"27C200B8";
        ram_buffer(42346) := X"00403021";
        ram_buffer(42347) := X"8FC501EC";
        ram_buffer(42348) := X"8FC401E8";
        ram_buffer(42349) := X"0C02EAF5";
        ram_buffer(42350) := X"00000000";
        ram_buffer(42351) := X"144004E4";
        ram_buffer(42352) := X"00000000";
        ram_buffer(42353) := X"27D000C4";
        ram_buffer(42354) := X"10000447";
        ram_buffer(42355) := X"00000000";
        ram_buffer(42356) := X"2A820066";
        ram_buffer(42357) := X"1440035A";
        ram_buffer(42358) := X"00000000";
        ram_buffer(42359) := X"8FC300A4";
        ram_buffer(42360) := X"8FC200A0";
        ram_buffer(42361) := X"00003821";
        ram_buffer(42362) := X"00003021";
        ram_buffer(42363) := X"00602821";
        ram_buffer(42364) := X"00402021";
        ram_buffer(42365) := X"0C03167F";
        ram_buffer(42366) := X"00000000";
        ram_buffer(42367) := X"14400089";
        ram_buffer(42368) := X"00000000";
        ram_buffer(42369) := X"3C02100D";
        ram_buffer(42370) := X"2442A760";
        ram_buffer(42371) := X"AE020000";
        ram_buffer(42372) := X"24020001";
        ram_buffer(42373) := X"AE020004";
        ram_buffer(42374) := X"8FC200C0";
        ram_buffer(42375) := X"00000000";
        ram_buffer(42376) := X"24420001";
        ram_buffer(42377) := X"AFC200C0";
        ram_buffer(42378) := X"26100008";
        ram_buffer(42379) := X"8FC200BC";
        ram_buffer(42380) := X"00000000";
        ram_buffer(42381) := X"24420001";
        ram_buffer(42382) := X"AFC200BC";
        ram_buffer(42383) := X"8FC200BC";
        ram_buffer(42384) := X"00000000";
        ram_buffer(42385) := X"28420008";
        ram_buffer(42386) := X"1440000A";
        ram_buffer(42387) := X"00000000";
        ram_buffer(42388) := X"27C200B8";
        ram_buffer(42389) := X"00403021";
        ram_buffer(42390) := X"8FC501EC";
        ram_buffer(42391) := X"8FC401E8";
        ram_buffer(42392) := X"0C02EAF5";
        ram_buffer(42393) := X"00000000";
        ram_buffer(42394) := X"144004BC";
        ram_buffer(42395) := X"00000000";
        ram_buffer(42396) := X"27D000C4";
        ram_buffer(42397) := X"8FC300A8";
        ram_buffer(42398) := X"8FC200B4";
        ram_buffer(42399) := X"00000000";
        ram_buffer(42400) := X"0062102A";
        ram_buffer(42401) := X"14400004";
        ram_buffer(42402) := X"00000000";
        ram_buffer(42403) := X"32420001";
        ram_buffer(42404) := X"10400415";
        ram_buffer(42405) := X"00000000";
        ram_buffer(42406) := X"8FC20084";
        ram_buffer(42407) := X"00000000";
        ram_buffer(42408) := X"AE020000";
        ram_buffer(42409) := X"8FC20088";
        ram_buffer(42410) := X"00000000";
        ram_buffer(42411) := X"AE020004";
        ram_buffer(42412) := X"8FC300C0";
        ram_buffer(42413) := X"8FC20088";
        ram_buffer(42414) := X"00000000";
        ram_buffer(42415) := X"00621021";
        ram_buffer(42416) := X"AFC200C0";
        ram_buffer(42417) := X"26100008";
        ram_buffer(42418) := X"8FC200BC";
        ram_buffer(42419) := X"00000000";
        ram_buffer(42420) := X"24420001";
        ram_buffer(42421) := X"AFC200BC";
        ram_buffer(42422) := X"8FC200BC";
        ram_buffer(42423) := X"00000000";
        ram_buffer(42424) := X"28420008";
        ram_buffer(42425) := X"1440000A";
        ram_buffer(42426) := X"00000000";
        ram_buffer(42427) := X"27C200B8";
        ram_buffer(42428) := X"00403021";
        ram_buffer(42429) := X"8FC501EC";
        ram_buffer(42430) := X"8FC401E8";
        ram_buffer(42431) := X"0C02EAF5";
        ram_buffer(42432) := X"00000000";
        ram_buffer(42433) := X"14400498";
        ram_buffer(42434) := X"00000000";
        ram_buffer(42435) := X"27D000C4";
        ram_buffer(42436) := X"8FC200B4";
        ram_buffer(42437) := X"00000000";
        ram_buffer(42438) := X"2451FFFF";
        ram_buffer(42439) := X"1A2003F2";
        ram_buffer(42440) := X"00000000";
        ram_buffer(42441) := X"1000001E";
        ram_buffer(42442) := X"00000000";
        ram_buffer(42443) := X"3C02100D";
        ram_buffer(42444) := X"2442A8E0";
        ram_buffer(42445) := X"AE020000";
        ram_buffer(42446) := X"24020010";
        ram_buffer(42447) := X"AE020004";
        ram_buffer(42448) := X"8FC200C0";
        ram_buffer(42449) := X"00000000";
        ram_buffer(42450) := X"24420010";
        ram_buffer(42451) := X"AFC200C0";
        ram_buffer(42452) := X"26100008";
        ram_buffer(42453) := X"8FC200BC";
        ram_buffer(42454) := X"00000000";
        ram_buffer(42455) := X"24420001";
        ram_buffer(42456) := X"AFC200BC";
        ram_buffer(42457) := X"8FC200BC";
        ram_buffer(42458) := X"00000000";
        ram_buffer(42459) := X"28420008";
        ram_buffer(42460) := X"1440000A";
        ram_buffer(42461) := X"00000000";
        ram_buffer(42462) := X"27C200B8";
        ram_buffer(42463) := X"00403021";
        ram_buffer(42464) := X"8FC501EC";
        ram_buffer(42465) := X"8FC401E8";
        ram_buffer(42466) := X"0C02EAF5";
        ram_buffer(42467) := X"00000000";
        ram_buffer(42468) := X"14400478";
        ram_buffer(42469) := X"00000000";
        ram_buffer(42470) := X"27D000C4";
        ram_buffer(42471) := X"2631FFF0";
        ram_buffer(42472) := X"2A220011";
        ram_buffer(42473) := X"1040FFE1";
        ram_buffer(42474) := X"00000000";
        ram_buffer(42475) := X"3C02100D";
        ram_buffer(42476) := X"2442A8E0";
        ram_buffer(42477) := X"AE020000";
        ram_buffer(42478) := X"02201021";
        ram_buffer(42479) := X"AE020004";
        ram_buffer(42480) := X"8FC300C0";
        ram_buffer(42481) := X"02201021";
        ram_buffer(42482) := X"00621021";
        ram_buffer(42483) := X"AFC200C0";
        ram_buffer(42484) := X"26100008";
        ram_buffer(42485) := X"8FC200BC";
        ram_buffer(42486) := X"00000000";
        ram_buffer(42487) := X"24420001";
        ram_buffer(42488) := X"AFC200BC";
        ram_buffer(42489) := X"8FC200BC";
        ram_buffer(42490) := X"00000000";
        ram_buffer(42491) := X"28420008";
        ram_buffer(42492) := X"144003BD";
        ram_buffer(42493) := X"00000000";
        ram_buffer(42494) := X"27C200B8";
        ram_buffer(42495) := X"00403021";
        ram_buffer(42496) := X"8FC501EC";
        ram_buffer(42497) := X"8FC401E8";
        ram_buffer(42498) := X"0C02EAF5";
        ram_buffer(42499) := X"00000000";
        ram_buffer(42500) := X"1440045B";
        ram_buffer(42501) := X"00000000";
        ram_buffer(42502) := X"27D000C4";
        ram_buffer(42503) := X"100003B2";
        ram_buffer(42504) := X"00000000";
        ram_buffer(42505) := X"8FC200A8";
        ram_buffer(42506) := X"00000000";
        ram_buffer(42507) := X"1C4000A7";
        ram_buffer(42508) := X"00000000";
        ram_buffer(42509) := X"3C02100D";
        ram_buffer(42510) := X"2442A760";
        ram_buffer(42511) := X"AE020000";
        ram_buffer(42512) := X"24020001";
        ram_buffer(42513) := X"AE020004";
        ram_buffer(42514) := X"8FC200C0";
        ram_buffer(42515) := X"00000000";
        ram_buffer(42516) := X"24420001";
        ram_buffer(42517) := X"AFC200C0";
        ram_buffer(42518) := X"26100008";
        ram_buffer(42519) := X"8FC200BC";
        ram_buffer(42520) := X"00000000";
        ram_buffer(42521) := X"24420001";
        ram_buffer(42522) := X"AFC200BC";
        ram_buffer(42523) := X"8FC200BC";
        ram_buffer(42524) := X"00000000";
        ram_buffer(42525) := X"28420008";
        ram_buffer(42526) := X"1440000A";
        ram_buffer(42527) := X"00000000";
        ram_buffer(42528) := X"27C200B8";
        ram_buffer(42529) := X"00403021";
        ram_buffer(42530) := X"8FC501EC";
        ram_buffer(42531) := X"8FC401E8";
        ram_buffer(42532) := X"0C02EAF5";
        ram_buffer(42533) := X"00000000";
        ram_buffer(42534) := X"1440043C";
        ram_buffer(42535) := X"00000000";
        ram_buffer(42536) := X"27D000C4";
        ram_buffer(42537) := X"8FC200A8";
        ram_buffer(42538) := X"00000000";
        ram_buffer(42539) := X"14400008";
        ram_buffer(42540) := X"00000000";
        ram_buffer(42541) := X"8FC200B4";
        ram_buffer(42542) := X"00000000";
        ram_buffer(42543) := X"14400004";
        ram_buffer(42544) := X"00000000";
        ram_buffer(42545) := X"32420001";
        ram_buffer(42546) := X"10400387";
        ram_buffer(42547) := X"00000000";
        ram_buffer(42548) := X"8FC20084";
        ram_buffer(42549) := X"00000000";
        ram_buffer(42550) := X"AE020000";
        ram_buffer(42551) := X"8FC20088";
        ram_buffer(42552) := X"00000000";
        ram_buffer(42553) := X"AE020004";
        ram_buffer(42554) := X"8FC300C0";
        ram_buffer(42555) := X"8FC20088";
        ram_buffer(42556) := X"00000000";
        ram_buffer(42557) := X"00621021";
        ram_buffer(42558) := X"AFC200C0";
        ram_buffer(42559) := X"26100008";
        ram_buffer(42560) := X"8FC200BC";
        ram_buffer(42561) := X"00000000";
        ram_buffer(42562) := X"24420001";
        ram_buffer(42563) := X"AFC200BC";
        ram_buffer(42564) := X"8FC200BC";
        ram_buffer(42565) := X"00000000";
        ram_buffer(42566) := X"28420008";
        ram_buffer(42567) := X"1440000A";
        ram_buffer(42568) := X"00000000";
        ram_buffer(42569) := X"27C200B8";
        ram_buffer(42570) := X"00403021";
        ram_buffer(42571) := X"8FC501EC";
        ram_buffer(42572) := X"8FC401E8";
        ram_buffer(42573) := X"0C02EAF5";
        ram_buffer(42574) := X"00000000";
        ram_buffer(42575) := X"14400416";
        ram_buffer(42576) := X"00000000";
        ram_buffer(42577) := X"27D000C4";
        ram_buffer(42578) := X"8FC200A8";
        ram_buffer(42579) := X"00000000";
        ram_buffer(42580) := X"00028823";
        ram_buffer(42581) := X"1A20003F";
        ram_buffer(42582) := X"00000000";
        ram_buffer(42583) := X"1000001E";
        ram_buffer(42584) := X"00000000";
        ram_buffer(42585) := X"3C02100D";
        ram_buffer(42586) := X"2442A8E0";
        ram_buffer(42587) := X"AE020000";
        ram_buffer(42588) := X"24020010";
        ram_buffer(42589) := X"AE020004";
        ram_buffer(42590) := X"8FC200C0";
        ram_buffer(42591) := X"00000000";
        ram_buffer(42592) := X"24420010";
        ram_buffer(42593) := X"AFC200C0";
        ram_buffer(42594) := X"26100008";
        ram_buffer(42595) := X"8FC200BC";
        ram_buffer(42596) := X"00000000";
        ram_buffer(42597) := X"24420001";
        ram_buffer(42598) := X"AFC200BC";
        ram_buffer(42599) := X"8FC200BC";
        ram_buffer(42600) := X"00000000";
        ram_buffer(42601) := X"28420008";
        ram_buffer(42602) := X"1440000A";
        ram_buffer(42603) := X"00000000";
        ram_buffer(42604) := X"27C200B8";
        ram_buffer(42605) := X"00403021";
        ram_buffer(42606) := X"8FC501EC";
        ram_buffer(42607) := X"8FC401E8";
        ram_buffer(42608) := X"0C02EAF5";
        ram_buffer(42609) := X"00000000";
        ram_buffer(42610) := X"144003F6";
        ram_buffer(42611) := X"00000000";
        ram_buffer(42612) := X"27D000C4";
        ram_buffer(42613) := X"2631FFF0";
        ram_buffer(42614) := X"2A220011";
        ram_buffer(42615) := X"1040FFE1";
        ram_buffer(42616) := X"00000000";
        ram_buffer(42617) := X"3C02100D";
        ram_buffer(42618) := X"2442A8E0";
        ram_buffer(42619) := X"AE020000";
        ram_buffer(42620) := X"02201021";
        ram_buffer(42621) := X"AE020004";
        ram_buffer(42622) := X"8FC300C0";
        ram_buffer(42623) := X"02201021";
        ram_buffer(42624) := X"00621021";
        ram_buffer(42625) := X"AFC200C0";
        ram_buffer(42626) := X"26100008";
        ram_buffer(42627) := X"8FC200BC";
        ram_buffer(42628) := X"00000000";
        ram_buffer(42629) := X"24420001";
        ram_buffer(42630) := X"AFC200BC";
        ram_buffer(42631) := X"8FC200BC";
        ram_buffer(42632) := X"00000000";
        ram_buffer(42633) := X"28420008";
        ram_buffer(42634) := X"1440000A";
        ram_buffer(42635) := X"00000000";
        ram_buffer(42636) := X"27C200B8";
        ram_buffer(42637) := X"00403021";
        ram_buffer(42638) := X"8FC501EC";
        ram_buffer(42639) := X"8FC401E8";
        ram_buffer(42640) := X"0C02EAF5";
        ram_buffer(42641) := X"00000000";
        ram_buffer(42642) := X"144003D9";
        ram_buffer(42643) := X"00000000";
        ram_buffer(42644) := X"27D000C4";
        ram_buffer(42645) := X"AE130000";
        ram_buffer(42646) := X"8FC200B4";
        ram_buffer(42647) := X"00000000";
        ram_buffer(42648) := X"AE020004";
        ram_buffer(42649) := X"8FC300C0";
        ram_buffer(42650) := X"8FC200B4";
        ram_buffer(42651) := X"00000000";
        ram_buffer(42652) := X"00621021";
        ram_buffer(42653) := X"AFC200C0";
        ram_buffer(42654) := X"26100008";
        ram_buffer(42655) := X"8FC200BC";
        ram_buffer(42656) := X"00000000";
        ram_buffer(42657) := X"24420001";
        ram_buffer(42658) := X"AFC200BC";
        ram_buffer(42659) := X"8FC200BC";
        ram_buffer(42660) := X"00000000";
        ram_buffer(42661) := X"28420008";
        ram_buffer(42662) := X"14400313";
        ram_buffer(42663) := X"00000000";
        ram_buffer(42664) := X"27C200B8";
        ram_buffer(42665) := X"00403021";
        ram_buffer(42666) := X"8FC501EC";
        ram_buffer(42667) := X"8FC401E8";
        ram_buffer(42668) := X"0C02EAF5";
        ram_buffer(42669) := X"00000000";
        ram_buffer(42670) := X"144003C0";
        ram_buffer(42671) := X"00000000";
        ram_buffer(42672) := X"27D000C4";
        ram_buffer(42673) := X"10000308";
        ram_buffer(42674) := X"00000000";
        ram_buffer(42675) := X"AFD30098";
        ram_buffer(42676) := X"8FC200B4";
        ram_buffer(42677) := X"00000000";
        ram_buffer(42678) := X"00401821";
        ram_buffer(42679) := X"8FC20098";
        ram_buffer(42680) := X"00000000";
        ram_buffer(42681) := X"00431021";
        ram_buffer(42682) := X"00401821";
        ram_buffer(42683) := X"02601021";
        ram_buffer(42684) := X"00621023";
        ram_buffer(42685) := X"AFC20078";
        ram_buffer(42686) := X"8FC30078";
        ram_buffer(42687) := X"8FC2004C";
        ram_buffer(42688) := X"00000000";
        ram_buffer(42689) := X"0043102A";
        ram_buffer(42690) := X"10400004";
        ram_buffer(42691) := X"00000000";
        ram_buffer(42692) := X"8FC2004C";
        ram_buffer(42693) := X"00000000";
        ram_buffer(42694) := X"AFC20078";
        ram_buffer(42695) := X"8FC20078";
        ram_buffer(42696) := X"00000000";
        ram_buffer(42697) := X"1840001D";
        ram_buffer(42698) := X"00000000";
        ram_buffer(42699) := X"AE130000";
        ram_buffer(42700) := X"8FC20078";
        ram_buffer(42701) := X"00000000";
        ram_buffer(42702) := X"AE020004";
        ram_buffer(42703) := X"8FC300C0";
        ram_buffer(42704) := X"8FC20078";
        ram_buffer(42705) := X"00000000";
        ram_buffer(42706) := X"00621021";
        ram_buffer(42707) := X"AFC200C0";
        ram_buffer(42708) := X"26100008";
        ram_buffer(42709) := X"8FC200BC";
        ram_buffer(42710) := X"00000000";
        ram_buffer(42711) := X"24420001";
        ram_buffer(42712) := X"AFC200BC";
        ram_buffer(42713) := X"8FC200BC";
        ram_buffer(42714) := X"00000000";
        ram_buffer(42715) := X"28420008";
        ram_buffer(42716) := X"1440000A";
        ram_buffer(42717) := X"00000000";
        ram_buffer(42718) := X"27C200B8";
        ram_buffer(42719) := X"00403021";
        ram_buffer(42720) := X"8FC501EC";
        ram_buffer(42721) := X"8FC401E8";
        ram_buffer(42722) := X"0C02EAF5";
        ram_buffer(42723) := X"00000000";
        ram_buffer(42724) := X"1440038D";
        ram_buffer(42725) := X"00000000";
        ram_buffer(42726) := X"27D000C4";
        ram_buffer(42727) := X"8FC30078";
        ram_buffer(42728) := X"00000000";
        ram_buffer(42729) := X"04610002";
        ram_buffer(42730) := X"00000000";
        ram_buffer(42731) := X"00001821";
        ram_buffer(42732) := X"8FC2004C";
        ram_buffer(42733) := X"00000000";
        ram_buffer(42734) := X"00431023";
        ram_buffer(42735) := X"AFC20078";
        ram_buffer(42736) := X"8FC20078";
        ram_buffer(42737) := X"00000000";
        ram_buffer(42738) := X"18400046";
        ram_buffer(42739) := X"00000000";
        ram_buffer(42740) := X"10000021";
        ram_buffer(42741) := X"00000000";
        ram_buffer(42742) := X"3C02100D";
        ram_buffer(42743) := X"2442A8E0";
        ram_buffer(42744) := X"AE020000";
        ram_buffer(42745) := X"24020010";
        ram_buffer(42746) := X"AE020004";
        ram_buffer(42747) := X"8FC200C0";
        ram_buffer(42748) := X"00000000";
        ram_buffer(42749) := X"24420010";
        ram_buffer(42750) := X"AFC200C0";
        ram_buffer(42751) := X"26100008";
        ram_buffer(42752) := X"8FC200BC";
        ram_buffer(42753) := X"00000000";
        ram_buffer(42754) := X"24420001";
        ram_buffer(42755) := X"AFC200BC";
        ram_buffer(42756) := X"8FC200BC";
        ram_buffer(42757) := X"00000000";
        ram_buffer(42758) := X"28420008";
        ram_buffer(42759) := X"1440000A";
        ram_buffer(42760) := X"00000000";
        ram_buffer(42761) := X"27C200B8";
        ram_buffer(42762) := X"00403021";
        ram_buffer(42763) := X"8FC501EC";
        ram_buffer(42764) := X"8FC401E8";
        ram_buffer(42765) := X"0C02EAF5";
        ram_buffer(42766) := X"00000000";
        ram_buffer(42767) := X"14400365";
        ram_buffer(42768) := X"00000000";
        ram_buffer(42769) := X"27D000C4";
        ram_buffer(42770) := X"8FC20078";
        ram_buffer(42771) := X"00000000";
        ram_buffer(42772) := X"2442FFF0";
        ram_buffer(42773) := X"AFC20078";
        ram_buffer(42774) := X"8FC20078";
        ram_buffer(42775) := X"00000000";
        ram_buffer(42776) := X"28420011";
        ram_buffer(42777) := X"1040FFDC";
        ram_buffer(42778) := X"00000000";
        ram_buffer(42779) := X"3C02100D";
        ram_buffer(42780) := X"2442A8E0";
        ram_buffer(42781) := X"AE020000";
        ram_buffer(42782) := X"8FC20078";
        ram_buffer(42783) := X"00000000";
        ram_buffer(42784) := X"AE020004";
        ram_buffer(42785) := X"8FC300C0";
        ram_buffer(42786) := X"8FC20078";
        ram_buffer(42787) := X"00000000";
        ram_buffer(42788) := X"00621021";
        ram_buffer(42789) := X"AFC200C0";
        ram_buffer(42790) := X"26100008";
        ram_buffer(42791) := X"8FC200BC";
        ram_buffer(42792) := X"00000000";
        ram_buffer(42793) := X"24420001";
        ram_buffer(42794) := X"AFC200BC";
        ram_buffer(42795) := X"8FC200BC";
        ram_buffer(42796) := X"00000000";
        ram_buffer(42797) := X"28420008";
        ram_buffer(42798) := X"1440000A";
        ram_buffer(42799) := X"00000000";
        ram_buffer(42800) := X"27C200B8";
        ram_buffer(42801) := X"00403021";
        ram_buffer(42802) := X"8FC501EC";
        ram_buffer(42803) := X"8FC401E8";
        ram_buffer(42804) := X"0C02EAF5";
        ram_buffer(42805) := X"00000000";
        ram_buffer(42806) := X"14400341";
        ram_buffer(42807) := X"00000000";
        ram_buffer(42808) := X"27D000C4";
        ram_buffer(42809) := X"8FC2004C";
        ram_buffer(42810) := X"00000000";
        ram_buffer(42811) := X"02629821";
        ram_buffer(42812) := X"32420400";
        ram_buffer(42813) := X"104000DD";
        ram_buffer(42814) := X"00000000";
        ram_buffer(42815) := X"100000C4";
        ram_buffer(42816) := X"00000000";
        ram_buffer(42817) := X"8FC20054";
        ram_buffer(42818) := X"00000000";
        ram_buffer(42819) := X"18400007";
        ram_buffer(42820) := X"00000000";
        ram_buffer(42821) := X"8FC20054";
        ram_buffer(42822) := X"00000000";
        ram_buffer(42823) := X"2442FFFF";
        ram_buffer(42824) := X"AFC20054";
        ram_buffer(42825) := X"10000009";
        ram_buffer(42826) := X"00000000";
        ram_buffer(42827) := X"8FC20044";
        ram_buffer(42828) := X"00000000";
        ram_buffer(42829) := X"2442FFFF";
        ram_buffer(42830) := X"AFC20044";
        ram_buffer(42831) := X"8FC20050";
        ram_buffer(42832) := X"00000000";
        ram_buffer(42833) := X"2442FFFF";
        ram_buffer(42834) := X"AFC20050";
        ram_buffer(42835) := X"8FC2003C";
        ram_buffer(42836) := X"00000000";
        ram_buffer(42837) := X"AE020000";
        ram_buffer(42838) := X"8FC20040";
        ram_buffer(42839) := X"00000000";
        ram_buffer(42840) := X"AE020004";
        ram_buffer(42841) := X"8FC300C0";
        ram_buffer(42842) := X"8FC20040";
        ram_buffer(42843) := X"00000000";
        ram_buffer(42844) := X"00621021";
        ram_buffer(42845) := X"AFC200C0";
        ram_buffer(42846) := X"26100008";
        ram_buffer(42847) := X"8FC200BC";
        ram_buffer(42848) := X"00000000";
        ram_buffer(42849) := X"24420001";
        ram_buffer(42850) := X"AFC200BC";
        ram_buffer(42851) := X"8FC200BC";
        ram_buffer(42852) := X"00000000";
        ram_buffer(42853) := X"28420008";
        ram_buffer(42854) := X"1440000A";
        ram_buffer(42855) := X"00000000";
        ram_buffer(42856) := X"27C200B8";
        ram_buffer(42857) := X"00403021";
        ram_buffer(42858) := X"8FC501EC";
        ram_buffer(42859) := X"8FC401E8";
        ram_buffer(42860) := X"0C02EAF5";
        ram_buffer(42861) := X"00000000";
        ram_buffer(42862) := X"1440030C";
        ram_buffer(42863) := X"00000000";
        ram_buffer(42864) := X"27D000C4";
        ram_buffer(42865) := X"8FC200B4";
        ram_buffer(42866) := X"00000000";
        ram_buffer(42867) := X"00401821";
        ram_buffer(42868) := X"8FC20098";
        ram_buffer(42869) := X"00000000";
        ram_buffer(42870) := X"00431021";
        ram_buffer(42871) := X"00401821";
        ram_buffer(42872) := X"02601021";
        ram_buffer(42873) := X"00621023";
        ram_buffer(42874) := X"AFC2007C";
        ram_buffer(42875) := X"8FC20044";
        ram_buffer(42876) := X"00000000";
        ram_buffer(42877) := X"80420000";
        ram_buffer(42878) := X"00000000";
        ram_buffer(42879) := X"00401821";
        ram_buffer(42880) := X"8FC2007C";
        ram_buffer(42881) := X"00000000";
        ram_buffer(42882) := X"0062102A";
        ram_buffer(42883) := X"10400006";
        ram_buffer(42884) := X"00000000";
        ram_buffer(42885) := X"8FC20044";
        ram_buffer(42886) := X"00000000";
        ram_buffer(42887) := X"80420000";
        ram_buffer(42888) := X"00000000";
        ram_buffer(42889) := X"AFC2007C";
        ram_buffer(42890) := X"8FC2007C";
        ram_buffer(42891) := X"00000000";
        ram_buffer(42892) := X"1840001D";
        ram_buffer(42893) := X"00000000";
        ram_buffer(42894) := X"AE130000";
        ram_buffer(42895) := X"8FC2007C";
        ram_buffer(42896) := X"00000000";
        ram_buffer(42897) := X"AE020004";
        ram_buffer(42898) := X"8FC300C0";
        ram_buffer(42899) := X"8FC2007C";
        ram_buffer(42900) := X"00000000";
        ram_buffer(42901) := X"00621021";
        ram_buffer(42902) := X"AFC200C0";
        ram_buffer(42903) := X"26100008";
        ram_buffer(42904) := X"8FC200BC";
        ram_buffer(42905) := X"00000000";
        ram_buffer(42906) := X"24420001";
        ram_buffer(42907) := X"AFC200BC";
        ram_buffer(42908) := X"8FC200BC";
        ram_buffer(42909) := X"00000000";
        ram_buffer(42910) := X"28420008";
        ram_buffer(42911) := X"1440000A";
        ram_buffer(42912) := X"00000000";
        ram_buffer(42913) := X"27C200B8";
        ram_buffer(42914) := X"00403021";
        ram_buffer(42915) := X"8FC501EC";
        ram_buffer(42916) := X"8FC401E8";
        ram_buffer(42917) := X"0C02EAF5";
        ram_buffer(42918) := X"00000000";
        ram_buffer(42919) := X"144002D6";
        ram_buffer(42920) := X"00000000";
        ram_buffer(42921) := X"27D000C4";
        ram_buffer(42922) := X"8FC20044";
        ram_buffer(42923) := X"00000000";
        ram_buffer(42924) := X"80420000";
        ram_buffer(42925) := X"00000000";
        ram_buffer(42926) := X"00401821";
        ram_buffer(42927) := X"8FC2007C";
        ram_buffer(42928) := X"00000000";
        ram_buffer(42929) := X"04410002";
        ram_buffer(42930) := X"00000000";
        ram_buffer(42931) := X"00001021";
        ram_buffer(42932) := X"00621023";
        ram_buffer(42933) := X"AFC2007C";
        ram_buffer(42934) := X"8FC2007C";
        ram_buffer(42935) := X"00000000";
        ram_buffer(42936) := X"18400046";
        ram_buffer(42937) := X"00000000";
        ram_buffer(42938) := X"10000021";
        ram_buffer(42939) := X"00000000";
        ram_buffer(42940) := X"3C02100D";
        ram_buffer(42941) := X"2442A8E0";
        ram_buffer(42942) := X"AE020000";
        ram_buffer(42943) := X"24020010";
        ram_buffer(42944) := X"AE020004";
        ram_buffer(42945) := X"8FC200C0";
        ram_buffer(42946) := X"00000000";
        ram_buffer(42947) := X"24420010";
        ram_buffer(42948) := X"AFC200C0";
        ram_buffer(42949) := X"26100008";
        ram_buffer(42950) := X"8FC200BC";
        ram_buffer(42951) := X"00000000";
        ram_buffer(42952) := X"24420001";
        ram_buffer(42953) := X"AFC200BC";
        ram_buffer(42954) := X"8FC200BC";
        ram_buffer(42955) := X"00000000";
        ram_buffer(42956) := X"28420008";
        ram_buffer(42957) := X"1440000A";
        ram_buffer(42958) := X"00000000";
        ram_buffer(42959) := X"27C200B8";
        ram_buffer(42960) := X"00403021";
        ram_buffer(42961) := X"8FC501EC";
        ram_buffer(42962) := X"8FC401E8";
        ram_buffer(42963) := X"0C02EAF5";
        ram_buffer(42964) := X"00000000";
        ram_buffer(42965) := X"144002AB";
        ram_buffer(42966) := X"00000000";
        ram_buffer(42967) := X"27D000C4";
        ram_buffer(42968) := X"8FC2007C";
        ram_buffer(42969) := X"00000000";
        ram_buffer(42970) := X"2442FFF0";
        ram_buffer(42971) := X"AFC2007C";
        ram_buffer(42972) := X"8FC2007C";
        ram_buffer(42973) := X"00000000";
        ram_buffer(42974) := X"28420011";
        ram_buffer(42975) := X"1040FFDC";
        ram_buffer(42976) := X"00000000";
        ram_buffer(42977) := X"3C02100D";
        ram_buffer(42978) := X"2442A8E0";
        ram_buffer(42979) := X"AE020000";
        ram_buffer(42980) := X"8FC2007C";
        ram_buffer(42981) := X"00000000";
        ram_buffer(42982) := X"AE020004";
        ram_buffer(42983) := X"8FC300C0";
        ram_buffer(42984) := X"8FC2007C";
        ram_buffer(42985) := X"00000000";
        ram_buffer(42986) := X"00621021";
        ram_buffer(42987) := X"AFC200C0";
        ram_buffer(42988) := X"26100008";
        ram_buffer(42989) := X"8FC200BC";
        ram_buffer(42990) := X"00000000";
        ram_buffer(42991) := X"24420001";
        ram_buffer(42992) := X"AFC200BC";
        ram_buffer(42993) := X"8FC200BC";
        ram_buffer(42994) := X"00000000";
        ram_buffer(42995) := X"28420008";
        ram_buffer(42996) := X"1440000A";
        ram_buffer(42997) := X"00000000";
        ram_buffer(42998) := X"27C200B8";
        ram_buffer(42999) := X"00403021";
        ram_buffer(43000) := X"8FC501EC";
        ram_buffer(43001) := X"8FC401E8";
        ram_buffer(43002) := X"0C02EAF5";
        ram_buffer(43003) := X"00000000";
        ram_buffer(43004) := X"14400287";
        ram_buffer(43005) := X"00000000";
        ram_buffer(43006) := X"27D000C4";
        ram_buffer(43007) := X"8FC20044";
        ram_buffer(43008) := X"00000000";
        ram_buffer(43009) := X"80420000";
        ram_buffer(43010) := X"00000000";
        ram_buffer(43011) := X"02629821";
        ram_buffer(43012) := X"8FC20050";
        ram_buffer(43013) := X"00000000";
        ram_buffer(43014) := X"1C40FF3A";
        ram_buffer(43015) := X"00000000";
        ram_buffer(43016) := X"8FC20054";
        ram_buffer(43017) := X"00000000";
        ram_buffer(43018) := X"1C40FF36";
        ram_buffer(43019) := X"00000000";
        ram_buffer(43020) := X"8FC200B4";
        ram_buffer(43021) := X"00000000";
        ram_buffer(43022) := X"00401821";
        ram_buffer(43023) := X"8FC20098";
        ram_buffer(43024) := X"00000000";
        ram_buffer(43025) := X"00431021";
        ram_buffer(43026) := X"0053102B";
        ram_buffer(43027) := X"10400007";
        ram_buffer(43028) := X"00000000";
        ram_buffer(43029) := X"8FC200B4";
        ram_buffer(43030) := X"00000000";
        ram_buffer(43031) := X"00401821";
        ram_buffer(43032) := X"8FC20098";
        ram_buffer(43033) := X"00000000";
        ram_buffer(43034) := X"00439821";
        ram_buffer(43035) := X"8FC300A8";
        ram_buffer(43036) := X"8FC200B4";
        ram_buffer(43037) := X"00000000";
        ram_buffer(43038) := X"0062102A";
        ram_buffer(43039) := X"14400004";
        ram_buffer(43040) := X"00000000";
        ram_buffer(43041) := X"32420001";
        ram_buffer(43042) := X"1040001F";
        ram_buffer(43043) := X"00000000";
        ram_buffer(43044) := X"8FC20084";
        ram_buffer(43045) := X"00000000";
        ram_buffer(43046) := X"AE020000";
        ram_buffer(43047) := X"8FC20088";
        ram_buffer(43048) := X"00000000";
        ram_buffer(43049) := X"AE020004";
        ram_buffer(43050) := X"8FC300C0";
        ram_buffer(43051) := X"8FC20088";
        ram_buffer(43052) := X"00000000";
        ram_buffer(43053) := X"00621021";
        ram_buffer(43054) := X"AFC200C0";
        ram_buffer(43055) := X"26100008";
        ram_buffer(43056) := X"8FC200BC";
        ram_buffer(43057) := X"00000000";
        ram_buffer(43058) := X"24420001";
        ram_buffer(43059) := X"AFC200BC";
        ram_buffer(43060) := X"8FC200BC";
        ram_buffer(43061) := X"00000000";
        ram_buffer(43062) := X"28420008";
        ram_buffer(43063) := X"1440000A";
        ram_buffer(43064) := X"00000000";
        ram_buffer(43065) := X"27C200B8";
        ram_buffer(43066) := X"00403021";
        ram_buffer(43067) := X"8FC501EC";
        ram_buffer(43068) := X"8FC401E8";
        ram_buffer(43069) := X"0C02EAF5";
        ram_buffer(43070) := X"00000000";
        ram_buffer(43071) := X"14400247";
        ram_buffer(43072) := X"00000000";
        ram_buffer(43073) := X"27D000C4";
        ram_buffer(43074) := X"8FC200B4";
        ram_buffer(43075) := X"00000000";
        ram_buffer(43076) := X"00401821";
        ram_buffer(43077) := X"8FC20098";
        ram_buffer(43078) := X"00000000";
        ram_buffer(43079) := X"00431021";
        ram_buffer(43080) := X"00401821";
        ram_buffer(43081) := X"02601021";
        ram_buffer(43082) := X"00621023";
        ram_buffer(43083) := X"AFC20080";
        ram_buffer(43084) := X"8FC300B4";
        ram_buffer(43085) := X"8FC200A8";
        ram_buffer(43086) := X"00000000";
        ram_buffer(43087) := X"00621823";
        ram_buffer(43088) := X"8FC20080";
        ram_buffer(43089) := X"00000000";
        ram_buffer(43090) := X"0062102A";
        ram_buffer(43091) := X"10400006";
        ram_buffer(43092) := X"00000000";
        ram_buffer(43093) := X"8FC300B4";
        ram_buffer(43094) := X"8FC200A8";
        ram_buffer(43095) := X"00000000";
        ram_buffer(43096) := X"00621023";
        ram_buffer(43097) := X"AFC20080";
        ram_buffer(43098) := X"8FC20080";
        ram_buffer(43099) := X"00000000";
        ram_buffer(43100) := X"1840001D";
        ram_buffer(43101) := X"00000000";
        ram_buffer(43102) := X"AE130000";
        ram_buffer(43103) := X"8FC20080";
        ram_buffer(43104) := X"00000000";
        ram_buffer(43105) := X"AE020004";
        ram_buffer(43106) := X"8FC300C0";
        ram_buffer(43107) := X"8FC20080";
        ram_buffer(43108) := X"00000000";
        ram_buffer(43109) := X"00621021";
        ram_buffer(43110) := X"AFC200C0";
        ram_buffer(43111) := X"26100008";
        ram_buffer(43112) := X"8FC200BC";
        ram_buffer(43113) := X"00000000";
        ram_buffer(43114) := X"24420001";
        ram_buffer(43115) := X"AFC200BC";
        ram_buffer(43116) := X"8FC200BC";
        ram_buffer(43117) := X"00000000";
        ram_buffer(43118) := X"28420008";
        ram_buffer(43119) := X"1440000A";
        ram_buffer(43120) := X"00000000";
        ram_buffer(43121) := X"27C200B8";
        ram_buffer(43122) := X"00403021";
        ram_buffer(43123) := X"8FC501EC";
        ram_buffer(43124) := X"8FC401E8";
        ram_buffer(43125) := X"0C02EAF5";
        ram_buffer(43126) := X"00000000";
        ram_buffer(43127) := X"14400212";
        ram_buffer(43128) := X"00000000";
        ram_buffer(43129) := X"27D000C4";
        ram_buffer(43130) := X"8FC300B4";
        ram_buffer(43131) := X"8FC200A8";
        ram_buffer(43132) := X"00000000";
        ram_buffer(43133) := X"00621823";
        ram_buffer(43134) := X"8FC20080";
        ram_buffer(43135) := X"00000000";
        ram_buffer(43136) := X"04410002";
        ram_buffer(43137) := X"00000000";
        ram_buffer(43138) := X"00001021";
        ram_buffer(43139) := X"00621023";
        ram_buffer(43140) := X"AFC20080";
        ram_buffer(43141) := X"8FC20080";
        ram_buffer(43142) := X"00000000";
        ram_buffer(43143) := X"18400132";
        ram_buffer(43144) := X"00000000";
        ram_buffer(43145) := X"10000021";
        ram_buffer(43146) := X"00000000";
        ram_buffer(43147) := X"3C02100D";
        ram_buffer(43148) := X"2442A8E0";
        ram_buffer(43149) := X"AE020000";
        ram_buffer(43150) := X"24020010";
        ram_buffer(43151) := X"AE020004";
        ram_buffer(43152) := X"8FC200C0";
        ram_buffer(43153) := X"00000000";
        ram_buffer(43154) := X"24420010";
        ram_buffer(43155) := X"AFC200C0";
        ram_buffer(43156) := X"26100008";
        ram_buffer(43157) := X"8FC200BC";
        ram_buffer(43158) := X"00000000";
        ram_buffer(43159) := X"24420001";
        ram_buffer(43160) := X"AFC200BC";
        ram_buffer(43161) := X"8FC200BC";
        ram_buffer(43162) := X"00000000";
        ram_buffer(43163) := X"28420008";
        ram_buffer(43164) := X"1440000A";
        ram_buffer(43165) := X"00000000";
        ram_buffer(43166) := X"27C200B8";
        ram_buffer(43167) := X"00403021";
        ram_buffer(43168) := X"8FC501EC";
        ram_buffer(43169) := X"8FC401E8";
        ram_buffer(43170) := X"0C02EAF5";
        ram_buffer(43171) := X"00000000";
        ram_buffer(43172) := X"144001E8";
        ram_buffer(43173) := X"00000000";
        ram_buffer(43174) := X"27D000C4";
        ram_buffer(43175) := X"8FC20080";
        ram_buffer(43176) := X"00000000";
        ram_buffer(43177) := X"2442FFF0";
        ram_buffer(43178) := X"AFC20080";
        ram_buffer(43179) := X"8FC20080";
        ram_buffer(43180) := X"00000000";
        ram_buffer(43181) := X"28420011";
        ram_buffer(43182) := X"1040FFDC";
        ram_buffer(43183) := X"00000000";
        ram_buffer(43184) := X"3C02100D";
        ram_buffer(43185) := X"2442A8E0";
        ram_buffer(43186) := X"AE020000";
        ram_buffer(43187) := X"8FC20080";
        ram_buffer(43188) := X"00000000";
        ram_buffer(43189) := X"AE020004";
        ram_buffer(43190) := X"8FC300C0";
        ram_buffer(43191) := X"8FC20080";
        ram_buffer(43192) := X"00000000";
        ram_buffer(43193) := X"00621021";
        ram_buffer(43194) := X"AFC200C0";
        ram_buffer(43195) := X"26100008";
        ram_buffer(43196) := X"8FC200BC";
        ram_buffer(43197) := X"00000000";
        ram_buffer(43198) := X"24420001";
        ram_buffer(43199) := X"AFC200BC";
        ram_buffer(43200) := X"8FC200BC";
        ram_buffer(43201) := X"00000000";
        ram_buffer(43202) := X"28420008";
        ram_buffer(43203) := X"144000F6";
        ram_buffer(43204) := X"00000000";
        ram_buffer(43205) := X"27C200B8";
        ram_buffer(43206) := X"00403021";
        ram_buffer(43207) := X"8FC501EC";
        ram_buffer(43208) := X"8FC401E8";
        ram_buffer(43209) := X"0C02EAF5";
        ram_buffer(43210) := X"00000000";
        ram_buffer(43211) := X"144001C4";
        ram_buffer(43212) := X"00000000";
        ram_buffer(43213) := X"27D000C4";
        ram_buffer(43214) := X"100000EB";
        ram_buffer(43215) := X"00000000";
        ram_buffer(43216) := X"8FC200B4";
        ram_buffer(43217) := X"00000000";
        ram_buffer(43218) := X"28420002";
        ram_buffer(43219) := X"10400004";
        ram_buffer(43220) := X"00000000";
        ram_buffer(43221) := X"32420001";
        ram_buffer(43222) := X"104000A9";
        ram_buffer(43223) := X"00000000";
        ram_buffer(43224) := X"AE130000";
        ram_buffer(43225) := X"24020001";
        ram_buffer(43226) := X"AE020004";
        ram_buffer(43227) := X"8FC200C0";
        ram_buffer(43228) := X"00000000";
        ram_buffer(43229) := X"24420001";
        ram_buffer(43230) := X"AFC200C0";
        ram_buffer(43231) := X"26100008";
        ram_buffer(43232) := X"8FC200BC";
        ram_buffer(43233) := X"00000000";
        ram_buffer(43234) := X"24420001";
        ram_buffer(43235) := X"AFC200BC";
        ram_buffer(43236) := X"8FC200BC";
        ram_buffer(43237) := X"00000000";
        ram_buffer(43238) := X"28420008";
        ram_buffer(43239) := X"1440000A";
        ram_buffer(43240) := X"00000000";
        ram_buffer(43241) := X"27C200B8";
        ram_buffer(43242) := X"00403021";
        ram_buffer(43243) := X"8FC501EC";
        ram_buffer(43244) := X"8FC401E8";
        ram_buffer(43245) := X"0C02EAF5";
        ram_buffer(43246) := X"00000000";
        ram_buffer(43247) := X"144001A3";
        ram_buffer(43248) := X"00000000";
        ram_buffer(43249) := X"27D000C4";
        ram_buffer(43250) := X"26730001";
        ram_buffer(43251) := X"8FC20084";
        ram_buffer(43252) := X"00000000";
        ram_buffer(43253) := X"AE020000";
        ram_buffer(43254) := X"8FC20088";
        ram_buffer(43255) := X"00000000";
        ram_buffer(43256) := X"AE020004";
        ram_buffer(43257) := X"8FC300C0";
        ram_buffer(43258) := X"8FC20088";
        ram_buffer(43259) := X"00000000";
        ram_buffer(43260) := X"00621021";
        ram_buffer(43261) := X"AFC200C0";
        ram_buffer(43262) := X"26100008";
        ram_buffer(43263) := X"8FC200BC";
        ram_buffer(43264) := X"00000000";
        ram_buffer(43265) := X"24420001";
        ram_buffer(43266) := X"AFC200BC";
        ram_buffer(43267) := X"8FC200BC";
        ram_buffer(43268) := X"00000000";
        ram_buffer(43269) := X"28420008";
        ram_buffer(43270) := X"1440000A";
        ram_buffer(43271) := X"00000000";
        ram_buffer(43272) := X"27C200B8";
        ram_buffer(43273) := X"00403021";
        ram_buffer(43274) := X"8FC501EC";
        ram_buffer(43275) := X"8FC401E8";
        ram_buffer(43276) := X"0C02EAF5";
        ram_buffer(43277) := X"00000000";
        ram_buffer(43278) := X"14400187";
        ram_buffer(43279) := X"00000000";
        ram_buffer(43280) := X"27D000C4";
        ram_buffer(43281) := X"8FC300A4";
        ram_buffer(43282) := X"8FC200A0";
        ram_buffer(43283) := X"00003821";
        ram_buffer(43284) := X"00003021";
        ram_buffer(43285) := X"00602821";
        ram_buffer(43286) := X"00402021";
        ram_buffer(43287) := X"0C03167F";
        ram_buffer(43288) := X"00000000";
        ram_buffer(43289) := X"10400021";
        ram_buffer(43290) := X"00000000";
        ram_buffer(43291) := X"AE130000";
        ram_buffer(43292) := X"8FC200B4";
        ram_buffer(43293) := X"00000000";
        ram_buffer(43294) := X"2442FFFF";
        ram_buffer(43295) := X"AE020004";
        ram_buffer(43296) := X"8FC300C0";
        ram_buffer(43297) := X"8FC200B4";
        ram_buffer(43298) := X"00000000";
        ram_buffer(43299) := X"00621021";
        ram_buffer(43300) := X"2442FFFF";
        ram_buffer(43301) := X"AFC200C0";
        ram_buffer(43302) := X"26100008";
        ram_buffer(43303) := X"8FC200BC";
        ram_buffer(43304) := X"00000000";
        ram_buffer(43305) := X"24420001";
        ram_buffer(43306) := X"AFC200BC";
        ram_buffer(43307) := X"8FC200BC";
        ram_buffer(43308) := X"00000000";
        ram_buffer(43309) := X"28420008";
        ram_buffer(43310) := X"1440006D";
        ram_buffer(43311) := X"00000000";
        ram_buffer(43312) := X"27C200B8";
        ram_buffer(43313) := X"00403021";
        ram_buffer(43314) := X"8FC501EC";
        ram_buffer(43315) := X"8FC401E8";
        ram_buffer(43316) := X"0C02EAF5";
        ram_buffer(43317) := X"00000000";
        ram_buffer(43318) := X"14400162";
        ram_buffer(43319) := X"00000000";
        ram_buffer(43320) := X"27D000C4";
        ram_buffer(43321) := X"10000062";
        ram_buffer(43322) := X"00000000";
        ram_buffer(43323) := X"8FC200B4";
        ram_buffer(43324) := X"00000000";
        ram_buffer(43325) := X"2451FFFF";
        ram_buffer(43326) := X"1A20005D";
        ram_buffer(43327) := X"00000000";
        ram_buffer(43328) := X"1000001E";
        ram_buffer(43329) := X"00000000";
        ram_buffer(43330) := X"3C02100D";
        ram_buffer(43331) := X"2442A8E0";
        ram_buffer(43332) := X"AE020000";
        ram_buffer(43333) := X"24020010";
        ram_buffer(43334) := X"AE020004";
        ram_buffer(43335) := X"8FC200C0";
        ram_buffer(43336) := X"00000000";
        ram_buffer(43337) := X"24420010";
        ram_buffer(43338) := X"AFC200C0";
        ram_buffer(43339) := X"26100008";
        ram_buffer(43340) := X"8FC200BC";
        ram_buffer(43341) := X"00000000";
        ram_buffer(43342) := X"24420001";
        ram_buffer(43343) := X"AFC200BC";
        ram_buffer(43344) := X"8FC200BC";
        ram_buffer(43345) := X"00000000";
        ram_buffer(43346) := X"28420008";
        ram_buffer(43347) := X"1440000A";
        ram_buffer(43348) := X"00000000";
        ram_buffer(43349) := X"27C200B8";
        ram_buffer(43350) := X"00403021";
        ram_buffer(43351) := X"8FC501EC";
        ram_buffer(43352) := X"8FC401E8";
        ram_buffer(43353) := X"0C02EAF5";
        ram_buffer(43354) := X"00000000";
        ram_buffer(43355) := X"14400140";
        ram_buffer(43356) := X"00000000";
        ram_buffer(43357) := X"27D000C4";
        ram_buffer(43358) := X"2631FFF0";
        ram_buffer(43359) := X"2A220011";
        ram_buffer(43360) := X"1040FFE1";
        ram_buffer(43361) := X"00000000";
        ram_buffer(43362) := X"3C02100D";
        ram_buffer(43363) := X"2442A8E0";
        ram_buffer(43364) := X"AE020000";
        ram_buffer(43365) := X"02201021";
        ram_buffer(43366) := X"AE020004";
        ram_buffer(43367) := X"8FC300C0";
        ram_buffer(43368) := X"02201021";
        ram_buffer(43369) := X"00621021";
        ram_buffer(43370) := X"AFC200C0";
        ram_buffer(43371) := X"26100008";
        ram_buffer(43372) := X"8FC200BC";
        ram_buffer(43373) := X"00000000";
        ram_buffer(43374) := X"24420001";
        ram_buffer(43375) := X"AFC200BC";
        ram_buffer(43376) := X"8FC200BC";
        ram_buffer(43377) := X"00000000";
        ram_buffer(43378) := X"28420008";
        ram_buffer(43379) := X"14400028";
        ram_buffer(43380) := X"00000000";
        ram_buffer(43381) := X"27C200B8";
        ram_buffer(43382) := X"00403021";
        ram_buffer(43383) := X"8FC501EC";
        ram_buffer(43384) := X"8FC401E8";
        ram_buffer(43385) := X"0C02EAF5";
        ram_buffer(43386) := X"00000000";
        ram_buffer(43387) := X"14400123";
        ram_buffer(43388) := X"00000000";
        ram_buffer(43389) := X"27D000C4";
        ram_buffer(43390) := X"1000001D";
        ram_buffer(43391) := X"00000000";
        ram_buffer(43392) := X"AE130000";
        ram_buffer(43393) := X"24020001";
        ram_buffer(43394) := X"AE020004";
        ram_buffer(43395) := X"8FC200C0";
        ram_buffer(43396) := X"00000000";
        ram_buffer(43397) := X"24420001";
        ram_buffer(43398) := X"AFC200C0";
        ram_buffer(43399) := X"26100008";
        ram_buffer(43400) := X"8FC200BC";
        ram_buffer(43401) := X"00000000";
        ram_buffer(43402) := X"24420001";
        ram_buffer(43403) := X"AFC200BC";
        ram_buffer(43404) := X"8FC200BC";
        ram_buffer(43405) := X"00000000";
        ram_buffer(43406) := X"28420008";
        ram_buffer(43407) := X"1440000D";
        ram_buffer(43408) := X"00000000";
        ram_buffer(43409) := X"27C200B8";
        ram_buffer(43410) := X"00403021";
        ram_buffer(43411) := X"8FC501EC";
        ram_buffer(43412) := X"8FC401E8";
        ram_buffer(43413) := X"0C02EAF5";
        ram_buffer(43414) := X"00000000";
        ram_buffer(43415) := X"1440010A";
        ram_buffer(43416) := X"00000000";
        ram_buffer(43417) := X"27D000C4";
        ram_buffer(43418) := X"10000002";
        ram_buffer(43419) := X"00000000";
        ram_buffer(43420) := X"00000000";
        ram_buffer(43421) := X"27C200AC";
        ram_buffer(43422) := X"AE020000";
        ram_buffer(43423) := X"8FC20048";
        ram_buffer(43424) := X"00000000";
        ram_buffer(43425) := X"AE020004";
        ram_buffer(43426) := X"8FC300C0";
        ram_buffer(43427) := X"8FC20048";
        ram_buffer(43428) := X"00000000";
        ram_buffer(43429) := X"00621021";
        ram_buffer(43430) := X"AFC200C0";
        ram_buffer(43431) := X"26100008";
        ram_buffer(43432) := X"8FC200BC";
        ram_buffer(43433) := X"00000000";
        ram_buffer(43434) := X"24420001";
        ram_buffer(43435) := X"AFC200BC";
        ram_buffer(43436) := X"8FC200BC";
        ram_buffer(43437) := X"00000000";
        ram_buffer(43438) := X"28420008";
        ram_buffer(43439) := X"1440000A";
        ram_buffer(43440) := X"00000000";
        ram_buffer(43441) := X"27C200B8";
        ram_buffer(43442) := X"00403021";
        ram_buffer(43443) := X"8FC501EC";
        ram_buffer(43444) := X"8FC401E8";
        ram_buffer(43445) := X"0C02EAF5";
        ram_buffer(43446) := X"00000000";
        ram_buffer(43447) := X"144000ED";
        ram_buffer(43448) := X"00000000";
        ram_buffer(43449) := X"27D000C4";
        ram_buffer(43450) := X"32420004";
        ram_buffer(43451) := X"10400045";
        ram_buffer(43452) := X"00000000";
        ram_buffer(43453) := X"8FC30034";
        ram_buffer(43454) := X"8FC20068";
        ram_buffer(43455) := X"00000000";
        ram_buffer(43456) := X"00628823";
        ram_buffer(43457) := X"1A20003F";
        ram_buffer(43458) := X"00000000";
        ram_buffer(43459) := X"1000001E";
        ram_buffer(43460) := X"00000000";
        ram_buffer(43461) := X"3C02100D";
        ram_buffer(43462) := X"2442A8D0";
        ram_buffer(43463) := X"AE020000";
        ram_buffer(43464) := X"24020010";
        ram_buffer(43465) := X"AE020004";
        ram_buffer(43466) := X"8FC200C0";
        ram_buffer(43467) := X"00000000";
        ram_buffer(43468) := X"24420010";
        ram_buffer(43469) := X"AFC200C0";
        ram_buffer(43470) := X"26100008";
        ram_buffer(43471) := X"8FC200BC";
        ram_buffer(43472) := X"00000000";
        ram_buffer(43473) := X"24420001";
        ram_buffer(43474) := X"AFC200BC";
        ram_buffer(43475) := X"8FC200BC";
        ram_buffer(43476) := X"00000000";
        ram_buffer(43477) := X"28420008";
        ram_buffer(43478) := X"1440000A";
        ram_buffer(43479) := X"00000000";
        ram_buffer(43480) := X"27C200B8";
        ram_buffer(43481) := X"00403021";
        ram_buffer(43482) := X"8FC501EC";
        ram_buffer(43483) := X"8FC401E8";
        ram_buffer(43484) := X"0C02EAF5";
        ram_buffer(43485) := X"00000000";
        ram_buffer(43486) := X"144000C9";
        ram_buffer(43487) := X"00000000";
        ram_buffer(43488) := X"27D000C4";
        ram_buffer(43489) := X"2631FFF0";
        ram_buffer(43490) := X"2A220011";
        ram_buffer(43491) := X"1040FFE1";
        ram_buffer(43492) := X"00000000";
        ram_buffer(43493) := X"3C02100D";
        ram_buffer(43494) := X"2442A8D0";
        ram_buffer(43495) := X"AE020000";
        ram_buffer(43496) := X"02201021";
        ram_buffer(43497) := X"AE020004";
        ram_buffer(43498) := X"8FC200C0";
        ram_buffer(43499) := X"02201821";
        ram_buffer(43500) := X"00431021";
        ram_buffer(43501) := X"AFC200C0";
        ram_buffer(43502) := X"26100008";
        ram_buffer(43503) := X"8FC200BC";
        ram_buffer(43504) := X"00000000";
        ram_buffer(43505) := X"24420001";
        ram_buffer(43506) := X"AFC200BC";
        ram_buffer(43507) := X"8FC200BC";
        ram_buffer(43508) := X"00000000";
        ram_buffer(43509) := X"28420008";
        ram_buffer(43510) := X"1440000A";
        ram_buffer(43511) := X"00000000";
        ram_buffer(43512) := X"27C200B8";
        ram_buffer(43513) := X"00403021";
        ram_buffer(43514) := X"8FC501EC";
        ram_buffer(43515) := X"8FC401E8";
        ram_buffer(43516) := X"0C02EAF5";
        ram_buffer(43517) := X"00000000";
        ram_buffer(43518) := X"144000AC";
        ram_buffer(43519) := X"00000000";
        ram_buffer(43520) := X"27D000C4";
        ram_buffer(43521) := X"8FC30034";
        ram_buffer(43522) := X"8FC20068";
        ram_buffer(43523) := X"00000000";
        ram_buffer(43524) := X"0043202A";
        ram_buffer(43525) := X"10800002";
        ram_buffer(43526) := X"00000000";
        ram_buffer(43527) := X"00601021";
        ram_buffer(43528) := X"8FC30030";
        ram_buffer(43529) := X"00000000";
        ram_buffer(43530) := X"00621021";
        ram_buffer(43531) := X"AFC20030";
        ram_buffer(43532) := X"8FC200C0";
        ram_buffer(43533) := X"00000000";
        ram_buffer(43534) := X"10400009";
        ram_buffer(43535) := X"00000000";
        ram_buffer(43536) := X"27C200B8";
        ram_buffer(43537) := X"00403021";
        ram_buffer(43538) := X"8FC501EC";
        ram_buffer(43539) := X"8FC401E8";
        ram_buffer(43540) := X"0C02EAF5";
        ram_buffer(43541) := X"00000000";
        ram_buffer(43542) := X"14400097";
        ram_buffer(43543) := X"00000000";
        ram_buffer(43544) := X"AFC000BC";
        ram_buffer(43545) := X"27D000C4";
        ram_buffer(43546) := X"8FC20074";
        ram_buffer(43547) := X"00000000";
        ram_buffer(43548) := X"1040F460";
        ram_buffer(43549) := X"00000000";
        ram_buffer(43550) := X"8FC50074";
        ram_buffer(43551) := X"8FC401E8";
        ram_buffer(43552) := X"0C027301";
        ram_buffer(43553) := X"00000000";
        ram_buffer(43554) := X"AFC00074";
        ram_buffer(43555) := X"1000F459";
        ram_buffer(43556) := X"00000000";
        ram_buffer(43557) := X"00000000";
        ram_buffer(43558) := X"10000002";
        ram_buffer(43559) := X"00000000";
        ram_buffer(43560) := X"00000000";
        ram_buffer(43561) := X"8FC200C0";
        ram_buffer(43562) := X"00000000";
        ram_buffer(43563) := X"10400009";
        ram_buffer(43564) := X"00000000";
        ram_buffer(43565) := X"27C200B8";
        ram_buffer(43566) := X"00403021";
        ram_buffer(43567) := X"8FC501EC";
        ram_buffer(43568) := X"8FC401E8";
        ram_buffer(43569) := X"0C02EAF5";
        ram_buffer(43570) := X"00000000";
        ram_buffer(43571) := X"1440007D";
        ram_buffer(43572) := X"00000000";
        ram_buffer(43573) := X"AFC000BC";
        ram_buffer(43574) := X"27D000C4";
        ram_buffer(43575) := X"1000007A";
        ram_buffer(43576) := X"00000000";
        ram_buffer(43577) := X"00000000";
        ram_buffer(43578) := X"10000077";
        ram_buffer(43579) := X"00000000";
        ram_buffer(43580) := X"00000000";
        ram_buffer(43581) := X"10000074";
        ram_buffer(43582) := X"00000000";
        ram_buffer(43583) := X"00000000";
        ram_buffer(43584) := X"10000071";
        ram_buffer(43585) := X"00000000";
        ram_buffer(43586) := X"00000000";
        ram_buffer(43587) := X"1000006E";
        ram_buffer(43588) := X"00000000";
        ram_buffer(43589) := X"00000000";
        ram_buffer(43590) := X"1000006B";
        ram_buffer(43591) := X"00000000";
        ram_buffer(43592) := X"00000000";
        ram_buffer(43593) := X"10000068";
        ram_buffer(43594) := X"00000000";
        ram_buffer(43595) := X"00000000";
        ram_buffer(43596) := X"10000065";
        ram_buffer(43597) := X"00000000";
        ram_buffer(43598) := X"00000000";
        ram_buffer(43599) := X"10000062";
        ram_buffer(43600) := X"00000000";
        ram_buffer(43601) := X"00000000";
        ram_buffer(43602) := X"1000005F";
        ram_buffer(43603) := X"00000000";
        ram_buffer(43604) := X"00000000";
        ram_buffer(43605) := X"1000005C";
        ram_buffer(43606) := X"00000000";
        ram_buffer(43607) := X"00000000";
        ram_buffer(43608) := X"10000059";
        ram_buffer(43609) := X"00000000";
        ram_buffer(43610) := X"00000000";
        ram_buffer(43611) := X"10000056";
        ram_buffer(43612) := X"00000000";
        ram_buffer(43613) := X"00000000";
        ram_buffer(43614) := X"10000053";
        ram_buffer(43615) := X"00000000";
        ram_buffer(43616) := X"00000000";
        ram_buffer(43617) := X"10000050";
        ram_buffer(43618) := X"00000000";
        ram_buffer(43619) := X"00000000";
        ram_buffer(43620) := X"1000004D";
        ram_buffer(43621) := X"00000000";
        ram_buffer(43622) := X"00000000";
        ram_buffer(43623) := X"1000004A";
        ram_buffer(43624) := X"00000000";
        ram_buffer(43625) := X"00000000";
        ram_buffer(43626) := X"10000047";
        ram_buffer(43627) := X"00000000";
        ram_buffer(43628) := X"00000000";
        ram_buffer(43629) := X"10000044";
        ram_buffer(43630) := X"00000000";
        ram_buffer(43631) := X"00000000";
        ram_buffer(43632) := X"10000041";
        ram_buffer(43633) := X"00000000";
        ram_buffer(43634) := X"00000000";
        ram_buffer(43635) := X"1000003E";
        ram_buffer(43636) := X"00000000";
        ram_buffer(43637) := X"00000000";
        ram_buffer(43638) := X"1000003B";
        ram_buffer(43639) := X"00000000";
        ram_buffer(43640) := X"00000000";
        ram_buffer(43641) := X"10000038";
        ram_buffer(43642) := X"00000000";
        ram_buffer(43643) := X"00000000";
        ram_buffer(43644) := X"10000035";
        ram_buffer(43645) := X"00000000";
        ram_buffer(43646) := X"00000000";
        ram_buffer(43647) := X"10000032";
        ram_buffer(43648) := X"00000000";
        ram_buffer(43649) := X"00000000";
        ram_buffer(43650) := X"1000002F";
        ram_buffer(43651) := X"00000000";
        ram_buffer(43652) := X"00000000";
        ram_buffer(43653) := X"1000002C";
        ram_buffer(43654) := X"00000000";
        ram_buffer(43655) := X"00000000";
        ram_buffer(43656) := X"10000029";
        ram_buffer(43657) := X"00000000";
        ram_buffer(43658) := X"00000000";
        ram_buffer(43659) := X"10000026";
        ram_buffer(43660) := X"00000000";
        ram_buffer(43661) := X"00000000";
        ram_buffer(43662) := X"10000023";
        ram_buffer(43663) := X"00000000";
        ram_buffer(43664) := X"00000000";
        ram_buffer(43665) := X"10000020";
        ram_buffer(43666) := X"00000000";
        ram_buffer(43667) := X"00000000";
        ram_buffer(43668) := X"1000001D";
        ram_buffer(43669) := X"00000000";
        ram_buffer(43670) := X"00000000";
        ram_buffer(43671) := X"1000001A";
        ram_buffer(43672) := X"00000000";
        ram_buffer(43673) := X"00000000";
        ram_buffer(43674) := X"10000017";
        ram_buffer(43675) := X"00000000";
        ram_buffer(43676) := X"00000000";
        ram_buffer(43677) := X"10000014";
        ram_buffer(43678) := X"00000000";
        ram_buffer(43679) := X"00000000";
        ram_buffer(43680) := X"10000011";
        ram_buffer(43681) := X"00000000";
        ram_buffer(43682) := X"00000000";
        ram_buffer(43683) := X"1000000E";
        ram_buffer(43684) := X"00000000";
        ram_buffer(43685) := X"00000000";
        ram_buffer(43686) := X"1000000B";
        ram_buffer(43687) := X"00000000";
        ram_buffer(43688) := X"00000000";
        ram_buffer(43689) := X"10000008";
        ram_buffer(43690) := X"00000000";
        ram_buffer(43691) := X"00000000";
        ram_buffer(43692) := X"10000005";
        ram_buffer(43693) := X"00000000";
        ram_buffer(43694) := X"00000000";
        ram_buffer(43695) := X"10000002";
        ram_buffer(43696) := X"00000000";
        ram_buffer(43697) := X"00000000";
        ram_buffer(43698) := X"8FC20074";
        ram_buffer(43699) := X"00000000";
        ram_buffer(43700) := X"10400005";
        ram_buffer(43701) := X"00000000";
        ram_buffer(43702) := X"8FC50074";
        ram_buffer(43703) := X"8FC401E8";
        ram_buffer(43704) := X"0C027301";
        ram_buffer(43705) := X"00000000";
        ram_buffer(43706) := X"8FC201EC";
        ram_buffer(43707) := X"00000000";
        ram_buffer(43708) := X"8442000C";
        ram_buffer(43709) := X"00000000";
        ram_buffer(43710) := X"3042FFFF";
        ram_buffer(43711) := X"30420040";
        ram_buffer(43712) := X"14400004";
        ram_buffer(43713) := X"00000000";
        ram_buffer(43714) := X"8FC20030";
        ram_buffer(43715) := X"10000003";
        ram_buffer(43716) := X"00000000";
        ram_buffer(43717) := X"2402FFFF";
        ram_buffer(43718) := X"00000000";
        ram_buffer(43719) := X"03C0E821";
        ram_buffer(43720) := X"8FBF01E4";
        ram_buffer(43721) := X"8FBE01E0";
        ram_buffer(43722) := X"8FB701DC";
        ram_buffer(43723) := X"8FB601D8";
        ram_buffer(43724) := X"8FB501D4";
        ram_buffer(43725) := X"8FB401D0";
        ram_buffer(43726) := X"8FB301CC";
        ram_buffer(43727) := X"8FB201C8";
        ram_buffer(43728) := X"8FB101C4";
        ram_buffer(43729) := X"8FB001C0";
        ram_buffer(43730) := X"27BD01E8";
        ram_buffer(43731) := X"03E00008";
        ram_buffer(43732) := X"00000000";
        ram_buffer(43733) := X"27BDFFB0";
        ram_buffer(43734) := X"AFBF004C";
        ram_buffer(43735) := X"AFBE0048";
        ram_buffer(43736) := X"03A0F021";
        ram_buffer(43737) := X"AFC40050";
        ram_buffer(43738) := X"AFC7005C";
        ram_buffer(43739) := X"AFC60058";
        ram_buffer(43740) := X"8FC3005C";
        ram_buffer(43741) := X"8FC20058";
        ram_buffer(43742) := X"AFC30044";
        ram_buffer(43743) := X"AFC20040";
        ram_buffer(43744) := X"8FC20040";
        ram_buffer(43745) := X"00000000";
        ram_buffer(43746) := X"0441000D";
        ram_buffer(43747) := X"00000000";
        ram_buffer(43748) := X"8FC30058";
        ram_buffer(43749) := X"3C028000";
        ram_buffer(43750) := X"00621026";
        ram_buffer(43751) := X"AFC20058";
        ram_buffer(43752) := X"8FC2005C";
        ram_buffer(43753) := X"00000000";
        ram_buffer(43754) := X"AFC2005C";
        ram_buffer(43755) := X"8FC20068";
        ram_buffer(43756) := X"2403002D";
        ram_buffer(43757) := X"A0430000";
        ram_buffer(43758) := X"10000004";
        ram_buffer(43759) := X"00000000";
        ram_buffer(43760) := X"8FC20068";
        ram_buffer(43761) := X"00000000";
        ram_buffer(43762) := X"A0400000";
        ram_buffer(43763) := X"8FC30070";
        ram_buffer(43764) := X"24020061";
        ram_buffer(43765) := X"10620005";
        ram_buffer(43766) := X"00000000";
        ram_buffer(43767) := X"8FC30070";
        ram_buffer(43768) := X"24020041";
        ram_buffer(43769) := X"146200B3";
        ram_buffer(43770) := X"00000000";
        ram_buffer(43771) := X"8FC6006C";
        ram_buffer(43772) := X"8FC5005C";
        ram_buffer(43773) := X"8FC40058";
        ram_buffer(43774) := X"0C02CB50";
        ram_buffer(43775) := X"00000000";
        ram_buffer(43776) := X"8F8780C4";
        ram_buffer(43777) := X"8F8680C0";
        ram_buffer(43778) := X"00602821";
        ram_buffer(43779) := X"00402021";
        ram_buffer(43780) := X"0C03144F";
        ram_buffer(43781) := X"00000000";
        ram_buffer(43782) := X"AFC3005C";
        ram_buffer(43783) := X"AFC20058";
        ram_buffer(43784) := X"00003821";
        ram_buffer(43785) := X"00003021";
        ram_buffer(43786) := X"8FC5005C";
        ram_buffer(43787) := X"8FC40058";
        ram_buffer(43788) := X"0C03167F";
        ram_buffer(43789) := X"00000000";
        ram_buffer(43790) := X"14400004";
        ram_buffer(43791) := X"00000000";
        ram_buffer(43792) := X"8FC2006C";
        ram_buffer(43793) := X"24030001";
        ram_buffer(43794) := X"AC430000";
        ram_buffer(43795) := X"8FC30070";
        ram_buffer(43796) := X"24020061";
        ram_buffer(43797) := X"14620005";
        ram_buffer(43798) := X"00000000";
        ram_buffer(43799) := X"3C02100D";
        ram_buffer(43800) := X"2442A714";
        ram_buffer(43801) := X"10000003";
        ram_buffer(43802) := X"00000000";
        ram_buffer(43803) := X"3C02100D";
        ram_buffer(43804) := X"2442A730";
        ram_buffer(43805) := X"AFC20030";
        ram_buffer(43806) := X"8FC20078";
        ram_buffer(43807) := X"00000000";
        ram_buffer(43808) := X"AFC2002C";
        ram_buffer(43809) := X"8F8780CC";
        ram_buffer(43810) := X"8F8680C8";
        ram_buffer(43811) := X"8FC5005C";
        ram_buffer(43812) := X"8FC40058";
        ram_buffer(43813) := X"0C03174A";
        ram_buffer(43814) := X"00000000";
        ram_buffer(43815) := X"AFC3005C";
        ram_buffer(43816) := X"AFC20058";
        ram_buffer(43817) := X"8FC5005C";
        ram_buffer(43818) := X"8FC40058";
        ram_buffer(43819) := X"0C031B37";
        ram_buffer(43820) := X"00000000";
        ram_buffer(43821) := X"AFC20028";
        ram_buffer(43822) := X"8FC40028";
        ram_buffer(43823) := X"0C031B7C";
        ram_buffer(43824) := X"00000000";
        ram_buffer(43825) := X"00603821";
        ram_buffer(43826) := X"00403021";
        ram_buffer(43827) := X"8FC5005C";
        ram_buffer(43828) := X"8FC40058";
        ram_buffer(43829) := X"0C0318D3";
        ram_buffer(43830) := X"00000000";
        ram_buffer(43831) := X"AFC3005C";
        ram_buffer(43832) := X"AFC20058";
        ram_buffer(43833) := X"8FC2002C";
        ram_buffer(43834) := X"00000000";
        ram_buffer(43835) := X"24430001";
        ram_buffer(43836) := X"AFC3002C";
        ram_buffer(43837) := X"8FC30028";
        ram_buffer(43838) := X"8FC40030";
        ram_buffer(43839) := X"00000000";
        ram_buffer(43840) := X"00831821";
        ram_buffer(43841) := X"80630000";
        ram_buffer(43842) := X"00000000";
        ram_buffer(43843) := X"A0430000";
        ram_buffer(43844) := X"8FC20060";
        ram_buffer(43845) := X"00000000";
        ram_buffer(43846) := X"2443FFFF";
        ram_buffer(43847) := X"AFC30060";
        ram_buffer(43848) := X"10400009";
        ram_buffer(43849) := X"00000000";
        ram_buffer(43850) := X"00003821";
        ram_buffer(43851) := X"00003021";
        ram_buffer(43852) := X"8FC5005C";
        ram_buffer(43853) := X"8FC40058";
        ram_buffer(43854) := X"0C03167F";
        ram_buffer(43855) := X"00000000";
        ram_buffer(43856) := X"1440FFD0";
        ram_buffer(43857) := X"00000000";
        ram_buffer(43858) := X"8F8780D4";
        ram_buffer(43859) := X"8F8680D0";
        ram_buffer(43860) := X"8FC5005C";
        ram_buffer(43861) := X"8FC40058";
        ram_buffer(43862) := X"0C0316AB";
        ram_buffer(43863) := X"00000000";
        ram_buffer(43864) := X"1C40000E";
        ram_buffer(43865) := X"00000000";
        ram_buffer(43866) := X"8F8780D4";
        ram_buffer(43867) := X"8F8680D0";
        ram_buffer(43868) := X"8FC5005C";
        ram_buffer(43869) := X"8FC40058";
        ram_buffer(43870) := X"0C03167F";
        ram_buffer(43871) := X"00000000";
        ram_buffer(43872) := X"14400034";
        ram_buffer(43873) := X"00000000";
        ram_buffer(43874) := X"8FC20028";
        ram_buffer(43875) := X"00000000";
        ram_buffer(43876) := X"30420001";
        ram_buffer(43877) := X"10400037";
        ram_buffer(43878) := X"00000000";
        ram_buffer(43879) := X"8FC2002C";
        ram_buffer(43880) := X"00000000";
        ram_buffer(43881) := X"AFC20038";
        ram_buffer(43882) := X"10000004";
        ram_buffer(43883) := X"00000000";
        ram_buffer(43884) := X"8FC20038";
        ram_buffer(43885) := X"24030030";
        ram_buffer(43886) := X"A0430000";
        ram_buffer(43887) := X"8FC20038";
        ram_buffer(43888) := X"00000000";
        ram_buffer(43889) := X"2442FFFF";
        ram_buffer(43890) := X"AFC20038";
        ram_buffer(43891) := X"8FC20038";
        ram_buffer(43892) := X"00000000";
        ram_buffer(43893) := X"80430000";
        ram_buffer(43894) := X"8FC20030";
        ram_buffer(43895) := X"00000000";
        ram_buffer(43896) := X"2442000F";
        ram_buffer(43897) := X"80420000";
        ram_buffer(43898) := X"00000000";
        ram_buffer(43899) := X"1062FFF0";
        ram_buffer(43900) := X"00000000";
        ram_buffer(43901) := X"8FC30038";
        ram_buffer(43902) := X"8FC20038";
        ram_buffer(43903) := X"00000000";
        ram_buffer(43904) := X"80440000";
        ram_buffer(43905) := X"24020039";
        ram_buffer(43906) := X"14820006";
        ram_buffer(43907) := X"00000000";
        ram_buffer(43908) := X"8FC20030";
        ram_buffer(43909) := X"00000000";
        ram_buffer(43910) := X"8042000A";
        ram_buffer(43911) := X"1000000A";
        ram_buffer(43912) := X"00000000";
        ram_buffer(43913) := X"8FC20038";
        ram_buffer(43914) := X"00000000";
        ram_buffer(43915) := X"80420000";
        ram_buffer(43916) := X"00000000";
        ram_buffer(43917) := X"304200FF";
        ram_buffer(43918) := X"24420001";
        ram_buffer(43919) := X"304200FF";
        ram_buffer(43920) := X"00021600";
        ram_buffer(43921) := X"00021603";
        ram_buffer(43922) := X"A0620000";
        ram_buffer(43923) := X"1000000F";
        ram_buffer(43924) := X"00000000";
        ram_buffer(43925) := X"10000007";
        ram_buffer(43926) := X"00000000";
        ram_buffer(43927) := X"8FC2002C";
        ram_buffer(43928) := X"00000000";
        ram_buffer(43929) := X"24430001";
        ram_buffer(43930) := X"AFC3002C";
        ram_buffer(43931) := X"24030030";
        ram_buffer(43932) := X"A0430000";
        ram_buffer(43933) := X"8FC20060";
        ram_buffer(43934) := X"00000000";
        ram_buffer(43935) := X"2443FFFF";
        ram_buffer(43936) := X"AFC30060";
        ram_buffer(43937) := X"0441FFF5";
        ram_buffer(43938) := X"00000000";
        ram_buffer(43939) := X"8FC3002C";
        ram_buffer(43940) := X"8FC20078";
        ram_buffer(43941) := X"00000000";
        ram_buffer(43942) := X"00621823";
        ram_buffer(43943) := X"8FC20074";
        ram_buffer(43944) := X"00000000";
        ram_buffer(43945) := X"AC430000";
        ram_buffer(43946) := X"8FC20078";
        ram_buffer(43947) := X"10000089";
        ram_buffer(43948) := X"00000000";
        ram_buffer(43949) := X"8FC30070";
        ram_buffer(43950) := X"24020066";
        ram_buffer(43951) := X"10620005";
        ram_buffer(43952) := X"00000000";
        ram_buffer(43953) := X"8FC30070";
        ram_buffer(43954) := X"24020046";
        ram_buffer(43955) := X"14620005";
        ram_buffer(43956) := X"00000000";
        ram_buffer(43957) := X"24020003";
        ram_buffer(43958) := X"AFC20028";
        ram_buffer(43959) := X"1000000F";
        ram_buffer(43960) := X"00000000";
        ram_buffer(43961) := X"8FC30070";
        ram_buffer(43962) := X"24020065";
        ram_buffer(43963) := X"10620005";
        ram_buffer(43964) := X"00000000";
        ram_buffer(43965) := X"8FC30070";
        ram_buffer(43966) := X"24020045";
        ram_buffer(43967) := X"14620005";
        ram_buffer(43968) := X"00000000";
        ram_buffer(43969) := X"8FC20060";
        ram_buffer(43970) := X"00000000";
        ram_buffer(43971) := X"24420001";
        ram_buffer(43972) := X"AFC20060";
        ram_buffer(43973) := X"24020002";
        ram_buffer(43974) := X"AFC20028";
        ram_buffer(43975) := X"27C20038";
        ram_buffer(43976) := X"AFA20020";
        ram_buffer(43977) := X"27C20034";
        ram_buffer(43978) := X"AFA2001C";
        ram_buffer(43979) := X"8FC2006C";
        ram_buffer(43980) := X"00000000";
        ram_buffer(43981) := X"AFA20018";
        ram_buffer(43982) := X"8FC20060";
        ram_buffer(43983) := X"00000000";
        ram_buffer(43984) := X"AFA20014";
        ram_buffer(43985) := X"8FC20028";
        ram_buffer(43986) := X"00000000";
        ram_buffer(43987) := X"AFA20010";
        ram_buffer(43988) := X"8FC7005C";
        ram_buffer(43989) := X"8FC60058";
        ram_buffer(43990) := X"8FC40050";
        ram_buffer(43991) := X"0C02AFA3";
        ram_buffer(43992) := X"00000000";
        ram_buffer(43993) := X"AFC20030";
        ram_buffer(43994) := X"8FC30070";
        ram_buffer(43995) := X"24020067";
        ram_buffer(43996) := X"10620005";
        ram_buffer(43997) := X"00000000";
        ram_buffer(43998) := X"8FC30070";
        ram_buffer(43999) := X"24020047";
        ram_buffer(44000) := X"14620006";
        ram_buffer(44001) := X"00000000";
        ram_buffer(44002) := X"8FC20064";
        ram_buffer(44003) := X"00000000";
        ram_buffer(44004) := X"30420001";
        ram_buffer(44005) := X"10400045";
        ram_buffer(44006) := X"00000000";
        ram_buffer(44007) := X"8FC20060";
        ram_buffer(44008) := X"8FC30030";
        ram_buffer(44009) := X"00000000";
        ram_buffer(44010) := X"00621021";
        ram_buffer(44011) := X"AFC2002C";
        ram_buffer(44012) := X"8FC30070";
        ram_buffer(44013) := X"24020066";
        ram_buffer(44014) := X"10620005";
        ram_buffer(44015) := X"00000000";
        ram_buffer(44016) := X"8FC30070";
        ram_buffer(44017) := X"24020046";
        ram_buffer(44018) := X"1462001F";
        ram_buffer(44019) := X"00000000";
        ram_buffer(44020) := X"8FC20030";
        ram_buffer(44021) := X"00000000";
        ram_buffer(44022) := X"80430000";
        ram_buffer(44023) := X"24020030";
        ram_buffer(44024) := X"14620010";
        ram_buffer(44025) := X"00000000";
        ram_buffer(44026) := X"00003821";
        ram_buffer(44027) := X"00003021";
        ram_buffer(44028) := X"8FC5005C";
        ram_buffer(44029) := X"8FC40058";
        ram_buffer(44030) := X"0C03167F";
        ram_buffer(44031) := X"00000000";
        ram_buffer(44032) := X"10400008";
        ram_buffer(44033) := X"00000000";
        ram_buffer(44034) := X"24030001";
        ram_buffer(44035) := X"8FC20060";
        ram_buffer(44036) := X"00000000";
        ram_buffer(44037) := X"00621823";
        ram_buffer(44038) := X"8FC2006C";
        ram_buffer(44039) := X"00000000";
        ram_buffer(44040) := X"AC430000";
        ram_buffer(44041) := X"8FC2006C";
        ram_buffer(44042) := X"00000000";
        ram_buffer(44043) := X"8C420000";
        ram_buffer(44044) := X"00000000";
        ram_buffer(44045) := X"00401821";
        ram_buffer(44046) := X"8FC2002C";
        ram_buffer(44047) := X"00000000";
        ram_buffer(44048) := X"00431021";
        ram_buffer(44049) := X"AFC2002C";
        ram_buffer(44050) := X"00003821";
        ram_buffer(44051) := X"00003021";
        ram_buffer(44052) := X"8FC5005C";
        ram_buffer(44053) := X"8FC40058";
        ram_buffer(44054) := X"0C03167F";
        ram_buffer(44055) := X"00000000";
        ram_buffer(44056) := X"14400004";
        ram_buffer(44057) := X"00000000";
        ram_buffer(44058) := X"8FC2002C";
        ram_buffer(44059) := X"00000000";
        ram_buffer(44060) := X"AFC20038";
        ram_buffer(44061) := X"10000007";
        ram_buffer(44062) := X"00000000";
        ram_buffer(44063) := X"8FC20038";
        ram_buffer(44064) := X"00000000";
        ram_buffer(44065) := X"24430001";
        ram_buffer(44066) := X"AFC30038";
        ram_buffer(44067) := X"24030030";
        ram_buffer(44068) := X"A0430000";
        ram_buffer(44069) := X"8FC30038";
        ram_buffer(44070) := X"8FC2002C";
        ram_buffer(44071) := X"00000000";
        ram_buffer(44072) := X"0062102B";
        ram_buffer(44073) := X"1440FFF5";
        ram_buffer(44074) := X"00000000";
        ram_buffer(44075) := X"8FC20038";
        ram_buffer(44076) := X"00000000";
        ram_buffer(44077) := X"00401821";
        ram_buffer(44078) := X"8FC20030";
        ram_buffer(44079) := X"00000000";
        ram_buffer(44080) := X"00621823";
        ram_buffer(44081) := X"8FC20074";
        ram_buffer(44082) := X"00000000";
        ram_buffer(44083) := X"AC430000";
        ram_buffer(44084) := X"8FC20030";
        ram_buffer(44085) := X"03C0E821";
        ram_buffer(44086) := X"8FBF004C";
        ram_buffer(44087) := X"8FBE0048";
        ram_buffer(44088) := X"27BD0050";
        ram_buffer(44089) := X"03E00008";
        ram_buffer(44090) := X"00000000";
        ram_buffer(44091) := X"27BDFFE0";
        ram_buffer(44092) := X"AFBE001C";
        ram_buffer(44093) := X"AFB10018";
        ram_buffer(44094) := X"AFB00014";
        ram_buffer(44095) := X"03A0F021";
        ram_buffer(44096) := X"AFC40020";
        ram_buffer(44097) := X"AFC50024";
        ram_buffer(44098) := X"AFC60028";
        ram_buffer(44099) := X"8FC30028";
        ram_buffer(44100) := X"24020061";
        ram_buffer(44101) := X"10620005";
        ram_buffer(44102) := X"00000000";
        ram_buffer(44103) := X"8FC30028";
        ram_buffer(44104) := X"24020041";
        ram_buffer(44105) := X"14620004";
        ram_buffer(44106) := X"00000000";
        ram_buffer(44107) := X"24020001";
        ram_buffer(44108) := X"10000002";
        ram_buffer(44109) := X"00000000";
        ram_buffer(44110) := X"00001021";
        ram_buffer(44111) := X"AFC20000";
        ram_buffer(44112) := X"8FD10020";
        ram_buffer(44113) := X"00000000";
        ram_buffer(44114) := X"02201821";
        ram_buffer(44115) := X"24710001";
        ram_buffer(44116) := X"8FC20000";
        ram_buffer(44117) := X"00000000";
        ram_buffer(44118) := X"1040000A";
        ram_buffer(44119) := X"00000000";
        ram_buffer(44120) := X"8FC20028";
        ram_buffer(44121) := X"00000000";
        ram_buffer(44122) := X"304200FF";
        ram_buffer(44123) := X"2442000F";
        ram_buffer(44124) := X"304200FF";
        ram_buffer(44125) := X"00021600";
        ram_buffer(44126) := X"00021603";
        ram_buffer(44127) := X"10000005";
        ram_buffer(44128) := X"00000000";
        ram_buffer(44129) := X"8FC20028";
        ram_buffer(44130) := X"00000000";
        ram_buffer(44131) := X"00021600";
        ram_buffer(44132) := X"00021603";
        ram_buffer(44133) := X"A0620000";
        ram_buffer(44134) := X"8FC20024";
        ram_buffer(44135) := X"00000000";
        ram_buffer(44136) := X"0441000B";
        ram_buffer(44137) := X"00000000";
        ram_buffer(44138) := X"8FC20024";
        ram_buffer(44139) := X"00000000";
        ram_buffer(44140) := X"00021023";
        ram_buffer(44141) := X"AFC20024";
        ram_buffer(44142) := X"02201021";
        ram_buffer(44143) := X"24510001";
        ram_buffer(44144) := X"2403002D";
        ram_buffer(44145) := X"A0430000";
        ram_buffer(44146) := X"10000005";
        ram_buffer(44147) := X"00000000";
        ram_buffer(44148) := X"02201021";
        ram_buffer(44149) := X"24510001";
        ram_buffer(44150) := X"2403002B";
        ram_buffer(44151) := X"A0430000";
        ram_buffer(44152) := X"27D00004";
        ram_buffer(44153) := X"26100007";
        ram_buffer(44154) := X"8FC20024";
        ram_buffer(44155) := X"00000000";
        ram_buffer(44156) := X"2842000A";
        ram_buffer(44157) := X"14400034";
        ram_buffer(44158) := X"00000000";
        ram_buffer(44159) := X"2610FFFF";
        ram_buffer(44160) := X"8FC30024";
        ram_buffer(44161) := X"2402000A";
        ram_buffer(44162) := X"14400002";
        ram_buffer(44163) := X"0062001A";
        ram_buffer(44164) := X"0007000D";
        ram_buffer(44165) := X"00001010";
        ram_buffer(44166) := X"304200FF";
        ram_buffer(44167) := X"24420030";
        ram_buffer(44168) := X"304200FF";
        ram_buffer(44169) := X"00021600";
        ram_buffer(44170) := X"00021603";
        ram_buffer(44171) := X"A2020000";
        ram_buffer(44172) := X"8FC30024";
        ram_buffer(44173) := X"2402000A";
        ram_buffer(44174) := X"14400002";
        ram_buffer(44175) := X"0062001A";
        ram_buffer(44176) := X"0007000D";
        ram_buffer(44177) := X"00001010";
        ram_buffer(44178) := X"00001012";
        ram_buffer(44179) := X"AFC20024";
        ram_buffer(44180) := X"8FC20024";
        ram_buffer(44181) := X"00000000";
        ram_buffer(44182) := X"2842000A";
        ram_buffer(44183) := X"1040FFE7";
        ram_buffer(44184) := X"00000000";
        ram_buffer(44185) := X"2610FFFF";
        ram_buffer(44186) := X"8FC20024";
        ram_buffer(44187) := X"00000000";
        ram_buffer(44188) := X"304200FF";
        ram_buffer(44189) := X"24420030";
        ram_buffer(44190) := X"304200FF";
        ram_buffer(44191) := X"00021600";
        ram_buffer(44192) := X"00021603";
        ram_buffer(44193) := X"A2020000";
        ram_buffer(44194) := X"10000008";
        ram_buffer(44195) := X"00000000";
        ram_buffer(44196) := X"02201021";
        ram_buffer(44197) := X"24510001";
        ram_buffer(44198) := X"02001821";
        ram_buffer(44199) := X"24700001";
        ram_buffer(44200) := X"80630000";
        ram_buffer(44201) := X"00000000";
        ram_buffer(44202) := X"A0430000";
        ram_buffer(44203) := X"27C20004";
        ram_buffer(44204) := X"24420007";
        ram_buffer(44205) := X"0202102B";
        ram_buffer(44206) := X"1440FFF5";
        ram_buffer(44207) := X"00000000";
        ram_buffer(44208) := X"10000013";
        ram_buffer(44209) := X"00000000";
        ram_buffer(44210) := X"8FC20000";
        ram_buffer(44211) := X"00000000";
        ram_buffer(44212) := X"14400005";
        ram_buffer(44213) := X"00000000";
        ram_buffer(44214) := X"02201021";
        ram_buffer(44215) := X"24510001";
        ram_buffer(44216) := X"24030030";
        ram_buffer(44217) := X"A0430000";
        ram_buffer(44218) := X"02201021";
        ram_buffer(44219) := X"24510001";
        ram_buffer(44220) := X"8FC30024";
        ram_buffer(44221) := X"00000000";
        ram_buffer(44222) := X"306300FF";
        ram_buffer(44223) := X"24630030";
        ram_buffer(44224) := X"306300FF";
        ram_buffer(44225) := X"00031E00";
        ram_buffer(44226) := X"00031E03";
        ram_buffer(44227) := X"A0430000";
        ram_buffer(44228) := X"02201821";
        ram_buffer(44229) := X"8FC20020";
        ram_buffer(44230) := X"00000000";
        ram_buffer(44231) := X"00621023";
        ram_buffer(44232) := X"03C0E821";
        ram_buffer(44233) := X"8FBE001C";
        ram_buffer(44234) := X"8FB10018";
        ram_buffer(44235) := X"8FB00014";
        ram_buffer(44236) := X"27BD0020";
        ram_buffer(44237) := X"03E00008";
        ram_buffer(44238) := X"00000000";
        ram_buffer(44239) := X"27BDFFE0";
        ram_buffer(44240) := X"AFBF001C";
        ram_buffer(44241) := X"AFBE0018";
        ram_buffer(44242) := X"03A0F021";
        ram_buffer(44243) := X"AFC40020";
        ram_buffer(44244) := X"AFC50024";
        ram_buffer(44245) := X"AFC60028";
        ram_buffer(44246) := X"AFC7002C";
        ram_buffer(44247) := X"AF8081EC";
        ram_buffer(44248) := X"8FC6002C";
        ram_buffer(44249) := X"8FC50028";
        ram_buffer(44250) := X"8FC40024";
        ram_buffer(44251) := X"0C02FCE3";
        ram_buffer(44252) := X"00000000";
        ram_buffer(44253) := X"AFC20010";
        ram_buffer(44254) := X"8FC30010";
        ram_buffer(44255) := X"2402FFFF";
        ram_buffer(44256) := X"14620009";
        ram_buffer(44257) := X"00000000";
        ram_buffer(44258) := X"8F8281EC";
        ram_buffer(44259) := X"00000000";
        ram_buffer(44260) := X"10400005";
        ram_buffer(44261) := X"00000000";
        ram_buffer(44262) := X"8F8381EC";
        ram_buffer(44263) := X"8FC20020";
        ram_buffer(44264) := X"00000000";
        ram_buffer(44265) := X"AC430000";
        ram_buffer(44266) := X"8FC20010";
        ram_buffer(44267) := X"03C0E821";
        ram_buffer(44268) := X"8FBF001C";
        ram_buffer(44269) := X"8FBE0018";
        ram_buffer(44270) := X"27BD0020";
        ram_buffer(44271) := X"03E00008";
        ram_buffer(44272) := X"00000000";
        ram_buffer(44273) := X"27BDFFD8";
        ram_buffer(44274) := X"AFBF0024";
        ram_buffer(44275) := X"AFBE0020";
        ram_buffer(44276) := X"AFB0001C";
        ram_buffer(44277) := X"03A0F021";
        ram_buffer(44278) := X"AFC40028";
        ram_buffer(44279) := X"00A08021";
        ram_buffer(44280) := X"8F828098";
        ram_buffer(44281) := X"00000000";
        ram_buffer(44282) := X"AFC20010";
        ram_buffer(44283) := X"8FC20010";
        ram_buffer(44284) := X"00000000";
        ram_buffer(44285) := X"1040000A";
        ram_buffer(44286) := X"00000000";
        ram_buffer(44287) := X"8FC20010";
        ram_buffer(44288) := X"00000000";
        ram_buffer(44289) := X"8C420038";
        ram_buffer(44290) := X"00000000";
        ram_buffer(44291) := X"14400004";
        ram_buffer(44292) := X"00000000";
        ram_buffer(44293) := X"8FC40010";
        ram_buffer(44294) := X"0C027069";
        ram_buffer(44295) := X"00000000";
        ram_buffer(44296) := X"8602000C";
        ram_buffer(44297) := X"00000000";
        ram_buffer(44298) := X"3042FFFF";
        ram_buffer(44299) := X"30420008";
        ram_buffer(44300) := X"14400038";
        ram_buffer(44301) := X"00000000";
        ram_buffer(44302) := X"8602000C";
        ram_buffer(44303) := X"00000000";
        ram_buffer(44304) := X"3042FFFF";
        ram_buffer(44305) := X"30420010";
        ram_buffer(44306) := X"1440000D";
        ram_buffer(44307) := X"00000000";
        ram_buffer(44308) := X"8FC20028";
        ram_buffer(44309) := X"24030009";
        ram_buffer(44310) := X"AC430000";
        ram_buffer(44311) := X"8602000C";
        ram_buffer(44312) := X"00000000";
        ram_buffer(44313) := X"34420040";
        ram_buffer(44314) := X"00021400";
        ram_buffer(44315) := X"00021403";
        ram_buffer(44316) := X"A602000C";
        ram_buffer(44317) := X"2402FFFF";
        ram_buffer(44318) := X"10000066";
        ram_buffer(44319) := X"00000000";
        ram_buffer(44320) := X"8602000C";
        ram_buffer(44321) := X"00000000";
        ram_buffer(44322) := X"3042FFFF";
        ram_buffer(44323) := X"30420004";
        ram_buffer(44324) := X"1040001A";
        ram_buffer(44325) := X"00000000";
        ram_buffer(44326) := X"8E020030";
        ram_buffer(44327) := X"00000000";
        ram_buffer(44328) := X"1040000C";
        ram_buffer(44329) := X"00000000";
        ram_buffer(44330) := X"8E030030";
        ram_buffer(44331) := X"26020040";
        ram_buffer(44332) := X"10620007";
        ram_buffer(44333) := X"00000000";
        ram_buffer(44334) := X"8E020030";
        ram_buffer(44335) := X"00000000";
        ram_buffer(44336) := X"00402821";
        ram_buffer(44337) := X"8FC40028";
        ram_buffer(44338) := X"0C027301";
        ram_buffer(44339) := X"00000000";
        ram_buffer(44340) := X"AE000030";
        ram_buffer(44341) := X"8603000C";
        ram_buffer(44342) := X"2402FFDB";
        ram_buffer(44343) := X"00621024";
        ram_buffer(44344) := X"00021400";
        ram_buffer(44345) := X"00021403";
        ram_buffer(44346) := X"A602000C";
        ram_buffer(44347) := X"AE000004";
        ram_buffer(44348) := X"8E020010";
        ram_buffer(44349) := X"00000000";
        ram_buffer(44350) := X"AE020000";
        ram_buffer(44351) := X"8602000C";
        ram_buffer(44352) := X"00000000";
        ram_buffer(44353) := X"34420008";
        ram_buffer(44354) := X"00021400";
        ram_buffer(44355) := X"00021403";
        ram_buffer(44356) := X"A602000C";
        ram_buffer(44357) := X"8E020010";
        ram_buffer(44358) := X"00000000";
        ram_buffer(44359) := X"14400011";
        ram_buffer(44360) := X"00000000";
        ram_buffer(44361) := X"8602000C";
        ram_buffer(44362) := X"00000000";
        ram_buffer(44363) := X"3042FFFF";
        ram_buffer(44364) := X"30420200";
        ram_buffer(44365) := X"10400007";
        ram_buffer(44366) := X"00000000";
        ram_buffer(44367) := X"8602000C";
        ram_buffer(44368) := X"00000000";
        ram_buffer(44369) := X"3042FFFF";
        ram_buffer(44370) := X"30420080";
        ram_buffer(44371) := X"10400005";
        ram_buffer(44372) := X"00000000";
        ram_buffer(44373) := X"02002821";
        ram_buffer(44374) := X"8FC40028";
        ram_buffer(44375) := X"0C027999";
        ram_buffer(44376) := X"00000000";
        ram_buffer(44377) := X"8602000C";
        ram_buffer(44378) := X"00000000";
        ram_buffer(44379) := X"3042FFFF";
        ram_buffer(44380) := X"30420001";
        ram_buffer(44381) := X"10400008";
        ram_buffer(44382) := X"00000000";
        ram_buffer(44383) := X"AE000008";
        ram_buffer(44384) := X"8E020014";
        ram_buffer(44385) := X"00000000";
        ram_buffer(44386) := X"00021023";
        ram_buffer(44387) := X"AE020018";
        ram_buffer(44388) := X"1000000C";
        ram_buffer(44389) := X"00000000";
        ram_buffer(44390) := X"8602000C";
        ram_buffer(44391) := X"00000000";
        ram_buffer(44392) := X"3042FFFF";
        ram_buffer(44393) := X"30420002";
        ram_buffer(44394) := X"14400004";
        ram_buffer(44395) := X"00000000";
        ram_buffer(44396) := X"8E020014";
        ram_buffer(44397) := X"10000002";
        ram_buffer(44398) := X"00000000";
        ram_buffer(44399) := X"00001021";
        ram_buffer(44400) := X"AE020008";
        ram_buffer(44401) := X"8E020010";
        ram_buffer(44402) := X"00000000";
        ram_buffer(44403) := X"14400010";
        ram_buffer(44404) := X"00000000";
        ram_buffer(44405) := X"8602000C";
        ram_buffer(44406) := X"00000000";
        ram_buffer(44407) := X"3042FFFF";
        ram_buffer(44408) := X"30420080";
        ram_buffer(44409) := X"1040000A";
        ram_buffer(44410) := X"00000000";
        ram_buffer(44411) := X"8602000C";
        ram_buffer(44412) := X"00000000";
        ram_buffer(44413) := X"34420040";
        ram_buffer(44414) := X"00021400";
        ram_buffer(44415) := X"00021403";
        ram_buffer(44416) := X"A602000C";
        ram_buffer(44417) := X"2402FFFF";
        ram_buffer(44418) := X"10000002";
        ram_buffer(44419) := X"00000000";
        ram_buffer(44420) := X"00001021";
        ram_buffer(44421) := X"03C0E821";
        ram_buffer(44422) := X"8FBF0024";
        ram_buffer(44423) := X"8FBE0020";
        ram_buffer(44424) := X"8FB0001C";
        ram_buffer(44425) := X"27BD0028";
        ram_buffer(44426) := X"03E00008";
        ram_buffer(44427) := X"00000000";
        ram_buffer(44428) := X"27BDFFC8";
        ram_buffer(44429) := X"AFBF0034";
        ram_buffer(44430) := X"AFBE0030";
        ram_buffer(44431) := X"AFB2002C";
        ram_buffer(44432) := X"AFB10028";
        ram_buffer(44433) := X"AFB00024";
        ram_buffer(44434) := X"03A0F021";
        ram_buffer(44435) := X"AFC40038";
        ram_buffer(44436) := X"AFC5003C";
        ram_buffer(44437) := X"8F82809C";
        ram_buffer(44438) := X"00000000";
        ram_buffer(44439) := X"8C500148";
        ram_buffer(44440) := X"8F82809C";
        ram_buffer(44441) := X"00000000";
        ram_buffer(44442) := X"24420148";
        ram_buffer(44443) := X"AFC20010";
        ram_buffer(44444) := X"10000088";
        ram_buffer(44445) := X"00000000";
        ram_buffer(44446) := X"26120088";
        ram_buffer(44447) := X"8E020004";
        ram_buffer(44448) := X"00000000";
        ram_buffer(44449) := X"2451FFFF";
        ram_buffer(44450) := X"10000065";
        ram_buffer(44451) := X"00000000";
        ram_buffer(44452) := X"24020001";
        ram_buffer(44453) := X"02221004";
        ram_buffer(44454) := X"AFC20014";
        ram_buffer(44455) := X"8FC2003C";
        ram_buffer(44456) := X"00000000";
        ram_buffer(44457) := X"1040000B";
        ram_buffer(44458) := X"00000000";
        ram_buffer(44459) := X"12400057";
        ram_buffer(44460) := X"00000000";
        ram_buffer(44461) := X"26220020";
        ram_buffer(44462) := X"00021080";
        ram_buffer(44463) := X"02421021";
        ram_buffer(44464) := X"8C430000";
        ram_buffer(44465) := X"8FC2003C";
        ram_buffer(44466) := X"00000000";
        ram_buffer(44467) := X"1462004F";
        ram_buffer(44468) := X"00000000";
        ram_buffer(44469) := X"26220002";
        ram_buffer(44470) := X"00021080";
        ram_buffer(44471) := X"02021021";
        ram_buffer(44472) := X"8C420000";
        ram_buffer(44473) := X"00000000";
        ram_buffer(44474) := X"AFC20018";
        ram_buffer(44475) := X"8E020004";
        ram_buffer(44476) := X"00000000";
        ram_buffer(44477) := X"2442FFFF";
        ram_buffer(44478) := X"14510007";
        ram_buffer(44479) := X"00000000";
        ram_buffer(44480) := X"8E020004";
        ram_buffer(44481) := X"00000000";
        ram_buffer(44482) := X"2442FFFF";
        ram_buffer(44483) := X"AE020004";
        ram_buffer(44484) := X"10000005";
        ram_buffer(44485) := X"00000000";
        ram_buffer(44486) := X"26220002";
        ram_buffer(44487) := X"00021080";
        ram_buffer(44488) := X"02021021";
        ram_buffer(44489) := X"AC400000";
        ram_buffer(44490) := X"8FC20018";
        ram_buffer(44491) := X"00000000";
        ram_buffer(44492) := X"10400039";
        ram_buffer(44493) := X"00000000";
        ram_buffer(44494) := X"8E020004";
        ram_buffer(44495) := X"00000000";
        ram_buffer(44496) := X"AFC2001C";
        ram_buffer(44497) := X"12400007";
        ram_buffer(44498) := X"00000000";
        ram_buffer(44499) := X"8E430100";
        ram_buffer(44500) := X"8FC20014";
        ram_buffer(44501) := X"00000000";
        ram_buffer(44502) := X"00621024";
        ram_buffer(44503) := X"14400007";
        ram_buffer(44504) := X"00000000";
        ram_buffer(44505) := X"8FC20018";
        ram_buffer(44506) := X"00000000";
        ram_buffer(44507) := X"0040F809";
        ram_buffer(44508) := X"00000000";
        ram_buffer(44509) := X"10000018";
        ram_buffer(44510) := X"00000000";
        ram_buffer(44511) := X"8E430104";
        ram_buffer(44512) := X"8FC20014";
        ram_buffer(44513) := X"00000000";
        ram_buffer(44514) := X"00621024";
        ram_buffer(44515) := X"1440000B";
        ram_buffer(44516) := X"00000000";
        ram_buffer(44517) := X"00111080";
        ram_buffer(44518) := X"02421021";
        ram_buffer(44519) := X"8C430000";
        ram_buffer(44520) := X"8FC20018";
        ram_buffer(44521) := X"00602821";
        ram_buffer(44522) := X"8FC40038";
        ram_buffer(44523) := X"0040F809";
        ram_buffer(44524) := X"00000000";
        ram_buffer(44525) := X"10000008";
        ram_buffer(44526) := X"00000000";
        ram_buffer(44527) := X"00111080";
        ram_buffer(44528) := X"02421021";
        ram_buffer(44529) := X"8C430000";
        ram_buffer(44530) := X"8FC20018";
        ram_buffer(44531) := X"00602021";
        ram_buffer(44532) := X"0040F809";
        ram_buffer(44533) := X"00000000";
        ram_buffer(44534) := X"8E030004";
        ram_buffer(44535) := X"8FC2001C";
        ram_buffer(44536) := X"00000000";
        ram_buffer(44537) := X"1462FF9B";
        ram_buffer(44538) := X"00000000";
        ram_buffer(44539) := X"8FC20010";
        ram_buffer(44540) := X"00000000";
        ram_buffer(44541) := X"8C420000";
        ram_buffer(44542) := X"00000000";
        ram_buffer(44543) := X"1450FF95";
        ram_buffer(44544) := X"00000000";
        ram_buffer(44545) := X"10000005";
        ram_buffer(44546) := X"00000000";
        ram_buffer(44547) := X"00000000";
        ram_buffer(44548) := X"10000002";
        ram_buffer(44549) := X"00000000";
        ram_buffer(44550) := X"00000000";
        ram_buffer(44551) := X"2631FFFF";
        ram_buffer(44552) := X"0621FF9B";
        ram_buffer(44553) := X"00000000";
        ram_buffer(44554) := X"3C02100A";
        ram_buffer(44555) := X"2442E934";
        ram_buffer(44556) := X"1040001C";
        ram_buffer(44557) := X"00000000";
        ram_buffer(44558) := X"8E020004";
        ram_buffer(44559) := X"00000000";
        ram_buffer(44560) := X"14400011";
        ram_buffer(44561) := X"00000000";
        ram_buffer(44562) := X"8E020000";
        ram_buffer(44563) := X"00000000";
        ram_buffer(44564) := X"1040000D";
        ram_buffer(44565) := X"00000000";
        ram_buffer(44566) := X"8E030000";
        ram_buffer(44567) := X"8FC20010";
        ram_buffer(44568) := X"00000000";
        ram_buffer(44569) := X"AC430000";
        ram_buffer(44570) := X"02002021";
        ram_buffer(44571) := X"0C027A4D";
        ram_buffer(44572) := X"00000000";
        ram_buffer(44573) := X"8FC20010";
        ram_buffer(44574) := X"00000000";
        ram_buffer(44575) := X"8C500000";
        ram_buffer(44576) := X"10000004";
        ram_buffer(44577) := X"00000000";
        ram_buffer(44578) := X"AFD00010";
        ram_buffer(44579) := X"8E100000";
        ram_buffer(44580) := X"00000000";
        ram_buffer(44581) := X"1600FF78";
        ram_buffer(44582) := X"00000000";
        ram_buffer(44583) := X"10000002";
        ram_buffer(44584) := X"00000000";
        ram_buffer(44585) := X"00000000";
        ram_buffer(44586) := X"00000000";
        ram_buffer(44587) := X"03C0E821";
        ram_buffer(44588) := X"8FBF0034";
        ram_buffer(44589) := X"8FBE0030";
        ram_buffer(44590) := X"8FB2002C";
        ram_buffer(44591) := X"8FB10028";
        ram_buffer(44592) := X"8FB00024";
        ram_buffer(44593) := X"27BD0038";
        ram_buffer(44594) := X"03E00008";
        ram_buffer(44595) := X"00000000";
        ram_buffer(44596) := X"27BDFFE0";
        ram_buffer(44597) := X"AFBF001C";
        ram_buffer(44598) := X"AFBE0018";
        ram_buffer(44599) := X"03A0F021";
        ram_buffer(44600) := X"AFC40020";
        ram_buffer(44601) := X"AFC50024";
        ram_buffer(44602) := X"AF8081EC";
        ram_buffer(44603) := X"8FC40024";
        ram_buffer(44604) := X"0C02FB69";
        ram_buffer(44605) := X"00000000";
        ram_buffer(44606) := X"AFC20010";
        ram_buffer(44607) := X"8FC30010";
        ram_buffer(44608) := X"2402FFFF";
        ram_buffer(44609) := X"14620009";
        ram_buffer(44610) := X"00000000";
        ram_buffer(44611) := X"8F8281EC";
        ram_buffer(44612) := X"00000000";
        ram_buffer(44613) := X"10400005";
        ram_buffer(44614) := X"00000000";
        ram_buffer(44615) := X"8F8381EC";
        ram_buffer(44616) := X"8FC20020";
        ram_buffer(44617) := X"00000000";
        ram_buffer(44618) := X"AC430000";
        ram_buffer(44619) := X"8FC20010";
        ram_buffer(44620) := X"03C0E821";
        ram_buffer(44621) := X"8FBF001C";
        ram_buffer(44622) := X"8FBE0018";
        ram_buffer(44623) := X"27BD0020";
        ram_buffer(44624) := X"03E00008";
        ram_buffer(44625) := X"00000000";
        ram_buffer(44626) := X"27BDFFB0";
        ram_buffer(44627) := X"AFBF004C";
        ram_buffer(44628) := X"AFBE0048";
        ram_buffer(44629) := X"03A0F021";
        ram_buffer(44630) := X"AFC40050";
        ram_buffer(44631) := X"AFC50054";
        ram_buffer(44632) := X"8FC20054";
        ram_buffer(44633) := X"00000000";
        ram_buffer(44634) := X"8C420010";
        ram_buffer(44635) := X"00000000";
        ram_buffer(44636) := X"AFC20010";
        ram_buffer(44637) := X"8FC20050";
        ram_buffer(44638) := X"00000000";
        ram_buffer(44639) := X"8C430010";
        ram_buffer(44640) := X"8FC20010";
        ram_buffer(44641) := X"00000000";
        ram_buffer(44642) := X"0062102A";
        ram_buffer(44643) := X"10400004";
        ram_buffer(44644) := X"00000000";
        ram_buffer(44645) := X"00001021";
        ram_buffer(44646) := X"10000136";
        ram_buffer(44647) := X"00000000";
        ram_buffer(44648) := X"8FC20054";
        ram_buffer(44649) := X"00000000";
        ram_buffer(44650) := X"24420014";
        ram_buffer(44651) := X"AFC20028";
        ram_buffer(44652) := X"8FC20010";
        ram_buffer(44653) := X"00000000";
        ram_buffer(44654) := X"2442FFFF";
        ram_buffer(44655) := X"AFC20010";
        ram_buffer(44656) := X"8FC20010";
        ram_buffer(44657) := X"00000000";
        ram_buffer(44658) := X"00021080";
        ram_buffer(44659) := X"8FC30028";
        ram_buffer(44660) := X"00000000";
        ram_buffer(44661) := X"00621021";
        ram_buffer(44662) := X"AFC2002C";
        ram_buffer(44663) := X"8FC20050";
        ram_buffer(44664) := X"00000000";
        ram_buffer(44665) := X"24420014";
        ram_buffer(44666) := X"AFC20020";
        ram_buffer(44667) := X"8FC20010";
        ram_buffer(44668) := X"00000000";
        ram_buffer(44669) := X"00021080";
        ram_buffer(44670) := X"8FC30020";
        ram_buffer(44671) := X"00000000";
        ram_buffer(44672) := X"00621021";
        ram_buffer(44673) := X"AFC20024";
        ram_buffer(44674) := X"8FC20024";
        ram_buffer(44675) := X"00000000";
        ram_buffer(44676) := X"8C430000";
        ram_buffer(44677) := X"8FC2002C";
        ram_buffer(44678) := X"00000000";
        ram_buffer(44679) := X"8C420000";
        ram_buffer(44680) := X"00000000";
        ram_buffer(44681) := X"24420001";
        ram_buffer(44682) := X"14400002";
        ram_buffer(44683) := X"0062001B";
        ram_buffer(44684) := X"0007000D";
        ram_buffer(44685) := X"00001010";
        ram_buffer(44686) := X"00001012";
        ram_buffer(44687) := X"AFC2001C";
        ram_buffer(44688) := X"8FC2001C";
        ram_buffer(44689) := X"00000000";
        ram_buffer(44690) := X"1040007C";
        ram_buffer(44691) := X"00000000";
        ram_buffer(44692) := X"AFC00014";
        ram_buffer(44693) := X"AFC00018";
        ram_buffer(44694) := X"8FC20028";
        ram_buffer(44695) := X"00000000";
        ram_buffer(44696) := X"24430004";
        ram_buffer(44697) := X"AFC30028";
        ram_buffer(44698) := X"8C420000";
        ram_buffer(44699) := X"00000000";
        ram_buffer(44700) := X"AFC20030";
        ram_buffer(44701) := X"8FC20030";
        ram_buffer(44702) := X"00000000";
        ram_buffer(44703) := X"3043FFFF";
        ram_buffer(44704) := X"8FC2001C";
        ram_buffer(44705) := X"00000000";
        ram_buffer(44706) := X"00620018";
        ram_buffer(44707) := X"8FC20018";
        ram_buffer(44708) := X"00001812";
        ram_buffer(44709) := X"00621021";
        ram_buffer(44710) := X"AFC20034";
        ram_buffer(44711) := X"8FC20030";
        ram_buffer(44712) := X"00000000";
        ram_buffer(44713) := X"00021C02";
        ram_buffer(44714) := X"8FC2001C";
        ram_buffer(44715) := X"00000000";
        ram_buffer(44716) := X"00620018";
        ram_buffer(44717) := X"8FC20034";
        ram_buffer(44718) := X"00000000";
        ram_buffer(44719) := X"00021402";
        ram_buffer(44720) := X"00001812";
        ram_buffer(44721) := X"00621021";
        ram_buffer(44722) := X"AFC20038";
        ram_buffer(44723) := X"8FC20038";
        ram_buffer(44724) := X"00000000";
        ram_buffer(44725) := X"00021402";
        ram_buffer(44726) := X"AFC20018";
        ram_buffer(44727) := X"8FC20020";
        ram_buffer(44728) := X"00000000";
        ram_buffer(44729) := X"8C420000";
        ram_buffer(44730) := X"00000000";
        ram_buffer(44731) := X"3043FFFF";
        ram_buffer(44732) := X"8FC20034";
        ram_buffer(44733) := X"00000000";
        ram_buffer(44734) := X"3042FFFF";
        ram_buffer(44735) := X"00621823";
        ram_buffer(44736) := X"8FC20014";
        ram_buffer(44737) := X"00000000";
        ram_buffer(44738) := X"00621021";
        ram_buffer(44739) := X"AFC2003C";
        ram_buffer(44740) := X"8FC2003C";
        ram_buffer(44741) := X"00000000";
        ram_buffer(44742) := X"00021403";
        ram_buffer(44743) := X"AFC20014";
        ram_buffer(44744) := X"8FC20020";
        ram_buffer(44745) := X"00000000";
        ram_buffer(44746) := X"8C420000";
        ram_buffer(44747) := X"00000000";
        ram_buffer(44748) := X"00021C02";
        ram_buffer(44749) := X"8FC20038";
        ram_buffer(44750) := X"00000000";
        ram_buffer(44751) := X"3042FFFF";
        ram_buffer(44752) := X"00621823";
        ram_buffer(44753) := X"8FC20014";
        ram_buffer(44754) := X"00000000";
        ram_buffer(44755) := X"00621021";
        ram_buffer(44756) := X"AFC20040";
        ram_buffer(44757) := X"8FC20040";
        ram_buffer(44758) := X"00000000";
        ram_buffer(44759) := X"00021403";
        ram_buffer(44760) := X"AFC20014";
        ram_buffer(44761) := X"8FC20020";
        ram_buffer(44762) := X"00000000";
        ram_buffer(44763) := X"24430004";
        ram_buffer(44764) := X"AFC30020";
        ram_buffer(44765) := X"8FC30040";
        ram_buffer(44766) := X"00000000";
        ram_buffer(44767) := X"00032400";
        ram_buffer(44768) := X"8FC3003C";
        ram_buffer(44769) := X"00000000";
        ram_buffer(44770) := X"3063FFFF";
        ram_buffer(44771) := X"00831825";
        ram_buffer(44772) := X"AC430000";
        ram_buffer(44773) := X"8FC30028";
        ram_buffer(44774) := X"8FC2002C";
        ram_buffer(44775) := X"00000000";
        ram_buffer(44776) := X"0043102B";
        ram_buffer(44777) := X"1040FFAC";
        ram_buffer(44778) := X"00000000";
        ram_buffer(44779) := X"8FC20024";
        ram_buffer(44780) := X"00000000";
        ram_buffer(44781) := X"8C420000";
        ram_buffer(44782) := X"00000000";
        ram_buffer(44783) := X"1440001F";
        ram_buffer(44784) := X"00000000";
        ram_buffer(44785) := X"8FC20050";
        ram_buffer(44786) := X"00000000";
        ram_buffer(44787) := X"24420014";
        ram_buffer(44788) := X"AFC20020";
        ram_buffer(44789) := X"10000005";
        ram_buffer(44790) := X"00000000";
        ram_buffer(44791) := X"8FC20010";
        ram_buffer(44792) := X"00000000";
        ram_buffer(44793) := X"2442FFFF";
        ram_buffer(44794) := X"AFC20010";
        ram_buffer(44795) := X"8FC20024";
        ram_buffer(44796) := X"00000000";
        ram_buffer(44797) := X"2442FFFC";
        ram_buffer(44798) := X"AFC20024";
        ram_buffer(44799) := X"8FC30024";
        ram_buffer(44800) := X"8FC20020";
        ram_buffer(44801) := X"00000000";
        ram_buffer(44802) := X"0043102B";
        ram_buffer(44803) := X"10400007";
        ram_buffer(44804) := X"00000000";
        ram_buffer(44805) := X"8FC20024";
        ram_buffer(44806) := X"00000000";
        ram_buffer(44807) := X"8C420000";
        ram_buffer(44808) := X"00000000";
        ram_buffer(44809) := X"1040FFED";
        ram_buffer(44810) := X"00000000";
        ram_buffer(44811) := X"8FC20050";
        ram_buffer(44812) := X"8FC30010";
        ram_buffer(44813) := X"00000000";
        ram_buffer(44814) := X"AC430010";
        ram_buffer(44815) := X"8FC50054";
        ram_buffer(44816) := X"8FC40050";
        ram_buffer(44817) := X"0C02C26D";
        ram_buffer(44818) := X"00000000";
        ram_buffer(44819) := X"04400088";
        ram_buffer(44820) := X"00000000";
        ram_buffer(44821) := X"8FC2001C";
        ram_buffer(44822) := X"00000000";
        ram_buffer(44823) := X"24420001";
        ram_buffer(44824) := X"AFC2001C";
        ram_buffer(44825) := X"AFC00014";
        ram_buffer(44826) := X"AFC00018";
        ram_buffer(44827) := X"8FC20050";
        ram_buffer(44828) := X"00000000";
        ram_buffer(44829) := X"24420014";
        ram_buffer(44830) := X"AFC20020";
        ram_buffer(44831) := X"8FC20054";
        ram_buffer(44832) := X"00000000";
        ram_buffer(44833) := X"24420014";
        ram_buffer(44834) := X"AFC20028";
        ram_buffer(44835) := X"8FC20028";
        ram_buffer(44836) := X"00000000";
        ram_buffer(44837) := X"24430004";
        ram_buffer(44838) := X"AFC30028";
        ram_buffer(44839) := X"8C420000";
        ram_buffer(44840) := X"00000000";
        ram_buffer(44841) := X"AFC20030";
        ram_buffer(44842) := X"8FC20030";
        ram_buffer(44843) := X"00000000";
        ram_buffer(44844) := X"3043FFFF";
        ram_buffer(44845) := X"8FC20018";
        ram_buffer(44846) := X"00000000";
        ram_buffer(44847) := X"00621021";
        ram_buffer(44848) := X"AFC20034";
        ram_buffer(44849) := X"8FC20030";
        ram_buffer(44850) := X"00000000";
        ram_buffer(44851) := X"00021C02";
        ram_buffer(44852) := X"8FC20034";
        ram_buffer(44853) := X"00000000";
        ram_buffer(44854) := X"00021402";
        ram_buffer(44855) := X"00621021";
        ram_buffer(44856) := X"AFC20038";
        ram_buffer(44857) := X"8FC20038";
        ram_buffer(44858) := X"00000000";
        ram_buffer(44859) := X"00021402";
        ram_buffer(44860) := X"AFC20018";
        ram_buffer(44861) := X"8FC20020";
        ram_buffer(44862) := X"00000000";
        ram_buffer(44863) := X"8C420000";
        ram_buffer(44864) := X"00000000";
        ram_buffer(44865) := X"3043FFFF";
        ram_buffer(44866) := X"8FC20034";
        ram_buffer(44867) := X"00000000";
        ram_buffer(44868) := X"3042FFFF";
        ram_buffer(44869) := X"00621823";
        ram_buffer(44870) := X"8FC20014";
        ram_buffer(44871) := X"00000000";
        ram_buffer(44872) := X"00621021";
        ram_buffer(44873) := X"AFC2003C";
        ram_buffer(44874) := X"8FC2003C";
        ram_buffer(44875) := X"00000000";
        ram_buffer(44876) := X"00021403";
        ram_buffer(44877) := X"AFC20014";
        ram_buffer(44878) := X"8FC20020";
        ram_buffer(44879) := X"00000000";
        ram_buffer(44880) := X"8C420000";
        ram_buffer(44881) := X"00000000";
        ram_buffer(44882) := X"00021C02";
        ram_buffer(44883) := X"8FC20038";
        ram_buffer(44884) := X"00000000";
        ram_buffer(44885) := X"3042FFFF";
        ram_buffer(44886) := X"00621823";
        ram_buffer(44887) := X"8FC20014";
        ram_buffer(44888) := X"00000000";
        ram_buffer(44889) := X"00621021";
        ram_buffer(44890) := X"AFC20040";
        ram_buffer(44891) := X"8FC20040";
        ram_buffer(44892) := X"00000000";
        ram_buffer(44893) := X"00021403";
        ram_buffer(44894) := X"AFC20014";
        ram_buffer(44895) := X"8FC20020";
        ram_buffer(44896) := X"00000000";
        ram_buffer(44897) := X"24430004";
        ram_buffer(44898) := X"AFC30020";
        ram_buffer(44899) := X"8FC30040";
        ram_buffer(44900) := X"00000000";
        ram_buffer(44901) := X"00032400";
        ram_buffer(44902) := X"8FC3003C";
        ram_buffer(44903) := X"00000000";
        ram_buffer(44904) := X"3063FFFF";
        ram_buffer(44905) := X"00831825";
        ram_buffer(44906) := X"AC430000";
        ram_buffer(44907) := X"8FC30028";
        ram_buffer(44908) := X"8FC2002C";
        ram_buffer(44909) := X"00000000";
        ram_buffer(44910) := X"0043102B";
        ram_buffer(44911) := X"1040FFB3";
        ram_buffer(44912) := X"00000000";
        ram_buffer(44913) := X"8FC20050";
        ram_buffer(44914) := X"00000000";
        ram_buffer(44915) := X"24420014";
        ram_buffer(44916) := X"AFC20020";
        ram_buffer(44917) := X"8FC20010";
        ram_buffer(44918) := X"00000000";
        ram_buffer(44919) := X"00021080";
        ram_buffer(44920) := X"8FC30020";
        ram_buffer(44921) := X"00000000";
        ram_buffer(44922) := X"00621021";
        ram_buffer(44923) := X"AFC20024";
        ram_buffer(44924) := X"8FC20024";
        ram_buffer(44925) := X"00000000";
        ram_buffer(44926) := X"8C420000";
        ram_buffer(44927) := X"00000000";
        ram_buffer(44928) := X"1440001B";
        ram_buffer(44929) := X"00000000";
        ram_buffer(44930) := X"10000005";
        ram_buffer(44931) := X"00000000";
        ram_buffer(44932) := X"8FC20010";
        ram_buffer(44933) := X"00000000";
        ram_buffer(44934) := X"2442FFFF";
        ram_buffer(44935) := X"AFC20010";
        ram_buffer(44936) := X"8FC20024";
        ram_buffer(44937) := X"00000000";
        ram_buffer(44938) := X"2442FFFC";
        ram_buffer(44939) := X"AFC20024";
        ram_buffer(44940) := X"8FC30024";
        ram_buffer(44941) := X"8FC20020";
        ram_buffer(44942) := X"00000000";
        ram_buffer(44943) := X"0043102B";
        ram_buffer(44944) := X"10400007";
        ram_buffer(44945) := X"00000000";
        ram_buffer(44946) := X"8FC20024";
        ram_buffer(44947) := X"00000000";
        ram_buffer(44948) := X"8C420000";
        ram_buffer(44949) := X"00000000";
        ram_buffer(44950) := X"1040FFED";
        ram_buffer(44951) := X"00000000";
        ram_buffer(44952) := X"8FC20050";
        ram_buffer(44953) := X"8FC30010";
        ram_buffer(44954) := X"00000000";
        ram_buffer(44955) := X"AC430010";
        ram_buffer(44956) := X"8FC2001C";
        ram_buffer(44957) := X"03C0E821";
        ram_buffer(44958) := X"8FBF004C";
        ram_buffer(44959) := X"8FBE0048";
        ram_buffer(44960) := X"27BD0050";
        ram_buffer(44961) := X"03E00008";
        ram_buffer(44962) := X"00000000";
        ram_buffer(44963) := X"27BDFF28";
        ram_buffer(44964) := X"AFBF00D4";
        ram_buffer(44965) := X"AFBE00D0";
        ram_buffer(44966) := X"AFB300CC";
        ram_buffer(44967) := X"AFB200C8";
        ram_buffer(44968) := X"AFB100C4";
        ram_buffer(44969) := X"AFB000C0";
        ram_buffer(44970) := X"03A0F021";
        ram_buffer(44971) := X"AFC400D8";
        ram_buffer(44972) := X"AFC700E4";
        ram_buffer(44973) := X"AFC600E0";
        ram_buffer(44974) := X"AFC00064";
        ram_buffer(44975) := X"8FC300E4";
        ram_buffer(44976) := X"8FC200E0";
        ram_buffer(44977) := X"AFC300AC";
        ram_buffer(44978) := X"AFC200A8";
        ram_buffer(44979) := X"8FC200D8";
        ram_buffer(44980) := X"00000000";
        ram_buffer(44981) := X"8C420040";
        ram_buffer(44982) := X"00000000";
        ram_buffer(44983) := X"1040001D";
        ram_buffer(44984) := X"00000000";
        ram_buffer(44985) := X"8FC200D8";
        ram_buffer(44986) := X"00000000";
        ram_buffer(44987) := X"8C420040";
        ram_buffer(44988) := X"8FC300D8";
        ram_buffer(44989) := X"00000000";
        ram_buffer(44990) := X"8C630044";
        ram_buffer(44991) := X"00000000";
        ram_buffer(44992) := X"AC430004";
        ram_buffer(44993) := X"8FC200D8";
        ram_buffer(44994) := X"00000000";
        ram_buffer(44995) := X"8C420040";
        ram_buffer(44996) := X"8FC300D8";
        ram_buffer(44997) := X"00000000";
        ram_buffer(44998) := X"8C630044";
        ram_buffer(44999) := X"24040001";
        ram_buffer(45000) := X"00641804";
        ram_buffer(45001) := X"AC430008";
        ram_buffer(45002) := X"8FC200D8";
        ram_buffer(45003) := X"00000000";
        ram_buffer(45004) := X"8C420040";
        ram_buffer(45005) := X"00000000";
        ram_buffer(45006) := X"00402821";
        ram_buffer(45007) := X"8FC400D8";
        ram_buffer(45008) := X"0C02BE10";
        ram_buffer(45009) := X"00000000";
        ram_buffer(45010) := X"8FC200D8";
        ram_buffer(45011) := X"00000000";
        ram_buffer(45012) := X"AC400040";
        ram_buffer(45013) := X"8FC200A8";
        ram_buffer(45014) := X"00000000";
        ram_buffer(45015) := X"0441000B";
        ram_buffer(45016) := X"00000000";
        ram_buffer(45017) := X"8FC200F4";
        ram_buffer(45018) := X"24030001";
        ram_buffer(45019) := X"AC430000";
        ram_buffer(45020) := X"8FC300A8";
        ram_buffer(45021) := X"3C027FFF";
        ram_buffer(45022) := X"3442FFFF";
        ram_buffer(45023) := X"00621024";
        ram_buffer(45024) := X"AFC200A8";
        ram_buffer(45025) := X"10000004";
        ram_buffer(45026) := X"00000000";
        ram_buffer(45027) := X"8FC200F4";
        ram_buffer(45028) := X"00000000";
        ram_buffer(45029) := X"AC400000";
        ram_buffer(45030) := X"8FC300A8";
        ram_buffer(45031) := X"3C027FF0";
        ram_buffer(45032) := X"00621824";
        ram_buffer(45033) := X"3C027FF0";
        ram_buffer(45034) := X"1462002E";
        ram_buffer(45035) := X"00000000";
        ram_buffer(45036) := X"8FC200F0";
        ram_buffer(45037) := X"2403270F";
        ram_buffer(45038) := X"AC430000";
        ram_buffer(45039) := X"8FC200AC";
        ram_buffer(45040) := X"00000000";
        ram_buffer(45041) := X"1440000B";
        ram_buffer(45042) := X"00000000";
        ram_buffer(45043) := X"8FC300A8";
        ram_buffer(45044) := X"3C02000F";
        ram_buffer(45045) := X"3442FFFF";
        ram_buffer(45046) := X"00621024";
        ram_buffer(45047) := X"14400005";
        ram_buffer(45048) := X"00000000";
        ram_buffer(45049) := X"3C02100D";
        ram_buffer(45050) := X"2442A8F0";
        ram_buffer(45051) := X"10000003";
        ram_buffer(45052) := X"00000000";
        ram_buffer(45053) := X"3C02100D";
        ram_buffer(45054) := X"2442A8FC";
        ram_buffer(45055) := X"AFC20078";
        ram_buffer(45056) := X"8FC200F8";
        ram_buffer(45057) := X"00000000";
        ram_buffer(45058) := X"10400013";
        ram_buffer(45059) := X"00000000";
        ram_buffer(45060) := X"8FC20078";
        ram_buffer(45061) := X"00000000";
        ram_buffer(45062) := X"24420003";
        ram_buffer(45063) := X"80420000";
        ram_buffer(45064) := X"00000000";
        ram_buffer(45065) := X"10400006";
        ram_buffer(45066) := X"00000000";
        ram_buffer(45067) := X"8FC20078";
        ram_buffer(45068) := X"00000000";
        ram_buffer(45069) := X"24420008";
        ram_buffer(45070) := X"10000004";
        ram_buffer(45071) := X"00000000";
        ram_buffer(45072) := X"8FC20078";
        ram_buffer(45073) := X"00000000";
        ram_buffer(45074) := X"24420003";
        ram_buffer(45075) := X"8FC300F8";
        ram_buffer(45076) := X"00000000";
        ram_buffer(45077) := X"AC620000";
        ram_buffer(45078) := X"8FC20078";
        ram_buffer(45079) := X"10000810";
        ram_buffer(45080) := X"00000000";
        ram_buffer(45081) := X"8FC300AC";
        ram_buffer(45082) := X"8FC200A8";
        ram_buffer(45083) := X"00003821";
        ram_buffer(45084) := X"00003021";
        ram_buffer(45085) := X"00602821";
        ram_buffer(45086) := X"00402021";
        ram_buffer(45087) := X"0C03167F";
        ram_buffer(45088) := X"00000000";
        ram_buffer(45089) := X"14400014";
        ram_buffer(45090) := X"00000000";
        ram_buffer(45091) := X"8FC200F0";
        ram_buffer(45092) := X"24030001";
        ram_buffer(45093) := X"AC430000";
        ram_buffer(45094) := X"3C02100D";
        ram_buffer(45095) := X"2442A900";
        ram_buffer(45096) := X"AFC20078";
        ram_buffer(45097) := X"8FC200F8";
        ram_buffer(45098) := X"00000000";
        ram_buffer(45099) := X"10400007";
        ram_buffer(45100) := X"00000000";
        ram_buffer(45101) := X"8FC20078";
        ram_buffer(45102) := X"00000000";
        ram_buffer(45103) := X"24430001";
        ram_buffer(45104) := X"8FC200F8";
        ram_buffer(45105) := X"00000000";
        ram_buffer(45106) := X"AC430000";
        ram_buffer(45107) := X"8FC20078";
        ram_buffer(45108) := X"100007F3";
        ram_buffer(45109) := X"00000000";
        ram_buffer(45110) := X"8FC300AC";
        ram_buffer(45111) := X"8FC200A8";
        ram_buffer(45112) := X"27C4009C";
        ram_buffer(45113) := X"AFA40014";
        ram_buffer(45114) := X"27C400A0";
        ram_buffer(45115) := X"AFA40010";
        ram_buffer(45116) := X"00603821";
        ram_buffer(45117) := X"00403021";
        ram_buffer(45118) := X"8FC400D8";
        ram_buffer(45119) := X"0C02C49D";
        ram_buffer(45120) := X"00000000";
        ram_buffer(45121) := X"AFC20060";
        ram_buffer(45122) := X"8FC200A8";
        ram_buffer(45123) := X"00000000";
        ram_buffer(45124) := X"00021502";
        ram_buffer(45125) := X"304207FF";
        ram_buffer(45126) := X"AFC20024";
        ram_buffer(45127) := X"8FC20024";
        ram_buffer(45128) := X"00000000";
        ram_buffer(45129) := X"10400015";
        ram_buffer(45130) := X"00000000";
        ram_buffer(45131) := X"8FC300AC";
        ram_buffer(45132) := X"8FC200A8";
        ram_buffer(45133) := X"AFC300B4";
        ram_buffer(45134) := X"AFC200B0";
        ram_buffer(45135) := X"8FC300B0";
        ram_buffer(45136) := X"3C02000F";
        ram_buffer(45137) := X"3442FFFF";
        ram_buffer(45138) := X"00621024";
        ram_buffer(45139) := X"AFC200B0";
        ram_buffer(45140) := X"8FC300B0";
        ram_buffer(45141) := X"3C023FF0";
        ram_buffer(45142) := X"00621025";
        ram_buffer(45143) := X"AFC200B0";
        ram_buffer(45144) := X"8FC20024";
        ram_buffer(45145) := X"00000000";
        ram_buffer(45146) := X"2442FC01";
        ram_buffer(45147) := X"AFC20024";
        ram_buffer(45148) := X"AFC0005C";
        ram_buffer(45149) := X"10000030";
        ram_buffer(45150) := X"00000000";
        ram_buffer(45151) := X"8FC3009C";
        ram_buffer(45152) := X"8FC200A0";
        ram_buffer(45153) := X"00000000";
        ram_buffer(45154) := X"00621021";
        ram_buffer(45155) := X"24420432";
        ram_buffer(45156) := X"AFC20024";
        ram_buffer(45157) := X"8FC20024";
        ram_buffer(45158) := X"00000000";
        ram_buffer(45159) := X"28420021";
        ram_buffer(45160) := X"1440000F";
        ram_buffer(45161) := X"00000000";
        ram_buffer(45162) := X"8FC300A8";
        ram_buffer(45163) := X"24040040";
        ram_buffer(45164) := X"8FC20024";
        ram_buffer(45165) := X"00000000";
        ram_buffer(45166) := X"00821023";
        ram_buffer(45167) := X"00431804";
        ram_buffer(45168) := X"8FC400AC";
        ram_buffer(45169) := X"8FC20024";
        ram_buffer(45170) := X"00000000";
        ram_buffer(45171) := X"2442FFE0";
        ram_buffer(45172) := X"00441006";
        ram_buffer(45173) := X"00621025";
        ram_buffer(45174) := X"10000007";
        ram_buffer(45175) := X"00000000";
        ram_buffer(45176) := X"8FC300AC";
        ram_buffer(45177) := X"24040020";
        ram_buffer(45178) := X"8FC20024";
        ram_buffer(45179) := X"00000000";
        ram_buffer(45180) := X"00821023";
        ram_buffer(45181) := X"00431004";
        ram_buffer(45182) := X"AFC2007C";
        ram_buffer(45183) := X"8FC4007C";
        ram_buffer(45184) := X"0C031BBD";
        ram_buffer(45185) := X"00000000";
        ram_buffer(45186) := X"AFC300B4";
        ram_buffer(45187) := X"AFC200B0";
        ram_buffer(45188) := X"8FC300B0";
        ram_buffer(45189) := X"3C02FE10";
        ram_buffer(45190) := X"00621021";
        ram_buffer(45191) := X"AFC200B0";
        ram_buffer(45192) := X"8FC20024";
        ram_buffer(45193) := X"00000000";
        ram_buffer(45194) := X"2442FBCD";
        ram_buffer(45195) := X"AFC20024";
        ram_buffer(45196) := X"24020001";
        ram_buffer(45197) := X"AFC2005C";
        ram_buffer(45198) := X"8FC300B4";
        ram_buffer(45199) := X"8FC200B0";
        ram_buffer(45200) := X"8F8780DC";
        ram_buffer(45201) := X"8F8680D8";
        ram_buffer(45202) := X"00602821";
        ram_buffer(45203) := X"00402021";
        ram_buffer(45204) := X"0C0318D3";
        ram_buffer(45205) := X"00000000";
        ram_buffer(45206) := X"8F8780E4";
        ram_buffer(45207) := X"8F8680E0";
        ram_buffer(45208) := X"00602821";
        ram_buffer(45209) := X"00402021";
        ram_buffer(45210) := X"0C03174A";
        ram_buffer(45211) := X"00000000";
        ram_buffer(45212) := X"8F8780EC";
        ram_buffer(45213) := X"8F8680E8";
        ram_buffer(45214) := X"00602821";
        ram_buffer(45215) := X"00402021";
        ram_buffer(45216) := X"0C0311FC";
        ram_buffer(45217) := X"00000000";
        ram_buffer(45218) := X"00609821";
        ram_buffer(45219) := X"00409021";
        ram_buffer(45220) := X"8FC40024";
        ram_buffer(45221) := X"0C031B7C";
        ram_buffer(45222) := X"00000000";
        ram_buffer(45223) := X"8F8780F4";
        ram_buffer(45224) := X"8F8680F0";
        ram_buffer(45225) := X"00602821";
        ram_buffer(45226) := X"00402021";
        ram_buffer(45227) := X"0C03174A";
        ram_buffer(45228) := X"00000000";
        ram_buffer(45229) := X"00603821";
        ram_buffer(45230) := X"00403021";
        ram_buffer(45231) := X"02602821";
        ram_buffer(45232) := X"02402021";
        ram_buffer(45233) := X"0C0311FC";
        ram_buffer(45234) := X"00000000";
        ram_buffer(45235) := X"AFC30074";
        ram_buffer(45236) := X"AFC20070";
        ram_buffer(45237) := X"8FC50074";
        ram_buffer(45238) := X"8FC40070";
        ram_buffer(45239) := X"0C031B37";
        ram_buffer(45240) := X"00000000";
        ram_buffer(45241) := X"AFC20038";
        ram_buffer(45242) := X"00003821";
        ram_buffer(45243) := X"00003021";
        ram_buffer(45244) := X"8FC50074";
        ram_buffer(45245) := X"8FC40070";
        ram_buffer(45246) := X"0C0316F7";
        ram_buffer(45247) := X"00000000";
        ram_buffer(45248) := X"04410010";
        ram_buffer(45249) := X"00000000";
        ram_buffer(45250) := X"8FC40038";
        ram_buffer(45251) := X"0C031B7C";
        ram_buffer(45252) := X"00000000";
        ram_buffer(45253) := X"8FC70074";
        ram_buffer(45254) := X"8FC60070";
        ram_buffer(45255) := X"00602821";
        ram_buffer(45256) := X"00402021";
        ram_buffer(45257) := X"0C03167F";
        ram_buffer(45258) := X"00000000";
        ram_buffer(45259) := X"10400005";
        ram_buffer(45260) := X"00000000";
        ram_buffer(45261) := X"8FC20038";
        ram_buffer(45262) := X"00000000";
        ram_buffer(45263) := X"2442FFFF";
        ram_buffer(45264) := X"AFC20038";
        ram_buffer(45265) := X"24020001";
        ram_buffer(45266) := X"AFC2003C";
        ram_buffer(45267) := X"8FC20038";
        ram_buffer(45268) := X"00000000";
        ram_buffer(45269) := X"0440001D";
        ram_buffer(45270) := X"00000000";
        ram_buffer(45271) := X"8FC20038";
        ram_buffer(45272) := X"00000000";
        ram_buffer(45273) := X"28420017";
        ram_buffer(45274) := X"10400018";
        ram_buffer(45275) := X"00000000";
        ram_buffer(45276) := X"8FC300AC";
        ram_buffer(45277) := X"8FC200A8";
        ram_buffer(45278) := X"3C04100D";
        ram_buffer(45279) := X"8FC50038";
        ram_buffer(45280) := X"00000000";
        ram_buffer(45281) := X"000528C0";
        ram_buffer(45282) := X"2484A938";
        ram_buffer(45283) := X"00A42021";
        ram_buffer(45284) := X"8C850004";
        ram_buffer(45285) := X"8C840000";
        ram_buffer(45286) := X"00A03821";
        ram_buffer(45287) := X"00803021";
        ram_buffer(45288) := X"00602821";
        ram_buffer(45289) := X"00402021";
        ram_buffer(45290) := X"0C0316F7";
        ram_buffer(45291) := X"00000000";
        ram_buffer(45292) := X"04410005";
        ram_buffer(45293) := X"00000000";
        ram_buffer(45294) := X"8FC20038";
        ram_buffer(45295) := X"00000000";
        ram_buffer(45296) := X"2442FFFF";
        ram_buffer(45297) := X"AFC20038";
        ram_buffer(45298) := X"AFC0003C";
        ram_buffer(45299) := X"8FC3009C";
        ram_buffer(45300) := X"8FC20024";
        ram_buffer(45301) := X"00000000";
        ram_buffer(45302) := X"00621023";
        ram_buffer(45303) := X"2442FFFF";
        ram_buffer(45304) := X"AFC20034";
        ram_buffer(45305) := X"8FC20034";
        ram_buffer(45306) := X"00000000";
        ram_buffer(45307) := X"04400007";
        ram_buffer(45308) := X"00000000";
        ram_buffer(45309) := X"AFC00018";
        ram_buffer(45310) := X"8FC20034";
        ram_buffer(45311) := X"00000000";
        ram_buffer(45312) := X"AFC2004C";
        ram_buffer(45313) := X"10000006";
        ram_buffer(45314) := X"00000000";
        ram_buffer(45315) := X"8FC20034";
        ram_buffer(45316) := X"00000000";
        ram_buffer(45317) := X"00021023";
        ram_buffer(45318) := X"AFC20018";
        ram_buffer(45319) := X"AFC0004C";
        ram_buffer(45320) := X"8FC20038";
        ram_buffer(45321) := X"00000000";
        ram_buffer(45322) := X"0440000C";
        ram_buffer(45323) := X"00000000";
        ram_buffer(45324) := X"AFC0001C";
        ram_buffer(45325) := X"8FC20038";
        ram_buffer(45326) := X"00000000";
        ram_buffer(45327) := X"AFC20050";
        ram_buffer(45328) := X"8FC3004C";
        ram_buffer(45329) := X"8FC20038";
        ram_buffer(45330) := X"00000000";
        ram_buffer(45331) := X"00621021";
        ram_buffer(45332) := X"AFC2004C";
        ram_buffer(45333) := X"1000000B";
        ram_buffer(45334) := X"00000000";
        ram_buffer(45335) := X"8FC30018";
        ram_buffer(45336) := X"8FC20038";
        ram_buffer(45337) := X"00000000";
        ram_buffer(45338) := X"00621023";
        ram_buffer(45339) := X"AFC20018";
        ram_buffer(45340) := X"8FC20038";
        ram_buffer(45341) := X"00000000";
        ram_buffer(45342) := X"00021023";
        ram_buffer(45343) := X"AFC2001C";
        ram_buffer(45344) := X"AFC00050";
        ram_buffer(45345) := X"8FC200E8";
        ram_buffer(45346) := X"00000000";
        ram_buffer(45347) := X"04400006";
        ram_buffer(45348) := X"00000000";
        ram_buffer(45349) := X"8FC200E8";
        ram_buffer(45350) := X"00000000";
        ram_buffer(45351) := X"2842000A";
        ram_buffer(45352) := X"14400002";
        ram_buffer(45353) := X"00000000";
        ram_buffer(45354) := X"AFC000E8";
        ram_buffer(45355) := X"24020001";
        ram_buffer(45356) := X"AFC20058";
        ram_buffer(45357) := X"8FC200E8";
        ram_buffer(45358) := X"00000000";
        ram_buffer(45359) := X"28420006";
        ram_buffer(45360) := X"14400006";
        ram_buffer(45361) := X"00000000";
        ram_buffer(45362) := X"8FC200E8";
        ram_buffer(45363) := X"00000000";
        ram_buffer(45364) := X"2442FFFC";
        ram_buffer(45365) := X"AFC200E8";
        ram_buffer(45366) := X"AFC00058";
        ram_buffer(45367) := X"24020001";
        ram_buffer(45368) := X"AFC20040";
        ram_buffer(45369) := X"2402FFFF";
        ram_buffer(45370) := X"AFC20030";
        ram_buffer(45371) := X"8FC20030";
        ram_buffer(45372) := X"00000000";
        ram_buffer(45373) := X"AFC2002C";
        ram_buffer(45374) := X"8FC200E8";
        ram_buffer(45375) := X"00000000";
        ram_buffer(45376) := X"2C420006";
        ram_buffer(45377) := X"10400036";
        ram_buffer(45378) := X"00000000";
        ram_buffer(45379) := X"8FC200E8";
        ram_buffer(45380) := X"00000000";
        ram_buffer(45381) := X"00021880";
        ram_buffer(45382) := X"3C02100D";
        ram_buffer(45383) := X"2442A904";
        ram_buffer(45384) := X"00621021";
        ram_buffer(45385) := X"8C420000";
        ram_buffer(45386) := X"00000000";
        ram_buffer(45387) := X"00400008";
        ram_buffer(45388) := X"00000000";
        ram_buffer(45389) := X"24020012";
        ram_buffer(45390) := X"AFC20024";
        ram_buffer(45391) := X"AFC000EC";
        ram_buffer(45392) := X"10000027";
        ram_buffer(45393) := X"00000000";
        ram_buffer(45394) := X"AFC00040";
        ram_buffer(45395) := X"8FC200EC";
        ram_buffer(45396) := X"00000000";
        ram_buffer(45397) := X"1C400003";
        ram_buffer(45398) := X"00000000";
        ram_buffer(45399) := X"24020001";
        ram_buffer(45400) := X"AFC200EC";
        ram_buffer(45401) := X"8FC200EC";
        ram_buffer(45402) := X"00000000";
        ram_buffer(45403) := X"AFC20024";
        ram_buffer(45404) := X"8FC20024";
        ram_buffer(45405) := X"00000000";
        ram_buffer(45406) := X"AFC20030";
        ram_buffer(45407) := X"8FC20030";
        ram_buffer(45408) := X"00000000";
        ram_buffer(45409) := X"AFC2002C";
        ram_buffer(45410) := X"10000015";
        ram_buffer(45411) := X"00000000";
        ram_buffer(45412) := X"AFC00040";
        ram_buffer(45413) := X"8FC300EC";
        ram_buffer(45414) := X"8FC20038";
        ram_buffer(45415) := X"00000000";
        ram_buffer(45416) := X"00621021";
        ram_buffer(45417) := X"24420001";
        ram_buffer(45418) := X"AFC20024";
        ram_buffer(45419) := X"8FC20024";
        ram_buffer(45420) := X"00000000";
        ram_buffer(45421) := X"AFC2002C";
        ram_buffer(45422) := X"8FC20024";
        ram_buffer(45423) := X"00000000";
        ram_buffer(45424) := X"2442FFFF";
        ram_buffer(45425) := X"AFC20030";
        ram_buffer(45426) := X"8FC20024";
        ram_buffer(45427) := X"00000000";
        ram_buffer(45428) := X"1C400003";
        ram_buffer(45429) := X"00000000";
        ram_buffer(45430) := X"24020001";
        ram_buffer(45431) := X"AFC20024";
        ram_buffer(45432) := X"24020004";
        ram_buffer(45433) := X"AFC20034";
        ram_buffer(45434) := X"8FC200D8";
        ram_buffer(45435) := X"00000000";
        ram_buffer(45436) := X"AC400044";
        ram_buffer(45437) := X"1000000D";
        ram_buffer(45438) := X"00000000";
        ram_buffer(45439) := X"8FC200D8";
        ram_buffer(45440) := X"00000000";
        ram_buffer(45441) := X"8C420044";
        ram_buffer(45442) := X"00000000";
        ram_buffer(45443) := X"24430001";
        ram_buffer(45444) := X"8FC200D8";
        ram_buffer(45445) := X"00000000";
        ram_buffer(45446) := X"AC430044";
        ram_buffer(45447) := X"8FC20034";
        ram_buffer(45448) := X"00000000";
        ram_buffer(45449) := X"00021040";
        ram_buffer(45450) := X"AFC20034";
        ram_buffer(45451) := X"8FC20034";
        ram_buffer(45452) := X"00000000";
        ram_buffer(45453) := X"24430014";
        ram_buffer(45454) := X"8FC20024";
        ram_buffer(45455) := X"00000000";
        ram_buffer(45456) := X"0043102B";
        ram_buffer(45457) := X"1040FFED";
        ram_buffer(45458) := X"00000000";
        ram_buffer(45459) := X"8FC200D8";
        ram_buffer(45460) := X"00000000";
        ram_buffer(45461) := X"8C420044";
        ram_buffer(45462) := X"00000000";
        ram_buffer(45463) := X"00402821";
        ram_buffer(45464) := X"8FC400D8";
        ram_buffer(45465) := X"0C02BDA8";
        ram_buffer(45466) := X"00000000";
        ram_buffer(45467) := X"00401821";
        ram_buffer(45468) := X"8FC200D8";
        ram_buffer(45469) := X"00000000";
        ram_buffer(45470) := X"AC430040";
        ram_buffer(45471) := X"8FC200D8";
        ram_buffer(45472) := X"00000000";
        ram_buffer(45473) := X"8C420040";
        ram_buffer(45474) := X"00000000";
        ram_buffer(45475) := X"AFC20080";
        ram_buffer(45476) := X"8FC20080";
        ram_buffer(45477) := X"00000000";
        ram_buffer(45478) := X"AFC20078";
        ram_buffer(45479) := X"8FC2002C";
        ram_buffer(45480) := X"00000000";
        ram_buffer(45481) := X"0440023C";
        ram_buffer(45482) := X"00000000";
        ram_buffer(45483) := X"8FC2002C";
        ram_buffer(45484) := X"00000000";
        ram_buffer(45485) := X"2842000F";
        ram_buffer(45486) := X"10400237";
        ram_buffer(45487) := X"00000000";
        ram_buffer(45488) := X"8FC20058";
        ram_buffer(45489) := X"00000000";
        ram_buffer(45490) := X"10400233";
        ram_buffer(45491) := X"00000000";
        ram_buffer(45492) := X"AFC00024";
        ram_buffer(45493) := X"8FC300AC";
        ram_buffer(45494) := X"8FC200A8";
        ram_buffer(45495) := X"AFC300B4";
        ram_buffer(45496) := X"AFC200B0";
        ram_buffer(45497) := X"8FC20038";
        ram_buffer(45498) := X"00000000";
        ram_buffer(45499) := X"AFC20084";
        ram_buffer(45500) := X"8FC2002C";
        ram_buffer(45501) := X"00000000";
        ram_buffer(45502) := X"AFC20088";
        ram_buffer(45503) := X"24020002";
        ram_buffer(45504) := X"AFC20028";
        ram_buffer(45505) := X"8FC20038";
        ram_buffer(45506) := X"00000000";
        ram_buffer(45507) := X"1840005E";
        ram_buffer(45508) := X"00000000";
        ram_buffer(45509) := X"8FC20038";
        ram_buffer(45510) := X"00000000";
        ram_buffer(45511) := X"3043000F";
        ram_buffer(45512) := X"3C02100D";
        ram_buffer(45513) := X"000318C0";
        ram_buffer(45514) := X"2442A938";
        ram_buffer(45515) := X"00621021";
        ram_buffer(45516) := X"8C430004";
        ram_buffer(45517) := X"8C420000";
        ram_buffer(45518) := X"AFC30074";
        ram_buffer(45519) := X"AFC20070";
        ram_buffer(45520) := X"8FC20038";
        ram_buffer(45521) := X"00000000";
        ram_buffer(45522) := X"00021103";
        ram_buffer(45523) := X"AFC20034";
        ram_buffer(45524) := X"8FC20034";
        ram_buffer(45525) := X"00000000";
        ram_buffer(45526) := X"30420010";
        ram_buffer(45527) := X"1040003A";
        ram_buffer(45528) := X"00000000";
        ram_buffer(45529) := X"8FC20034";
        ram_buffer(45530) := X"00000000";
        ram_buffer(45531) := X"3042000F";
        ram_buffer(45532) := X"AFC20034";
        ram_buffer(45533) := X"8FC300AC";
        ram_buffer(45534) := X"8FC200A8";
        ram_buffer(45535) := X"3C04100D";
        ram_buffer(45536) := X"2484AA00";
        ram_buffer(45537) := X"8C850024";
        ram_buffer(45538) := X"8C840020";
        ram_buffer(45539) := X"00A03821";
        ram_buffer(45540) := X"00803021";
        ram_buffer(45541) := X"00602821";
        ram_buffer(45542) := X"00402021";
        ram_buffer(45543) := X"0C03144F";
        ram_buffer(45544) := X"00000000";
        ram_buffer(45545) := X"AFC300AC";
        ram_buffer(45546) := X"AFC200A8";
        ram_buffer(45547) := X"8FC20028";
        ram_buffer(45548) := X"00000000";
        ram_buffer(45549) := X"24420001";
        ram_buffer(45550) := X"AFC20028";
        ram_buffer(45551) := X"10000022";
        ram_buffer(45552) := X"00000000";
        ram_buffer(45553) := X"8FC20034";
        ram_buffer(45554) := X"00000000";
        ram_buffer(45555) := X"30420001";
        ram_buffer(45556) := X"10400015";
        ram_buffer(45557) := X"00000000";
        ram_buffer(45558) := X"8FC20028";
        ram_buffer(45559) := X"00000000";
        ram_buffer(45560) := X"24420001";
        ram_buffer(45561) := X"AFC20028";
        ram_buffer(45562) := X"3C02100D";
        ram_buffer(45563) := X"8FC30024";
        ram_buffer(45564) := X"00000000";
        ram_buffer(45565) := X"000318C0";
        ram_buffer(45566) := X"2442AA00";
        ram_buffer(45567) := X"00621021";
        ram_buffer(45568) := X"8C430004";
        ram_buffer(45569) := X"8C420000";
        ram_buffer(45570) := X"00603821";
        ram_buffer(45571) := X"00403021";
        ram_buffer(45572) := X"8FC50074";
        ram_buffer(45573) := X"8FC40070";
        ram_buffer(45574) := X"0C03174A";
        ram_buffer(45575) := X"00000000";
        ram_buffer(45576) := X"AFC30074";
        ram_buffer(45577) := X"AFC20070";
        ram_buffer(45578) := X"8FC20034";
        ram_buffer(45579) := X"00000000";
        ram_buffer(45580) := X"00021043";
        ram_buffer(45581) := X"AFC20034";
        ram_buffer(45582) := X"8FC20024";
        ram_buffer(45583) := X"00000000";
        ram_buffer(45584) := X"24420001";
        ram_buffer(45585) := X"AFC20024";
        ram_buffer(45586) := X"8FC20034";
        ram_buffer(45587) := X"00000000";
        ram_buffer(45588) := X"1440FFDC";
        ram_buffer(45589) := X"00000000";
        ram_buffer(45590) := X"8FC300AC";
        ram_buffer(45591) := X"8FC200A8";
        ram_buffer(45592) := X"8FC70074";
        ram_buffer(45593) := X"8FC60070";
        ram_buffer(45594) := X"00602821";
        ram_buffer(45595) := X"00402021";
        ram_buffer(45596) := X"0C03144F";
        ram_buffer(45597) := X"00000000";
        ram_buffer(45598) := X"AFC300AC";
        ram_buffer(45599) := X"AFC200A8";
        ram_buffer(45600) := X"10000049";
        ram_buffer(45601) := X"00000000";
        ram_buffer(45602) := X"8FC20038";
        ram_buffer(45603) := X"00000000";
        ram_buffer(45604) := X"00021023";
        ram_buffer(45605) := X"AFC2008C";
        ram_buffer(45606) := X"8FC2008C";
        ram_buffer(45607) := X"00000000";
        ram_buffer(45608) := X"10400041";
        ram_buffer(45609) := X"00000000";
        ram_buffer(45610) := X"8FC300AC";
        ram_buffer(45611) := X"8FC200A8";
        ram_buffer(45612) := X"8FC4008C";
        ram_buffer(45613) := X"00000000";
        ram_buffer(45614) := X"3085000F";
        ram_buffer(45615) := X"3C04100D";
        ram_buffer(45616) := X"000528C0";
        ram_buffer(45617) := X"2484A938";
        ram_buffer(45618) := X"00A42021";
        ram_buffer(45619) := X"8C850004";
        ram_buffer(45620) := X"8C840000";
        ram_buffer(45621) := X"00A03821";
        ram_buffer(45622) := X"00803021";
        ram_buffer(45623) := X"00602821";
        ram_buffer(45624) := X"00402021";
        ram_buffer(45625) := X"0C03174A";
        ram_buffer(45626) := X"00000000";
        ram_buffer(45627) := X"AFC300AC";
        ram_buffer(45628) := X"AFC200A8";
        ram_buffer(45629) := X"8FC2008C";
        ram_buffer(45630) := X"00000000";
        ram_buffer(45631) := X"00021103";
        ram_buffer(45632) := X"AFC20034";
        ram_buffer(45633) := X"10000024";
        ram_buffer(45634) := X"00000000";
        ram_buffer(45635) := X"8FC20034";
        ram_buffer(45636) := X"00000000";
        ram_buffer(45637) := X"30420001";
        ram_buffer(45638) := X"10400017";
        ram_buffer(45639) := X"00000000";
        ram_buffer(45640) := X"8FC20028";
        ram_buffer(45641) := X"00000000";
        ram_buffer(45642) := X"24420001";
        ram_buffer(45643) := X"AFC20028";
        ram_buffer(45644) := X"8FC300AC";
        ram_buffer(45645) := X"8FC200A8";
        ram_buffer(45646) := X"3C04100D";
        ram_buffer(45647) := X"8FC50024";
        ram_buffer(45648) := X"00000000";
        ram_buffer(45649) := X"000528C0";
        ram_buffer(45650) := X"2484AA00";
        ram_buffer(45651) := X"00A42021";
        ram_buffer(45652) := X"8C850004";
        ram_buffer(45653) := X"8C840000";
        ram_buffer(45654) := X"00A03821";
        ram_buffer(45655) := X"00803021";
        ram_buffer(45656) := X"00602821";
        ram_buffer(45657) := X"00402021";
        ram_buffer(45658) := X"0C03174A";
        ram_buffer(45659) := X"00000000";
        ram_buffer(45660) := X"AFC300AC";
        ram_buffer(45661) := X"AFC200A8";
        ram_buffer(45662) := X"8FC20034";
        ram_buffer(45663) := X"00000000";
        ram_buffer(45664) := X"00021043";
        ram_buffer(45665) := X"AFC20034";
        ram_buffer(45666) := X"8FC20024";
        ram_buffer(45667) := X"00000000";
        ram_buffer(45668) := X"24420001";
        ram_buffer(45669) := X"AFC20024";
        ram_buffer(45670) := X"8FC20034";
        ram_buffer(45671) := X"00000000";
        ram_buffer(45672) := X"1440FFDA";
        ram_buffer(45673) := X"00000000";
        ram_buffer(45674) := X"8FC2003C";
        ram_buffer(45675) := X"00000000";
        ram_buffer(45676) := X"10400028";
        ram_buffer(45677) := X"00000000";
        ram_buffer(45678) := X"8FC300AC";
        ram_buffer(45679) := X"8FC200A8";
        ram_buffer(45680) := X"8F8780FC";
        ram_buffer(45681) := X"8F8680F8";
        ram_buffer(45682) := X"00602821";
        ram_buffer(45683) := X"00402021";
        ram_buffer(45684) := X"0C0316F7";
        ram_buffer(45685) := X"00000000";
        ram_buffer(45686) := X"0441001E";
        ram_buffer(45687) := X"00000000";
        ram_buffer(45688) := X"8FC2002C";
        ram_buffer(45689) := X"00000000";
        ram_buffer(45690) := X"1840001A";
        ram_buffer(45691) := X"00000000";
        ram_buffer(45692) := X"8FC20030";
        ram_buffer(45693) := X"00000000";
        ram_buffer(45694) := X"18400156";
        ram_buffer(45695) := X"00000000";
        ram_buffer(45696) := X"8FC20030";
        ram_buffer(45697) := X"00000000";
        ram_buffer(45698) := X"AFC2002C";
        ram_buffer(45699) := X"8FC20038";
        ram_buffer(45700) := X"00000000";
        ram_buffer(45701) := X"2442FFFF";
        ram_buffer(45702) := X"AFC20038";
        ram_buffer(45703) := X"8FC300AC";
        ram_buffer(45704) := X"8FC200A8";
        ram_buffer(45705) := X"8F878104";
        ram_buffer(45706) := X"8F868100";
        ram_buffer(45707) := X"00602821";
        ram_buffer(45708) := X"00402021";
        ram_buffer(45709) := X"0C03174A";
        ram_buffer(45710) := X"00000000";
        ram_buffer(45711) := X"AFC300AC";
        ram_buffer(45712) := X"AFC200A8";
        ram_buffer(45713) := X"8FC20028";
        ram_buffer(45714) := X"00000000";
        ram_buffer(45715) := X"24420001";
        ram_buffer(45716) := X"AFC20028";
        ram_buffer(45717) := X"8FC40028";
        ram_buffer(45718) := X"0C031B7C";
        ram_buffer(45719) := X"00000000";
        ram_buffer(45720) := X"00602821";
        ram_buffer(45721) := X"00402021";
        ram_buffer(45722) := X"8FC300AC";
        ram_buffer(45723) := X"8FC200A8";
        ram_buffer(45724) := X"00603821";
        ram_buffer(45725) := X"00403021";
        ram_buffer(45726) := X"0C03174A";
        ram_buffer(45727) := X"00000000";
        ram_buffer(45728) := X"8F87810C";
        ram_buffer(45729) := X"8F868108";
        ram_buffer(45730) := X"00602821";
        ram_buffer(45731) := X"00402021";
        ram_buffer(45732) := X"0C0311FC";
        ram_buffer(45733) := X"00000000";
        ram_buffer(45734) := X"AFC300BC";
        ram_buffer(45735) := X"AFC200B8";
        ram_buffer(45736) := X"8FC300B8";
        ram_buffer(45737) := X"3C02FCC0";
        ram_buffer(45738) := X"00621021";
        ram_buffer(45739) := X"AFC200B8";
        ram_buffer(45740) := X"8FC2002C";
        ram_buffer(45741) := X"00000000";
        ram_buffer(45742) := X"1440002A";
        ram_buffer(45743) := X"00000000";
        ram_buffer(45744) := X"AFC00068";
        ram_buffer(45745) := X"8FC20068";
        ram_buffer(45746) := X"00000000";
        ram_buffer(45747) := X"AFC2006C";
        ram_buffer(45748) := X"8FC300AC";
        ram_buffer(45749) := X"8FC200A8";
        ram_buffer(45750) := X"8F878114";
        ram_buffer(45751) := X"8F868110";
        ram_buffer(45752) := X"00602821";
        ram_buffer(45753) := X"00402021";
        ram_buffer(45754) := X"0C0318D3";
        ram_buffer(45755) := X"00000000";
        ram_buffer(45756) := X"AFC300AC";
        ram_buffer(45757) := X"AFC200A8";
        ram_buffer(45758) := X"8FC300AC";
        ram_buffer(45759) := X"8FC200A8";
        ram_buffer(45760) := X"8FC500BC";
        ram_buffer(45761) := X"8FC400B8";
        ram_buffer(45762) := X"00A03821";
        ram_buffer(45763) := X"00803021";
        ram_buffer(45764) := X"00602821";
        ram_buffer(45765) := X"00402021";
        ram_buffer(45766) := X"0C0316AB";
        ram_buffer(45767) := X"00000000";
        ram_buffer(45768) := X"1C40038C";
        ram_buffer(45769) := X"00000000";
        ram_buffer(45770) := X"8FC500AC";
        ram_buffer(45771) := X"8FC400A8";
        ram_buffer(45772) := X"8FC300BC";
        ram_buffer(45773) := X"8FC200B8";
        ram_buffer(45774) := X"3C068000";
        ram_buffer(45775) := X"00468026";
        ram_buffer(45776) := X"00608821";
        ram_buffer(45777) := X"02203821";
        ram_buffer(45778) := X"02003021";
        ram_buffer(45779) := X"0C0316F7";
        ram_buffer(45780) := X"00000000";
        ram_buffer(45781) := X"04400378";
        ram_buffer(45782) := X"00000000";
        ram_buffer(45783) := X"10000101";
        ram_buffer(45784) := X"00000000";
        ram_buffer(45785) := X"8FC20040";
        ram_buffer(45786) := X"00000000";
        ram_buffer(45787) := X"10400079";
        ram_buffer(45788) := X"00000000";
        ram_buffer(45789) := X"8FC2002C";
        ram_buffer(45790) := X"00000000";
        ram_buffer(45791) := X"2443FFFF";
        ram_buffer(45792) := X"3C02100D";
        ram_buffer(45793) := X"000318C0";
        ram_buffer(45794) := X"2442A938";
        ram_buffer(45795) := X"00621021";
        ram_buffer(45796) := X"8C430004";
        ram_buffer(45797) := X"8C420000";
        ram_buffer(45798) := X"00603821";
        ram_buffer(45799) := X"00403021";
        ram_buffer(45800) := X"8F85811C";
        ram_buffer(45801) := X"8F848118";
        ram_buffer(45802) := X"0C03144F";
        ram_buffer(45803) := X"00000000";
        ram_buffer(45804) := X"00602821";
        ram_buffer(45805) := X"00402021";
        ram_buffer(45806) := X"8FC300BC";
        ram_buffer(45807) := X"8FC200B8";
        ram_buffer(45808) := X"00603821";
        ram_buffer(45809) := X"00403021";
        ram_buffer(45810) := X"0C0318D3";
        ram_buffer(45811) := X"00000000";
        ram_buffer(45812) := X"AFC300BC";
        ram_buffer(45813) := X"AFC200B8";
        ram_buffer(45814) := X"AFC00024";
        ram_buffer(45815) := X"8FC300AC";
        ram_buffer(45816) := X"8FC200A8";
        ram_buffer(45817) := X"00602821";
        ram_buffer(45818) := X"00402021";
        ram_buffer(45819) := X"0C031B37";
        ram_buffer(45820) := X"00000000";
        ram_buffer(45821) := X"AFC20090";
        ram_buffer(45822) := X"8FD100AC";
        ram_buffer(45823) := X"8FD000A8";
        ram_buffer(45824) := X"8FC40090";
        ram_buffer(45825) := X"0C031B7C";
        ram_buffer(45826) := X"00000000";
        ram_buffer(45827) := X"00603821";
        ram_buffer(45828) := X"00403021";
        ram_buffer(45829) := X"02202821";
        ram_buffer(45830) := X"02002021";
        ram_buffer(45831) := X"0C0318D3";
        ram_buffer(45832) := X"00000000";
        ram_buffer(45833) := X"AFC300AC";
        ram_buffer(45834) := X"AFC200A8";
        ram_buffer(45835) := X"8FC20078";
        ram_buffer(45836) := X"00000000";
        ram_buffer(45837) := X"24430001";
        ram_buffer(45838) := X"AFC30078";
        ram_buffer(45839) := X"8FC30090";
        ram_buffer(45840) := X"00000000";
        ram_buffer(45841) := X"306300FF";
        ram_buffer(45842) := X"24630030";
        ram_buffer(45843) := X"306300FF";
        ram_buffer(45844) := X"00031E00";
        ram_buffer(45845) := X"00031E03";
        ram_buffer(45846) := X"A0430000";
        ram_buffer(45847) := X"8FC300AC";
        ram_buffer(45848) := X"8FC200A8";
        ram_buffer(45849) := X"8FC500BC";
        ram_buffer(45850) := X"8FC400B8";
        ram_buffer(45851) := X"00A03821";
        ram_buffer(45852) := X"00803021";
        ram_buffer(45853) := X"00602821";
        ram_buffer(45854) := X"00402021";
        ram_buffer(45855) := X"0C0316F7";
        ram_buffer(45856) := X"00000000";
        ram_buffer(45857) := X"044004EF";
        ram_buffer(45858) := X"00000000";
        ram_buffer(45859) := X"8FC300AC";
        ram_buffer(45860) := X"8FC200A8";
        ram_buffer(45861) := X"00603821";
        ram_buffer(45862) := X"00403021";
        ram_buffer(45863) := X"8F8580FC";
        ram_buffer(45864) := X"8F8480F8";
        ram_buffer(45865) := X"0C0318D3";
        ram_buffer(45866) := X"00000000";
        ram_buffer(45867) := X"00602821";
        ram_buffer(45868) := X"00402021";
        ram_buffer(45869) := X"8FC300BC";
        ram_buffer(45870) := X"8FC200B8";
        ram_buffer(45871) := X"00603821";
        ram_buffer(45872) := X"00403021";
        ram_buffer(45873) := X"0C0316F7";
        ram_buffer(45874) := X"00000000";
        ram_buffer(45875) := X"04400141";
        ram_buffer(45876) := X"00000000";
        ram_buffer(45877) := X"8FC20024";
        ram_buffer(45878) := X"00000000";
        ram_buffer(45879) := X"24420001";
        ram_buffer(45880) := X"AFC20024";
        ram_buffer(45881) := X"8FC30024";
        ram_buffer(45882) := X"8FC2002C";
        ram_buffer(45883) := X"00000000";
        ram_buffer(45884) := X"0062102A";
        ram_buffer(45885) := X"1040009A";
        ram_buffer(45886) := X"00000000";
        ram_buffer(45887) := X"8FC300BC";
        ram_buffer(45888) := X"8FC200B8";
        ram_buffer(45889) := X"8F878104";
        ram_buffer(45890) := X"8F868100";
        ram_buffer(45891) := X"00602821";
        ram_buffer(45892) := X"00402021";
        ram_buffer(45893) := X"0C03174A";
        ram_buffer(45894) := X"00000000";
        ram_buffer(45895) := X"AFC300BC";
        ram_buffer(45896) := X"AFC200B8";
        ram_buffer(45897) := X"8FC300AC";
        ram_buffer(45898) := X"8FC200A8";
        ram_buffer(45899) := X"8F878104";
        ram_buffer(45900) := X"8F868100";
        ram_buffer(45901) := X"00602821";
        ram_buffer(45902) := X"00402021";
        ram_buffer(45903) := X"0C03174A";
        ram_buffer(45904) := X"00000000";
        ram_buffer(45905) := X"AFC300AC";
        ram_buffer(45906) := X"AFC200A8";
        ram_buffer(45907) := X"1000FFA3";
        ram_buffer(45908) := X"00000000";
        ram_buffer(45909) := X"8FC300BC";
        ram_buffer(45910) := X"8FC200B8";
        ram_buffer(45911) := X"8FC4002C";
        ram_buffer(45912) := X"00000000";
        ram_buffer(45913) := X"2485FFFF";
        ram_buffer(45914) := X"3C04100D";
        ram_buffer(45915) := X"000528C0";
        ram_buffer(45916) := X"2484A938";
        ram_buffer(45917) := X"00A42021";
        ram_buffer(45918) := X"8C850004";
        ram_buffer(45919) := X"8C840000";
        ram_buffer(45920) := X"00A03821";
        ram_buffer(45921) := X"00803021";
        ram_buffer(45922) := X"00602821";
        ram_buffer(45923) := X"00402021";
        ram_buffer(45924) := X"0C03174A";
        ram_buffer(45925) := X"00000000";
        ram_buffer(45926) := X"AFC300BC";
        ram_buffer(45927) := X"AFC200B8";
        ram_buffer(45928) := X"24020001";
        ram_buffer(45929) := X"AFC20024";
        ram_buffer(45930) := X"8FC300AC";
        ram_buffer(45931) := X"8FC200A8";
        ram_buffer(45932) := X"00602821";
        ram_buffer(45933) := X"00402021";
        ram_buffer(45934) := X"0C031B37";
        ram_buffer(45935) := X"00000000";
        ram_buffer(45936) := X"AFC20090";
        ram_buffer(45937) := X"8FD100AC";
        ram_buffer(45938) := X"8FD000A8";
        ram_buffer(45939) := X"8FC40090";
        ram_buffer(45940) := X"0C031B7C";
        ram_buffer(45941) := X"00000000";
        ram_buffer(45942) := X"00603821";
        ram_buffer(45943) := X"00403021";
        ram_buffer(45944) := X"02202821";
        ram_buffer(45945) := X"02002021";
        ram_buffer(45946) := X"0C0318D3";
        ram_buffer(45947) := X"00000000";
        ram_buffer(45948) := X"AFC300AC";
        ram_buffer(45949) := X"AFC200A8";
        ram_buffer(45950) := X"8FC20078";
        ram_buffer(45951) := X"00000000";
        ram_buffer(45952) := X"24430001";
        ram_buffer(45953) := X"AFC30078";
        ram_buffer(45954) := X"8FC30090";
        ram_buffer(45955) := X"00000000";
        ram_buffer(45956) := X"306300FF";
        ram_buffer(45957) := X"24630030";
        ram_buffer(45958) := X"306300FF";
        ram_buffer(45959) := X"00031E00";
        ram_buffer(45960) := X"00031E03";
        ram_buffer(45961) := X"A0430000";
        ram_buffer(45962) := X"8FC30024";
        ram_buffer(45963) := X"8FC2002C";
        ram_buffer(45964) := X"00000000";
        ram_buffer(45965) := X"14620037";
        ram_buffer(45966) := X"00000000";
        ram_buffer(45967) := X"8FD100AC";
        ram_buffer(45968) := X"8FD000A8";
        ram_buffer(45969) := X"8FC300BC";
        ram_buffer(45970) := X"8FC200B8";
        ram_buffer(45971) := X"8F87811C";
        ram_buffer(45972) := X"8F868118";
        ram_buffer(45973) := X"00602821";
        ram_buffer(45974) := X"00402021";
        ram_buffer(45975) := X"0C0311FC";
        ram_buffer(45976) := X"00000000";
        ram_buffer(45977) := X"00603821";
        ram_buffer(45978) := X"00403021";
        ram_buffer(45979) := X"02202821";
        ram_buffer(45980) := X"02002021";
        ram_buffer(45981) := X"0C0316AB";
        ram_buffer(45982) := X"00000000";
        ram_buffer(45983) := X"1C4000D8";
        ram_buffer(45984) := X"00000000";
        ram_buffer(45985) := X"8FD100AC";
        ram_buffer(45986) := X"8FD000A8";
        ram_buffer(45987) := X"8FC300BC";
        ram_buffer(45988) := X"8FC200B8";
        ram_buffer(45989) := X"00603821";
        ram_buffer(45990) := X"00403021";
        ram_buffer(45991) := X"8F85811C";
        ram_buffer(45992) := X"8F848118";
        ram_buffer(45993) := X"0C0318D3";
        ram_buffer(45994) := X"00000000";
        ram_buffer(45995) := X"00603821";
        ram_buffer(45996) := X"00403021";
        ram_buffer(45997) := X"02202821";
        ram_buffer(45998) := X"02002021";
        ram_buffer(45999) := X"0C0316F7";
        ram_buffer(46000) := X"00000000";
        ram_buffer(46001) := X"04400003";
        ram_buffer(46002) := X"00000000";
        ram_buffer(46003) := X"10000025";
        ram_buffer(46004) := X"00000000";
        ram_buffer(46005) := X"8FC20078";
        ram_buffer(46006) := X"00000000";
        ram_buffer(46007) := X"2442FFFF";
        ram_buffer(46008) := X"AFC20078";
        ram_buffer(46009) := X"8FC20078";
        ram_buffer(46010) := X"00000000";
        ram_buffer(46011) := X"80430000";
        ram_buffer(46012) := X"24020030";
        ram_buffer(46013) := X"1062FFF7";
        ram_buffer(46014) := X"00000000";
        ram_buffer(46015) := X"8FC20078";
        ram_buffer(46016) := X"00000000";
        ram_buffer(46017) := X"24420001";
        ram_buffer(46018) := X"AFC20078";
        ram_buffer(46019) := X"1000044E";
        ram_buffer(46020) := X"00000000";
        ram_buffer(46021) := X"8FC20024";
        ram_buffer(46022) := X"00000000";
        ram_buffer(46023) := X"24420001";
        ram_buffer(46024) := X"AFC20024";
        ram_buffer(46025) := X"8FC300AC";
        ram_buffer(46026) := X"8FC200A8";
        ram_buffer(46027) := X"8F878104";
        ram_buffer(46028) := X"8F868100";
        ram_buffer(46029) := X"00602821";
        ram_buffer(46030) := X"00402021";
        ram_buffer(46031) := X"0C03174A";
        ram_buffer(46032) := X"00000000";
        ram_buffer(46033) := X"AFC300AC";
        ram_buffer(46034) := X"AFC200A8";
        ram_buffer(46035) := X"1000FF96";
        ram_buffer(46036) := X"00000000";
        ram_buffer(46037) := X"00000000";
        ram_buffer(46038) := X"10000002";
        ram_buffer(46039) := X"00000000";
        ram_buffer(46040) := X"00000000";
        ram_buffer(46041) := X"8FC20080";
        ram_buffer(46042) := X"00000000";
        ram_buffer(46043) := X"AFC20078";
        ram_buffer(46044) := X"8FC300B4";
        ram_buffer(46045) := X"8FC200B0";
        ram_buffer(46046) := X"AFC300AC";
        ram_buffer(46047) := X"AFC200A8";
        ram_buffer(46048) := X"8FC20084";
        ram_buffer(46049) := X"00000000";
        ram_buffer(46050) := X"AFC20038";
        ram_buffer(46051) := X"8FC20088";
        ram_buffer(46052) := X"00000000";
        ram_buffer(46053) := X"AFC2002C";
        ram_buffer(46054) := X"8FC200A0";
        ram_buffer(46055) := X"00000000";
        ram_buffer(46056) := X"044000D8";
        ram_buffer(46057) := X"00000000";
        ram_buffer(46058) := X"8FC20038";
        ram_buffer(46059) := X"00000000";
        ram_buffer(46060) := X"2842000F";
        ram_buffer(46061) := X"104000D3";
        ram_buffer(46062) := X"00000000";
        ram_buffer(46063) := X"3C02100D";
        ram_buffer(46064) := X"8FC30038";
        ram_buffer(46065) := X"00000000";
        ram_buffer(46066) := X"000318C0";
        ram_buffer(46067) := X"2442A938";
        ram_buffer(46068) := X"00621021";
        ram_buffer(46069) := X"8C430004";
        ram_buffer(46070) := X"8C420000";
        ram_buffer(46071) := X"AFC30074";
        ram_buffer(46072) := X"AFC20070";
        ram_buffer(46073) := X"8FC200EC";
        ram_buffer(46074) := X"00000000";
        ram_buffer(46075) := X"0441001F";
        ram_buffer(46076) := X"00000000";
        ram_buffer(46077) := X"8FC2002C";
        ram_buffer(46078) := X"00000000";
        ram_buffer(46079) := X"1C40001B";
        ram_buffer(46080) := X"00000000";
        ram_buffer(46081) := X"AFC00068";
        ram_buffer(46082) := X"8FC20068";
        ram_buffer(46083) := X"00000000";
        ram_buffer(46084) := X"AFC2006C";
        ram_buffer(46085) := X"8FC2002C";
        ram_buffer(46086) := X"00000000";
        ram_buffer(46087) := X"04400247";
        ram_buffer(46088) := X"00000000";
        ram_buffer(46089) := X"8FD100AC";
        ram_buffer(46090) := X"8FD000A8";
        ram_buffer(46091) := X"8F878114";
        ram_buffer(46092) := X"8F868110";
        ram_buffer(46093) := X"8FC50074";
        ram_buffer(46094) := X"8FC40070";
        ram_buffer(46095) := X"0C03174A";
        ram_buffer(46096) := X"00000000";
        ram_buffer(46097) := X"00603821";
        ram_buffer(46098) := X"00403021";
        ram_buffer(46099) := X"02202821";
        ram_buffer(46100) := X"02002021";
        ram_buffer(46101) := X"0C0316F7";
        ram_buffer(46102) := X"00000000";
        ram_buffer(46103) := X"18400237";
        ram_buffer(46104) := X"00000000";
        ram_buffer(46105) := X"1000023C";
        ram_buffer(46106) := X"00000000";
        ram_buffer(46107) := X"24020001";
        ram_buffer(46108) := X"AFC20024";
        ram_buffer(46109) := X"8FC300AC";
        ram_buffer(46110) := X"8FC200A8";
        ram_buffer(46111) := X"8FC70074";
        ram_buffer(46112) := X"8FC60070";
        ram_buffer(46113) := X"00602821";
        ram_buffer(46114) := X"00402021";
        ram_buffer(46115) := X"0C03144F";
        ram_buffer(46116) := X"00000000";
        ram_buffer(46117) := X"00602821";
        ram_buffer(46118) := X"00402021";
        ram_buffer(46119) := X"0C031B37";
        ram_buffer(46120) := X"00000000";
        ram_buffer(46121) := X"AFC20090";
        ram_buffer(46122) := X"8FD100AC";
        ram_buffer(46123) := X"8FD000A8";
        ram_buffer(46124) := X"8FC40090";
        ram_buffer(46125) := X"0C031B7C";
        ram_buffer(46126) := X"00000000";
        ram_buffer(46127) := X"8FC70074";
        ram_buffer(46128) := X"8FC60070";
        ram_buffer(46129) := X"00602821";
        ram_buffer(46130) := X"00402021";
        ram_buffer(46131) := X"0C03174A";
        ram_buffer(46132) := X"00000000";
        ram_buffer(46133) := X"00603821";
        ram_buffer(46134) := X"00403021";
        ram_buffer(46135) := X"02202821";
        ram_buffer(46136) := X"02002021";
        ram_buffer(46137) := X"0C0318D3";
        ram_buffer(46138) := X"00000000";
        ram_buffer(46139) := X"AFC300AC";
        ram_buffer(46140) := X"AFC200A8";
        ram_buffer(46141) := X"8FC20078";
        ram_buffer(46142) := X"00000000";
        ram_buffer(46143) := X"24430001";
        ram_buffer(46144) := X"AFC30078";
        ram_buffer(46145) := X"8FC30090";
        ram_buffer(46146) := X"00000000";
        ram_buffer(46147) := X"306300FF";
        ram_buffer(46148) := X"24630030";
        ram_buffer(46149) := X"306300FF";
        ram_buffer(46150) := X"00031E00";
        ram_buffer(46151) := X"00031E03";
        ram_buffer(46152) := X"A0430000";
        ram_buffer(46153) := X"8FC30024";
        ram_buffer(46154) := X"8FC2002C";
        ram_buffer(46155) := X"00000000";
        ram_buffer(46156) := X"14620054";
        ram_buffer(46157) := X"00000000";
        ram_buffer(46158) := X"8FC300AC";
        ram_buffer(46159) := X"8FC200A8";
        ram_buffer(46160) := X"00603821";
        ram_buffer(46161) := X"00403021";
        ram_buffer(46162) := X"00602821";
        ram_buffer(46163) := X"00402021";
        ram_buffer(46164) := X"0C0311FC";
        ram_buffer(46165) := X"00000000";
        ram_buffer(46166) := X"AFC300AC";
        ram_buffer(46167) := X"AFC200A8";
        ram_buffer(46168) := X"8FC300AC";
        ram_buffer(46169) := X"8FC200A8";
        ram_buffer(46170) := X"8FC70074";
        ram_buffer(46171) := X"8FC60070";
        ram_buffer(46172) := X"00602821";
        ram_buffer(46173) := X"00402021";
        ram_buffer(46174) := X"0C0316AB";
        ram_buffer(46175) := X"00000000";
        ram_buffer(46176) := X"1C400028";
        ram_buffer(46177) := X"00000000";
        ram_buffer(46178) := X"8FC300AC";
        ram_buffer(46179) := X"8FC200A8";
        ram_buffer(46180) := X"8FC70074";
        ram_buffer(46181) := X"8FC60070";
        ram_buffer(46182) := X"00602821";
        ram_buffer(46183) := X"00402021";
        ram_buffer(46184) := X"0C03167F";
        ram_buffer(46185) := X"00000000";
        ram_buffer(46186) := X"10400003";
        ram_buffer(46187) := X"00000000";
        ram_buffer(46188) := X"1000004E";
        ram_buffer(46189) := X"00000000";
        ram_buffer(46190) := X"8FC20090";
        ram_buffer(46191) := X"00000000";
        ram_buffer(46192) := X"30420001";
        ram_buffer(46193) := X"10400049";
        ram_buffer(46194) := X"00000000";
        ram_buffer(46195) := X"10000015";
        ram_buffer(46196) := X"00000000";
        ram_buffer(46197) := X"00000000";
        ram_buffer(46198) := X"10000012";
        ram_buffer(46199) := X"00000000";
        ram_buffer(46200) := X"00000000";
        ram_buffer(46201) := X"1000000F";
        ram_buffer(46202) := X"00000000";
        ram_buffer(46203) := X"8FC30078";
        ram_buffer(46204) := X"8FC20080";
        ram_buffer(46205) := X"00000000";
        ram_buffer(46206) := X"1462000A";
        ram_buffer(46207) := X"00000000";
        ram_buffer(46208) := X"8FC20038";
        ram_buffer(46209) := X"00000000";
        ram_buffer(46210) := X"24420001";
        ram_buffer(46211) := X"AFC20038";
        ram_buffer(46212) := X"8FC20078";
        ram_buffer(46213) := X"24030030";
        ram_buffer(46214) := X"A0430000";
        ram_buffer(46215) := X"1000000B";
        ram_buffer(46216) := X"00000000";
        ram_buffer(46217) := X"8FC20078";
        ram_buffer(46218) := X"00000000";
        ram_buffer(46219) := X"2442FFFF";
        ram_buffer(46220) := X"AFC20078";
        ram_buffer(46221) := X"8FC20078";
        ram_buffer(46222) := X"00000000";
        ram_buffer(46223) := X"80430000";
        ram_buffer(46224) := X"24020039";
        ram_buffer(46225) := X"1062FFE9";
        ram_buffer(46226) := X"00000000";
        ram_buffer(46227) := X"8FC20078";
        ram_buffer(46228) := X"00000000";
        ram_buffer(46229) := X"24430001";
        ram_buffer(46230) := X"AFC30078";
        ram_buffer(46231) := X"80430000";
        ram_buffer(46232) := X"00000000";
        ram_buffer(46233) := X"306300FF";
        ram_buffer(46234) := X"24630001";
        ram_buffer(46235) := X"306300FF";
        ram_buffer(46236) := X"00031E00";
        ram_buffer(46237) := X"00031E03";
        ram_buffer(46238) := X"A0430000";
        ram_buffer(46239) := X"1000001B";
        ram_buffer(46240) := X"00000000";
        ram_buffer(46241) := X"8FC300AC";
        ram_buffer(46242) := X"8FC200A8";
        ram_buffer(46243) := X"8F878104";
        ram_buffer(46244) := X"8F868100";
        ram_buffer(46245) := X"00602821";
        ram_buffer(46246) := X"00402021";
        ram_buffer(46247) := X"0C03174A";
        ram_buffer(46248) := X"00000000";
        ram_buffer(46249) := X"AFC300AC";
        ram_buffer(46250) := X"AFC200A8";
        ram_buffer(46251) := X"8FC300AC";
        ram_buffer(46252) := X"8FC200A8";
        ram_buffer(46253) := X"00003821";
        ram_buffer(46254) := X"00003021";
        ram_buffer(46255) := X"00602821";
        ram_buffer(46256) := X"00402021";
        ram_buffer(46257) := X"0C03167F";
        ram_buffer(46258) := X"00000000";
        ram_buffer(46259) := X"1040000A";
        ram_buffer(46260) := X"00000000";
        ram_buffer(46261) := X"8FC20024";
        ram_buffer(46262) := X"00000000";
        ram_buffer(46263) := X"24420001";
        ram_buffer(46264) := X"AFC20024";
        ram_buffer(46265) := X"1000FF63";
        ram_buffer(46266) := X"00000000";
        ram_buffer(46267) := X"00000000";
        ram_buffer(46268) := X"10000355";
        ram_buffer(46269) := X"00000000";
        ram_buffer(46270) := X"00000000";
        ram_buffer(46271) := X"10000352";
        ram_buffer(46272) := X"00000000";
        ram_buffer(46273) := X"8FC20018";
        ram_buffer(46274) := X"00000000";
        ram_buffer(46275) := X"AFC20044";
        ram_buffer(46276) := X"8FC2001C";
        ram_buffer(46277) := X"00000000";
        ram_buffer(46278) := X"AFC20048";
        ram_buffer(46279) := X"AFC00064";
        ram_buffer(46280) := X"8FC20064";
        ram_buffer(46281) := X"00000000";
        ram_buffer(46282) := X"AFC20068";
        ram_buffer(46283) := X"8FC20040";
        ram_buffer(46284) := X"00000000";
        ram_buffer(46285) := X"10400052";
        ram_buffer(46286) := X"00000000";
        ram_buffer(46287) := X"8FC200E8";
        ram_buffer(46288) := X"00000000";
        ram_buffer(46289) := X"28420002";
        ram_buffer(46290) := X"10400010";
        ram_buffer(46291) := X"00000000";
        ram_buffer(46292) := X"8FC2005C";
        ram_buffer(46293) := X"00000000";
        ram_buffer(46294) := X"10400006";
        ram_buffer(46295) := X"00000000";
        ram_buffer(46296) := X"8FC200A0";
        ram_buffer(46297) := X"00000000";
        ram_buffer(46298) := X"24420433";
        ram_buffer(46299) := X"10000004";
        ram_buffer(46300) := X"00000000";
        ram_buffer(46301) := X"8FC2009C";
        ram_buffer(46302) := X"24030036";
        ram_buffer(46303) := X"00621023";
        ram_buffer(46304) := X"AFC20024";
        ram_buffer(46305) := X"1000002F";
        ram_buffer(46306) := X"00000000";
        ram_buffer(46307) := X"8FC2002C";
        ram_buffer(46308) := X"00000000";
        ram_buffer(46309) := X"2442FFFF";
        ram_buffer(46310) := X"AFC20034";
        ram_buffer(46311) := X"8FC30048";
        ram_buffer(46312) := X"8FC20034";
        ram_buffer(46313) := X"00000000";
        ram_buffer(46314) := X"0062102A";
        ram_buffer(46315) := X"14400008";
        ram_buffer(46316) := X"00000000";
        ram_buffer(46317) := X"8FC30048";
        ram_buffer(46318) := X"8FC20034";
        ram_buffer(46319) := X"00000000";
        ram_buffer(46320) := X"00621023";
        ram_buffer(46321) := X"AFC20048";
        ram_buffer(46322) := X"10000011";
        ram_buffer(46323) := X"00000000";
        ram_buffer(46324) := X"8FC30034";
        ram_buffer(46325) := X"8FC20048";
        ram_buffer(46326) := X"00000000";
        ram_buffer(46327) := X"00621023";
        ram_buffer(46328) := X"AFC20034";
        ram_buffer(46329) := X"8FC20034";
        ram_buffer(46330) := X"8FC30050";
        ram_buffer(46331) := X"00000000";
        ram_buffer(46332) := X"00621021";
        ram_buffer(46333) := X"AFC20050";
        ram_buffer(46334) := X"8FC3001C";
        ram_buffer(46335) := X"8FC20034";
        ram_buffer(46336) := X"00000000";
        ram_buffer(46337) := X"00621021";
        ram_buffer(46338) := X"AFC2001C";
        ram_buffer(46339) := X"AFC00048";
        ram_buffer(46340) := X"8FC2002C";
        ram_buffer(46341) := X"00000000";
        ram_buffer(46342) := X"AFC20024";
        ram_buffer(46343) := X"8FC20024";
        ram_buffer(46344) := X"00000000";
        ram_buffer(46345) := X"04410007";
        ram_buffer(46346) := X"00000000";
        ram_buffer(46347) := X"8FC30044";
        ram_buffer(46348) := X"8FC20024";
        ram_buffer(46349) := X"00000000";
        ram_buffer(46350) := X"00621023";
        ram_buffer(46351) := X"AFC20044";
        ram_buffer(46352) := X"AFC00024";
        ram_buffer(46353) := X"8FC30018";
        ram_buffer(46354) := X"8FC20024";
        ram_buffer(46355) := X"00000000";
        ram_buffer(46356) := X"00621021";
        ram_buffer(46357) := X"AFC20018";
        ram_buffer(46358) := X"8FC3004C";
        ram_buffer(46359) := X"8FC20024";
        ram_buffer(46360) := X"00000000";
        ram_buffer(46361) := X"00621021";
        ram_buffer(46362) := X"AFC2004C";
        ram_buffer(46363) := X"24050001";
        ram_buffer(46364) := X"8FC400D8";
        ram_buffer(46365) := X"0C02BFBF";
        ram_buffer(46366) := X"00000000";
        ram_buffer(46367) := X"AFC20068";
        ram_buffer(46368) := X"8FC20044";
        ram_buffer(46369) := X"00000000";
        ram_buffer(46370) := X"1840001C";
        ram_buffer(46371) := X"00000000";
        ram_buffer(46372) := X"8FC2004C";
        ram_buffer(46373) := X"00000000";
        ram_buffer(46374) := X"18400018";
        ram_buffer(46375) := X"00000000";
        ram_buffer(46376) := X"8FC30044";
        ram_buffer(46377) := X"8FC2004C";
        ram_buffer(46378) := X"00000000";
        ram_buffer(46379) := X"0062202A";
        ram_buffer(46380) := X"10800002";
        ram_buffer(46381) := X"00000000";
        ram_buffer(46382) := X"00601021";
        ram_buffer(46383) := X"AFC20024";
        ram_buffer(46384) := X"8FC30018";
        ram_buffer(46385) := X"8FC20024";
        ram_buffer(46386) := X"00000000";
        ram_buffer(46387) := X"00621023";
        ram_buffer(46388) := X"AFC20018";
        ram_buffer(46389) := X"8FC30044";
        ram_buffer(46390) := X"8FC20024";
        ram_buffer(46391) := X"00000000";
        ram_buffer(46392) := X"00621023";
        ram_buffer(46393) := X"AFC20044";
        ram_buffer(46394) := X"8FC3004C";
        ram_buffer(46395) := X"8FC20024";
        ram_buffer(46396) := X"00000000";
        ram_buffer(46397) := X"00621023";
        ram_buffer(46398) := X"AFC2004C";
        ram_buffer(46399) := X"8FC2001C";
        ram_buffer(46400) := X"00000000";
        ram_buffer(46401) := X"18400033";
        ram_buffer(46402) := X"00000000";
        ram_buffer(46403) := X"8FC20040";
        ram_buffer(46404) := X"00000000";
        ram_buffer(46405) := X"10400029";
        ram_buffer(46406) := X"00000000";
        ram_buffer(46407) := X"8FC20048";
        ram_buffer(46408) := X"00000000";
        ram_buffer(46409) := X"18400014";
        ram_buffer(46410) := X"00000000";
        ram_buffer(46411) := X"8FC60048";
        ram_buffer(46412) := X"8FC50068";
        ram_buffer(46413) := X"8FC400D8";
        ram_buffer(46414) := X"0C02C138";
        ram_buffer(46415) := X"00000000";
        ram_buffer(46416) := X"AFC20068";
        ram_buffer(46417) := X"8FC60060";
        ram_buffer(46418) := X"8FC50068";
        ram_buffer(46419) := X"8FC400D8";
        ram_buffer(46420) := X"0C02BFD8";
        ram_buffer(46421) := X"00000000";
        ram_buffer(46422) := X"AFC20094";
        ram_buffer(46423) := X"8FC50060";
        ram_buffer(46424) := X"8FC400D8";
        ram_buffer(46425) := X"0C02BE10";
        ram_buffer(46426) := X"00000000";
        ram_buffer(46427) := X"8FC20094";
        ram_buffer(46428) := X"00000000";
        ram_buffer(46429) := X"AFC20060";
        ram_buffer(46430) := X"8FC3001C";
        ram_buffer(46431) := X"8FC20048";
        ram_buffer(46432) := X"00000000";
        ram_buffer(46433) := X"00621023";
        ram_buffer(46434) := X"AFC20034";
        ram_buffer(46435) := X"8FC20034";
        ram_buffer(46436) := X"00000000";
        ram_buffer(46437) := X"1040000F";
        ram_buffer(46438) := X"00000000";
        ram_buffer(46439) := X"8FC60034";
        ram_buffer(46440) := X"8FC50060";
        ram_buffer(46441) := X"8FC400D8";
        ram_buffer(46442) := X"0C02C138";
        ram_buffer(46443) := X"00000000";
        ram_buffer(46444) := X"AFC20060";
        ram_buffer(46445) := X"10000007";
        ram_buffer(46446) := X"00000000";
        ram_buffer(46447) := X"8FC6001C";
        ram_buffer(46448) := X"8FC50060";
        ram_buffer(46449) := X"8FC400D8";
        ram_buffer(46450) := X"0C02C138";
        ram_buffer(46451) := X"00000000";
        ram_buffer(46452) := X"AFC20060";
        ram_buffer(46453) := X"24050001";
        ram_buffer(46454) := X"8FC400D8";
        ram_buffer(46455) := X"0C02BFBF";
        ram_buffer(46456) := X"00000000";
        ram_buffer(46457) := X"AFC2006C";
        ram_buffer(46458) := X"8FC20050";
        ram_buffer(46459) := X"00000000";
        ram_buffer(46460) := X"18400007";
        ram_buffer(46461) := X"00000000";
        ram_buffer(46462) := X"8FC60050";
        ram_buffer(46463) := X"8FC5006C";
        ram_buffer(46464) := X"8FC400D8";
        ram_buffer(46465) := X"0C02C138";
        ram_buffer(46466) := X"00000000";
        ram_buffer(46467) := X"AFC2006C";
        ram_buffer(46468) := X"AFC00054";
        ram_buffer(46469) := X"8FC200E8";
        ram_buffer(46470) := X"00000000";
        ram_buffer(46471) := X"28420002";
        ram_buffer(46472) := X"1040001A";
        ram_buffer(46473) := X"00000000";
        ram_buffer(46474) := X"8FC200AC";
        ram_buffer(46475) := X"00000000";
        ram_buffer(46476) := X"14400016";
        ram_buffer(46477) := X"00000000";
        ram_buffer(46478) := X"8FC300A8";
        ram_buffer(46479) := X"3C02000F";
        ram_buffer(46480) := X"3442FFFF";
        ram_buffer(46481) := X"00621024";
        ram_buffer(46482) := X"14400010";
        ram_buffer(46483) := X"00000000";
        ram_buffer(46484) := X"8FC300A8";
        ram_buffer(46485) := X"3C027FF0";
        ram_buffer(46486) := X"00621024";
        ram_buffer(46487) := X"1040000B";
        ram_buffer(46488) := X"00000000";
        ram_buffer(46489) := X"8FC20018";
        ram_buffer(46490) := X"00000000";
        ram_buffer(46491) := X"24420001";
        ram_buffer(46492) := X"AFC20018";
        ram_buffer(46493) := X"8FC2004C";
        ram_buffer(46494) := X"00000000";
        ram_buffer(46495) := X"24420001";
        ram_buffer(46496) := X"AFC2004C";
        ram_buffer(46497) := X"24020001";
        ram_buffer(46498) := X"AFC20054";
        ram_buffer(46499) := X"8FC20050";
        ram_buffer(46500) := X"00000000";
        ram_buffer(46501) := X"10400014";
        ram_buffer(46502) := X"00000000";
        ram_buffer(46503) := X"8FC2006C";
        ram_buffer(46504) := X"00000000";
        ram_buffer(46505) := X"8C420010";
        ram_buffer(46506) := X"00000000";
        ram_buffer(46507) := X"2442FFFF";
        ram_buffer(46508) := X"8FC3006C";
        ram_buffer(46509) := X"24420004";
        ram_buffer(46510) := X"00021080";
        ram_buffer(46511) := X"00621021";
        ram_buffer(46512) := X"8C420004";
        ram_buffer(46513) := X"00000000";
        ram_buffer(46514) := X"00402021";
        ram_buffer(46515) := X"0C02BF41";
        ram_buffer(46516) := X"00000000";
        ram_buffer(46517) := X"00401821";
        ram_buffer(46518) := X"24020020";
        ram_buffer(46519) := X"00431023";
        ram_buffer(46520) := X"10000002";
        ram_buffer(46521) := X"00000000";
        ram_buffer(46522) := X"24020001";
        ram_buffer(46523) := X"8FC3004C";
        ram_buffer(46524) := X"00000000";
        ram_buffer(46525) := X"00431021";
        ram_buffer(46526) := X"3042001F";
        ram_buffer(46527) := X"AFC20024";
        ram_buffer(46528) := X"8FC20024";
        ram_buffer(46529) := X"00000000";
        ram_buffer(46530) := X"10400006";
        ram_buffer(46531) := X"00000000";
        ram_buffer(46532) := X"24030020";
        ram_buffer(46533) := X"8FC20024";
        ram_buffer(46534) := X"00000000";
        ram_buffer(46535) := X"00621023";
        ram_buffer(46536) := X"AFC20024";
        ram_buffer(46537) := X"8FC20024";
        ram_buffer(46538) := X"00000000";
        ram_buffer(46539) := X"28420005";
        ram_buffer(46540) := X"14400016";
        ram_buffer(46541) := X"00000000";
        ram_buffer(46542) := X"8FC20024";
        ram_buffer(46543) := X"00000000";
        ram_buffer(46544) := X"2442FFFC";
        ram_buffer(46545) := X"AFC20024";
        ram_buffer(46546) := X"8FC30018";
        ram_buffer(46547) := X"8FC20024";
        ram_buffer(46548) := X"00000000";
        ram_buffer(46549) := X"00621021";
        ram_buffer(46550) := X"AFC20018";
        ram_buffer(46551) := X"8FC30044";
        ram_buffer(46552) := X"8FC20024";
        ram_buffer(46553) := X"00000000";
        ram_buffer(46554) := X"00621021";
        ram_buffer(46555) := X"AFC20044";
        ram_buffer(46556) := X"8FC3004C";
        ram_buffer(46557) := X"8FC20024";
        ram_buffer(46558) := X"00000000";
        ram_buffer(46559) := X"00621021";
        ram_buffer(46560) := X"AFC2004C";
        ram_buffer(46561) := X"10000019";
        ram_buffer(46562) := X"00000000";
        ram_buffer(46563) := X"8FC20024";
        ram_buffer(46564) := X"00000000";
        ram_buffer(46565) := X"28420004";
        ram_buffer(46566) := X"10400014";
        ram_buffer(46567) := X"00000000";
        ram_buffer(46568) := X"8FC20024";
        ram_buffer(46569) := X"00000000";
        ram_buffer(46570) := X"2442001C";
        ram_buffer(46571) := X"AFC20024";
        ram_buffer(46572) := X"8FC30018";
        ram_buffer(46573) := X"8FC20024";
        ram_buffer(46574) := X"00000000";
        ram_buffer(46575) := X"00621021";
        ram_buffer(46576) := X"AFC20018";
        ram_buffer(46577) := X"8FC30044";
        ram_buffer(46578) := X"8FC20024";
        ram_buffer(46579) := X"00000000";
        ram_buffer(46580) := X"00621021";
        ram_buffer(46581) := X"AFC20044";
        ram_buffer(46582) := X"8FC3004C";
        ram_buffer(46583) := X"8FC20024";
        ram_buffer(46584) := X"00000000";
        ram_buffer(46585) := X"00621021";
        ram_buffer(46586) := X"AFC2004C";
        ram_buffer(46587) := X"8FC20018";
        ram_buffer(46588) := X"00000000";
        ram_buffer(46589) := X"18400007";
        ram_buffer(46590) := X"00000000";
        ram_buffer(46591) := X"8FC60018";
        ram_buffer(46592) := X"8FC50060";
        ram_buffer(46593) := X"8FC400D8";
        ram_buffer(46594) := X"0C02C1BB";
        ram_buffer(46595) := X"00000000";
        ram_buffer(46596) := X"AFC20060";
        ram_buffer(46597) := X"8FC2004C";
        ram_buffer(46598) := X"00000000";
        ram_buffer(46599) := X"18400007";
        ram_buffer(46600) := X"00000000";
        ram_buffer(46601) := X"8FC6004C";
        ram_buffer(46602) := X"8FC5006C";
        ram_buffer(46603) := X"8FC400D8";
        ram_buffer(46604) := X"0C02C1BB";
        ram_buffer(46605) := X"00000000";
        ram_buffer(46606) := X"AFC2006C";
        ram_buffer(46607) := X"8FC2003C";
        ram_buffer(46608) := X"00000000";
        ram_buffer(46609) := X"10400020";
        ram_buffer(46610) := X"00000000";
        ram_buffer(46611) := X"8FC5006C";
        ram_buffer(46612) := X"8FC40060";
        ram_buffer(46613) := X"0C02C26D";
        ram_buffer(46614) := X"00000000";
        ram_buffer(46615) := X"0441001A";
        ram_buffer(46616) := X"00000000";
        ram_buffer(46617) := X"8FC20038";
        ram_buffer(46618) := X"00000000";
        ram_buffer(46619) := X"2442FFFF";
        ram_buffer(46620) := X"AFC20038";
        ram_buffer(46621) := X"00003821";
        ram_buffer(46622) := X"2406000A";
        ram_buffer(46623) := X"8FC50060";
        ram_buffer(46624) := X"8FC400D8";
        ram_buffer(46625) := X"0C02BE38";
        ram_buffer(46626) := X"00000000";
        ram_buffer(46627) := X"AFC20060";
        ram_buffer(46628) := X"8FC20040";
        ram_buffer(46629) := X"00000000";
        ram_buffer(46630) := X"10400008";
        ram_buffer(46631) := X"00000000";
        ram_buffer(46632) := X"00003821";
        ram_buffer(46633) := X"2406000A";
        ram_buffer(46634) := X"8FC50068";
        ram_buffer(46635) := X"8FC400D8";
        ram_buffer(46636) := X"0C02BE38";
        ram_buffer(46637) := X"00000000";
        ram_buffer(46638) := X"AFC20068";
        ram_buffer(46639) := X"8FC20030";
        ram_buffer(46640) := X"00000000";
        ram_buffer(46641) := X"AFC2002C";
        ram_buffer(46642) := X"8FC2002C";
        ram_buffer(46643) := X"00000000";
        ram_buffer(46644) := X"1C40002D";
        ram_buffer(46645) := X"00000000";
        ram_buffer(46646) := X"8FC200E8";
        ram_buffer(46647) := X"00000000";
        ram_buffer(46648) := X"28420003";
        ram_buffer(46649) := X"14400028";
        ram_buffer(46650) := X"00000000";
        ram_buffer(46651) := X"8FC2002C";
        ram_buffer(46652) := X"00000000";
        ram_buffer(46653) := X"04400011";
        ram_buffer(46654) := X"00000000";
        ram_buffer(46655) := X"00003821";
        ram_buffer(46656) := X"24060005";
        ram_buffer(46657) := X"8FC5006C";
        ram_buffer(46658) := X"8FC400D8";
        ram_buffer(46659) := X"0C02BE38";
        ram_buffer(46660) := X"00000000";
        ram_buffer(46661) := X"AFC2006C";
        ram_buffer(46662) := X"8FC5006C";
        ram_buffer(46663) := X"8FC40060";
        ram_buffer(46664) := X"0C02C26D";
        ram_buffer(46665) := X"00000000";
        ram_buffer(46666) := X"1C40000B";
        ram_buffer(46667) := X"00000000";
        ram_buffer(46668) := X"10000002";
        ram_buffer(46669) := X"00000000";
        ram_buffer(46670) := X"00000000";
        ram_buffer(46671) := X"8FC200EC";
        ram_buffer(46672) := X"00000000";
        ram_buffer(46673) := X"00021027";
        ram_buffer(46674) := X"AFC20038";
        ram_buffer(46675) := X"100001A2";
        ram_buffer(46676) := X"00000000";
        ram_buffer(46677) := X"00000000";
        ram_buffer(46678) := X"8FC20078";
        ram_buffer(46679) := X"00000000";
        ram_buffer(46680) := X"24430001";
        ram_buffer(46681) := X"AFC30078";
        ram_buffer(46682) := X"24030031";
        ram_buffer(46683) := X"A0430000";
        ram_buffer(46684) := X"8FC20038";
        ram_buffer(46685) := X"00000000";
        ram_buffer(46686) := X"24420001";
        ram_buffer(46687) := X"AFC20038";
        ram_buffer(46688) := X"10000195";
        ram_buffer(46689) := X"00000000";
        ram_buffer(46690) := X"8FC20040";
        ram_buffer(46691) := X"00000000";
        ram_buffer(46692) := X"10400118";
        ram_buffer(46693) := X"00000000";
        ram_buffer(46694) := X"8FC20044";
        ram_buffer(46695) := X"00000000";
        ram_buffer(46696) := X"18400007";
        ram_buffer(46697) := X"00000000";
        ram_buffer(46698) := X"8FC60044";
        ram_buffer(46699) := X"8FC50068";
        ram_buffer(46700) := X"8FC400D8";
        ram_buffer(46701) := X"0C02C1BB";
        ram_buffer(46702) := X"00000000";
        ram_buffer(46703) := X"AFC20068";
        ram_buffer(46704) := X"8FC20068";
        ram_buffer(46705) := X"00000000";
        ram_buffer(46706) := X"AFC20064";
        ram_buffer(46707) := X"8FC20054";
        ram_buffer(46708) := X"00000000";
        ram_buffer(46709) := X"10400021";
        ram_buffer(46710) := X"00000000";
        ram_buffer(46711) := X"8FC20068";
        ram_buffer(46712) := X"00000000";
        ram_buffer(46713) := X"8C420004";
        ram_buffer(46714) := X"00000000";
        ram_buffer(46715) := X"00402821";
        ram_buffer(46716) := X"8FC400D8";
        ram_buffer(46717) := X"0C02BDA8";
        ram_buffer(46718) := X"00000000";
        ram_buffer(46719) := X"AFC20068";
        ram_buffer(46720) := X"8FC20068";
        ram_buffer(46721) := X"00000000";
        ram_buffer(46722) := X"2443000C";
        ram_buffer(46723) := X"8FC20064";
        ram_buffer(46724) := X"00000000";
        ram_buffer(46725) := X"2444000C";
        ram_buffer(46726) := X"8FC20064";
        ram_buffer(46727) := X"00000000";
        ram_buffer(46728) := X"8C420010";
        ram_buffer(46729) := X"00000000";
        ram_buffer(46730) := X"24420002";
        ram_buffer(46731) := X"00021080";
        ram_buffer(46732) := X"00403021";
        ram_buffer(46733) := X"00802821";
        ram_buffer(46734) := X"00602021";
        ram_buffer(46735) := X"0C027F93";
        ram_buffer(46736) := X"00000000";
        ram_buffer(46737) := X"24060001";
        ram_buffer(46738) := X"8FC50068";
        ram_buffer(46739) := X"8FC400D8";
        ram_buffer(46740) := X"0C02C1BB";
        ram_buffer(46741) := X"00000000";
        ram_buffer(46742) := X"AFC20068";
        ram_buffer(46743) := X"24020001";
        ram_buffer(46744) := X"AFC20024";
        ram_buffer(46745) := X"8FC5006C";
        ram_buffer(46746) := X"8FC40060";
        ram_buffer(46747) := X"0C02AE52";
        ram_buffer(46748) := X"00000000";
        ram_buffer(46749) := X"24420030";
        ram_buffer(46750) := X"AFC20020";
        ram_buffer(46751) := X"8FC50064";
        ram_buffer(46752) := X"8FC40060";
        ram_buffer(46753) := X"0C02C26D";
        ram_buffer(46754) := X"00000000";
        ram_buffer(46755) := X"AFC20034";
        ram_buffer(46756) := X"8FC60068";
        ram_buffer(46757) := X"8FC5006C";
        ram_buffer(46758) := X"8FC400D8";
        ram_buffer(46759) := X"0C02C2CE";
        ram_buffer(46760) := X"00000000";
        ram_buffer(46761) := X"AFC20098";
        ram_buffer(46762) := X"8FC20098";
        ram_buffer(46763) := X"00000000";
        ram_buffer(46764) := X"8C42000C";
        ram_buffer(46765) := X"00000000";
        ram_buffer(46766) := X"14400007";
        ram_buffer(46767) := X"00000000";
        ram_buffer(46768) := X"8FC50098";
        ram_buffer(46769) := X"8FC40060";
        ram_buffer(46770) := X"0C02C26D";
        ram_buffer(46771) := X"00000000";
        ram_buffer(46772) := X"10000002";
        ram_buffer(46773) := X"00000000";
        ram_buffer(46774) := X"24020001";
        ram_buffer(46775) := X"AFC2008C";
        ram_buffer(46776) := X"8FC50098";
        ram_buffer(46777) := X"8FC400D8";
        ram_buffer(46778) := X"0C02BE10";
        ram_buffer(46779) := X"00000000";
        ram_buffer(46780) := X"8FC2008C";
        ram_buffer(46781) := X"00000000";
        ram_buffer(46782) := X"14400021";
        ram_buffer(46783) := X"00000000";
        ram_buffer(46784) := X"8FC200E8";
        ram_buffer(46785) := X"00000000";
        ram_buffer(46786) := X"1440001D";
        ram_buffer(46787) := X"00000000";
        ram_buffer(46788) := X"8FC200AC";
        ram_buffer(46789) := X"00000000";
        ram_buffer(46790) := X"30420001";
        ram_buffer(46791) := X"14400018";
        ram_buffer(46792) := X"00000000";
        ram_buffer(46793) := X"8FC30020";
        ram_buffer(46794) := X"24020039";
        ram_buffer(46795) := X"1062005D";
        ram_buffer(46796) := X"00000000";
        ram_buffer(46797) := X"8FC20034";
        ram_buffer(46798) := X"00000000";
        ram_buffer(46799) := X"18400005";
        ram_buffer(46800) := X"00000000";
        ram_buffer(46801) := X"8FC20020";
        ram_buffer(46802) := X"00000000";
        ram_buffer(46803) := X"24420001";
        ram_buffer(46804) := X"AFC20020";
        ram_buffer(46805) := X"8FC20078";
        ram_buffer(46806) := X"00000000";
        ram_buffer(46807) := X"24430001";
        ram_buffer(46808) := X"AFC30078";
        ram_buffer(46809) := X"8FC30020";
        ram_buffer(46810) := X"00000000";
        ram_buffer(46811) := X"00031E00";
        ram_buffer(46812) := X"00031E03";
        ram_buffer(46813) := X"A0430000";
        ram_buffer(46814) := X"10000117";
        ram_buffer(46815) := X"00000000";
        ram_buffer(46816) := X"8FC20034";
        ram_buffer(46817) := X"00000000";
        ram_buffer(46818) := X"0440000E";
        ram_buffer(46819) := X"00000000";
        ram_buffer(46820) := X"8FC20034";
        ram_buffer(46821) := X"00000000";
        ram_buffer(46822) := X"14400038";
        ram_buffer(46823) := X"00000000";
        ram_buffer(46824) := X"8FC200E8";
        ram_buffer(46825) := X"00000000";
        ram_buffer(46826) := X"14400034";
        ram_buffer(46827) := X"00000000";
        ram_buffer(46828) := X"8FC200AC";
        ram_buffer(46829) := X"00000000";
        ram_buffer(46830) := X"30420001";
        ram_buffer(46831) := X"1440002F";
        ram_buffer(46832) := X"00000000";
        ram_buffer(46833) := X"8FC2008C";
        ram_buffer(46834) := X"00000000";
        ram_buffer(46835) := X"18400020";
        ram_buffer(46836) := X"00000000";
        ram_buffer(46837) := X"24060001";
        ram_buffer(46838) := X"8FC50060";
        ram_buffer(46839) := X"8FC400D8";
        ram_buffer(46840) := X"0C02C1BB";
        ram_buffer(46841) := X"00000000";
        ram_buffer(46842) := X"AFC20060";
        ram_buffer(46843) := X"8FC5006C";
        ram_buffer(46844) := X"8FC40060";
        ram_buffer(46845) := X"0C02C26D";
        ram_buffer(46846) := X"00000000";
        ram_buffer(46847) := X"AFC2008C";
        ram_buffer(46848) := X"8FC2008C";
        ram_buffer(46849) := X"00000000";
        ram_buffer(46850) := X"1C40000A";
        ram_buffer(46851) := X"00000000";
        ram_buffer(46852) := X"8FC2008C";
        ram_buffer(46853) := X"00000000";
        ram_buffer(46854) := X"1440000D";
        ram_buffer(46855) := X"00000000";
        ram_buffer(46856) := X"8FC20020";
        ram_buffer(46857) := X"00000000";
        ram_buffer(46858) := X"30420001";
        ram_buffer(46859) := X"10400008";
        ram_buffer(46860) := X"00000000";
        ram_buffer(46861) := X"8FC20020";
        ram_buffer(46862) := X"00000000";
        ram_buffer(46863) := X"24430001";
        ram_buffer(46864) := X"AFC30020";
        ram_buffer(46865) := X"24030039";
        ram_buffer(46866) := X"10430019";
        ram_buffer(46867) := X"00000000";
        ram_buffer(46868) := X"8FC20078";
        ram_buffer(46869) := X"00000000";
        ram_buffer(46870) := X"24430001";
        ram_buffer(46871) := X"AFC30078";
        ram_buffer(46872) := X"8FC30020";
        ram_buffer(46873) := X"00000000";
        ram_buffer(46874) := X"00031E00";
        ram_buffer(46875) := X"00031E03";
        ram_buffer(46876) := X"A0430000";
        ram_buffer(46877) := X"100000D8";
        ram_buffer(46878) := X"00000000";
        ram_buffer(46879) := X"8FC2008C";
        ram_buffer(46880) := X"00000000";
        ram_buffer(46881) := X"18400021";
        ram_buffer(46882) := X"00000000";
        ram_buffer(46883) := X"8FC30020";
        ram_buffer(46884) := X"24020039";
        ram_buffer(46885) := X"1462000F";
        ram_buffer(46886) := X"00000000";
        ram_buffer(46887) := X"10000005";
        ram_buffer(46888) := X"00000000";
        ram_buffer(46889) := X"00000000";
        ram_buffer(46890) := X"10000002";
        ram_buffer(46891) := X"00000000";
        ram_buffer(46892) := X"00000000";
        ram_buffer(46893) := X"8FC20078";
        ram_buffer(46894) := X"00000000";
        ram_buffer(46895) := X"24430001";
        ram_buffer(46896) := X"AFC30078";
        ram_buffer(46897) := X"24030039";
        ram_buffer(46898) := X"A0430000";
        ram_buffer(46899) := X"10000089";
        ram_buffer(46900) := X"00000000";
        ram_buffer(46901) := X"8FC20078";
        ram_buffer(46902) := X"00000000";
        ram_buffer(46903) := X"24430001";
        ram_buffer(46904) := X"AFC30078";
        ram_buffer(46905) := X"8FC30020";
        ram_buffer(46906) := X"00000000";
        ram_buffer(46907) := X"306300FF";
        ram_buffer(46908) := X"24630001";
        ram_buffer(46909) := X"306300FF";
        ram_buffer(46910) := X"00031E00";
        ram_buffer(46911) := X"00031E03";
        ram_buffer(46912) := X"A0430000";
        ram_buffer(46913) := X"100000B4";
        ram_buffer(46914) := X"00000000";
        ram_buffer(46915) := X"8FC20078";
        ram_buffer(46916) := X"00000000";
        ram_buffer(46917) := X"24430001";
        ram_buffer(46918) := X"AFC30078";
        ram_buffer(46919) := X"8FC30020";
        ram_buffer(46920) := X"00000000";
        ram_buffer(46921) := X"00031E00";
        ram_buffer(46922) := X"00031E03";
        ram_buffer(46923) := X"A0430000";
        ram_buffer(46924) := X"8FC30024";
        ram_buffer(46925) := X"8FC2002C";
        ram_buffer(46926) := X"00000000";
        ram_buffer(46927) := X"10620051";
        ram_buffer(46928) := X"00000000";
        ram_buffer(46929) := X"00003821";
        ram_buffer(46930) := X"2406000A";
        ram_buffer(46931) := X"8FC50060";
        ram_buffer(46932) := X"8FC400D8";
        ram_buffer(46933) := X"0C02BE38";
        ram_buffer(46934) := X"00000000";
        ram_buffer(46935) := X"AFC20060";
        ram_buffer(46936) := X"8FC30064";
        ram_buffer(46937) := X"8FC20068";
        ram_buffer(46938) := X"00000000";
        ram_buffer(46939) := X"1462000D";
        ram_buffer(46940) := X"00000000";
        ram_buffer(46941) := X"00003821";
        ram_buffer(46942) := X"2406000A";
        ram_buffer(46943) := X"8FC50068";
        ram_buffer(46944) := X"8FC400D8";
        ram_buffer(46945) := X"0C02BE38";
        ram_buffer(46946) := X"00000000";
        ram_buffer(46947) := X"AFC20068";
        ram_buffer(46948) := X"8FC20068";
        ram_buffer(46949) := X"00000000";
        ram_buffer(46950) := X"AFC20064";
        ram_buffer(46951) := X"1000000F";
        ram_buffer(46952) := X"00000000";
        ram_buffer(46953) := X"00003821";
        ram_buffer(46954) := X"2406000A";
        ram_buffer(46955) := X"8FC50064";
        ram_buffer(46956) := X"8FC400D8";
        ram_buffer(46957) := X"0C02BE38";
        ram_buffer(46958) := X"00000000";
        ram_buffer(46959) := X"AFC20064";
        ram_buffer(46960) := X"00003821";
        ram_buffer(46961) := X"2406000A";
        ram_buffer(46962) := X"8FC50068";
        ram_buffer(46963) := X"8FC400D8";
        ram_buffer(46964) := X"0C02BE38";
        ram_buffer(46965) := X"00000000";
        ram_buffer(46966) := X"AFC20068";
        ram_buffer(46967) := X"8FC20024";
        ram_buffer(46968) := X"00000000";
        ram_buffer(46969) := X"24420001";
        ram_buffer(46970) := X"AFC20024";
        ram_buffer(46971) := X"1000FF1D";
        ram_buffer(46972) := X"00000000";
        ram_buffer(46973) := X"24020001";
        ram_buffer(46974) := X"AFC20024";
        ram_buffer(46975) := X"8FD00078";
        ram_buffer(46976) := X"00000000";
        ram_buffer(46977) := X"26020001";
        ram_buffer(46978) := X"AFC20078";
        ram_buffer(46979) := X"8FC5006C";
        ram_buffer(46980) := X"8FC40060";
        ram_buffer(46981) := X"0C02AE52";
        ram_buffer(46982) := X"00000000";
        ram_buffer(46983) := X"24420030";
        ram_buffer(46984) := X"AFC20020";
        ram_buffer(46985) := X"8FC20020";
        ram_buffer(46986) := X"00000000";
        ram_buffer(46987) := X"00021600";
        ram_buffer(46988) := X"00021603";
        ram_buffer(46989) := X"A2020000";
        ram_buffer(46990) := X"8FC30024";
        ram_buffer(46991) := X"8FC2002C";
        ram_buffer(46992) := X"00000000";
        ram_buffer(46993) := X"0062102A";
        ram_buffer(46994) := X"10400011";
        ram_buffer(46995) := X"00000000";
        ram_buffer(46996) := X"00003821";
        ram_buffer(46997) := X"2406000A";
        ram_buffer(46998) := X"8FC50060";
        ram_buffer(46999) := X"8FC400D8";
        ram_buffer(47000) := X"0C02BE38";
        ram_buffer(47001) := X"00000000";
        ram_buffer(47002) := X"AFC20060";
        ram_buffer(47003) := X"8FC20024";
        ram_buffer(47004) := X"00000000";
        ram_buffer(47005) := X"24420001";
        ram_buffer(47006) := X"AFC20024";
        ram_buffer(47007) := X"1000FFDF";
        ram_buffer(47008) := X"00000000";
        ram_buffer(47009) := X"00000000";
        ram_buffer(47010) := X"10000002";
        ram_buffer(47011) := X"00000000";
        ram_buffer(47012) := X"00000000";
        ram_buffer(47013) := X"24060001";
        ram_buffer(47014) := X"8FC50060";
        ram_buffer(47015) := X"8FC400D8";
        ram_buffer(47016) := X"0C02C1BB";
        ram_buffer(47017) := X"00000000";
        ram_buffer(47018) := X"AFC20060";
        ram_buffer(47019) := X"8FC5006C";
        ram_buffer(47020) := X"8FC40060";
        ram_buffer(47021) := X"0C02C26D";
        ram_buffer(47022) := X"00000000";
        ram_buffer(47023) := X"AFC20034";
        ram_buffer(47024) := X"8FC20034";
        ram_buffer(47025) := X"00000000";
        ram_buffer(47026) := X"1C40001D";
        ram_buffer(47027) := X"00000000";
        ram_buffer(47028) := X"8FC20034";
        ram_buffer(47029) := X"00000000";
        ram_buffer(47030) := X"14400031";
        ram_buffer(47031) := X"00000000";
        ram_buffer(47032) := X"8FC20020";
        ram_buffer(47033) := X"00000000";
        ram_buffer(47034) := X"30420001";
        ram_buffer(47035) := X"1040002C";
        ram_buffer(47036) := X"00000000";
        ram_buffer(47037) := X"10000012";
        ram_buffer(47038) := X"00000000";
        ram_buffer(47039) := X"8FC30078";
        ram_buffer(47040) := X"8FC20080";
        ram_buffer(47041) := X"00000000";
        ram_buffer(47042) := X"1462000D";
        ram_buffer(47043) := X"00000000";
        ram_buffer(47044) := X"8FC20038";
        ram_buffer(47045) := X"00000000";
        ram_buffer(47046) := X"24420001";
        ram_buffer(47047) := X"AFC20038";
        ram_buffer(47048) := X"8FC20078";
        ram_buffer(47049) := X"00000000";
        ram_buffer(47050) := X"24430001";
        ram_buffer(47051) := X"AFC30078";
        ram_buffer(47052) := X"24030031";
        ram_buffer(47053) := X"A0430000";
        ram_buffer(47054) := X"10000027";
        ram_buffer(47055) := X"00000000";
        ram_buffer(47056) := X"8FC20078";
        ram_buffer(47057) := X"00000000";
        ram_buffer(47058) := X"2442FFFF";
        ram_buffer(47059) := X"AFC20078";
        ram_buffer(47060) := X"8FC20078";
        ram_buffer(47061) := X"00000000";
        ram_buffer(47062) := X"80430000";
        ram_buffer(47063) := X"24020039";
        ram_buffer(47064) := X"1062FFE6";
        ram_buffer(47065) := X"00000000";
        ram_buffer(47066) := X"8FC20078";
        ram_buffer(47067) := X"00000000";
        ram_buffer(47068) := X"24430001";
        ram_buffer(47069) := X"AFC30078";
        ram_buffer(47070) := X"80430000";
        ram_buffer(47071) := X"00000000";
        ram_buffer(47072) := X"306300FF";
        ram_buffer(47073) := X"24630001";
        ram_buffer(47074) := X"306300FF";
        ram_buffer(47075) := X"00031E00";
        ram_buffer(47076) := X"00031E03";
        ram_buffer(47077) := X"A0430000";
        ram_buffer(47078) := X"1000000F";
        ram_buffer(47079) := X"00000000";
        ram_buffer(47080) := X"8FC20078";
        ram_buffer(47081) := X"00000000";
        ram_buffer(47082) := X"2442FFFF";
        ram_buffer(47083) := X"AFC20078";
        ram_buffer(47084) := X"8FC20078";
        ram_buffer(47085) := X"00000000";
        ram_buffer(47086) := X"80430000";
        ram_buffer(47087) := X"24020030";
        ram_buffer(47088) := X"1062FFF7";
        ram_buffer(47089) := X"00000000";
        ram_buffer(47090) := X"8FC20078";
        ram_buffer(47091) := X"00000000";
        ram_buffer(47092) := X"24420001";
        ram_buffer(47093) := X"AFC20078";
        ram_buffer(47094) := X"8FC5006C";
        ram_buffer(47095) := X"8FC400D8";
        ram_buffer(47096) := X"0C02BE10";
        ram_buffer(47097) := X"00000000";
        ram_buffer(47098) := X"8FC20068";
        ram_buffer(47099) := X"00000000";
        ram_buffer(47100) := X"10400015";
        ram_buffer(47101) := X"00000000";
        ram_buffer(47102) := X"8FC20064";
        ram_buffer(47103) := X"00000000";
        ram_buffer(47104) := X"1040000A";
        ram_buffer(47105) := X"00000000";
        ram_buffer(47106) := X"8FC30064";
        ram_buffer(47107) := X"8FC20068";
        ram_buffer(47108) := X"00000000";
        ram_buffer(47109) := X"10620005";
        ram_buffer(47110) := X"00000000";
        ram_buffer(47111) := X"8FC50064";
        ram_buffer(47112) := X"8FC400D8";
        ram_buffer(47113) := X"0C02BE10";
        ram_buffer(47114) := X"00000000";
        ram_buffer(47115) := X"8FC50068";
        ram_buffer(47116) := X"8FC400D8";
        ram_buffer(47117) := X"0C02BE10";
        ram_buffer(47118) := X"00000000";
        ram_buffer(47119) := X"10000002";
        ram_buffer(47120) := X"00000000";
        ram_buffer(47121) := X"00000000";
        ram_buffer(47122) := X"8FC50060";
        ram_buffer(47123) := X"8FC400D8";
        ram_buffer(47124) := X"0C02BE10";
        ram_buffer(47125) := X"00000000";
        ram_buffer(47126) := X"8FC20078";
        ram_buffer(47127) := X"00000000";
        ram_buffer(47128) := X"A0400000";
        ram_buffer(47129) := X"8FC20038";
        ram_buffer(47130) := X"00000000";
        ram_buffer(47131) := X"24430001";
        ram_buffer(47132) := X"8FC200F0";
        ram_buffer(47133) := X"00000000";
        ram_buffer(47134) := X"AC430000";
        ram_buffer(47135) := X"8FC200F8";
        ram_buffer(47136) := X"00000000";
        ram_buffer(47137) := X"10400005";
        ram_buffer(47138) := X"00000000";
        ram_buffer(47139) := X"8FC200F8";
        ram_buffer(47140) := X"8FC30078";
        ram_buffer(47141) := X"00000000";
        ram_buffer(47142) := X"AC430000";
        ram_buffer(47143) := X"8FC20080";
        ram_buffer(47144) := X"03C0E821";
        ram_buffer(47145) := X"8FBF00D4";
        ram_buffer(47146) := X"8FBE00D0";
        ram_buffer(47147) := X"8FB300CC";
        ram_buffer(47148) := X"8FB200C8";
        ram_buffer(47149) := X"8FB100C4";
        ram_buffer(47150) := X"8FB000C0";
        ram_buffer(47151) := X"27BD00D8";
        ram_buffer(47152) := X"03E00008";
        ram_buffer(47153) := X"00000000";
        ram_buffer(47154) := X"27BDFFF8";
        ram_buffer(47155) := X"AFBE0004";
        ram_buffer(47156) := X"03A0F021";
        ram_buffer(47157) := X"AFC40008";
        ram_buffer(47158) := X"00000000";
        ram_buffer(47159) := X"03C0E821";
        ram_buffer(47160) := X"8FBE0004";
        ram_buffer(47161) := X"27BD0008";
        ram_buffer(47162) := X"03E00008";
        ram_buffer(47163) := X"00000000";
        ram_buffer(47164) := X"27BDFFF8";
        ram_buffer(47165) := X"AFBE0004";
        ram_buffer(47166) := X"03A0F021";
        ram_buffer(47167) := X"AFC40008";
        ram_buffer(47168) := X"00000000";
        ram_buffer(47169) := X"03C0E821";
        ram_buffer(47170) := X"8FBE0004";
        ram_buffer(47171) := X"27BD0008";
        ram_buffer(47172) := X"03E00008";
        ram_buffer(47173) := X"00000000";
        ram_buffer(47174) := X"27BDFFF0";
        ram_buffer(47175) := X"AFBE000C";
        ram_buffer(47176) := X"AFB20008";
        ram_buffer(47177) := X"AFB10004";
        ram_buffer(47178) := X"AFB00000";
        ram_buffer(47179) := X"03A0F021";
        ram_buffer(47180) := X"AFC40010";
        ram_buffer(47181) := X"00A01021";
        ram_buffer(47182) := X"AFC60018";
        ram_buffer(47183) := X"80430000";
        ram_buffer(47184) := X"24040072";
        ram_buffer(47185) := X"10640009";
        ram_buffer(47186) := X"00000000";
        ram_buffer(47187) := X"24040077";
        ram_buffer(47188) := X"1064000B";
        ram_buffer(47189) := X"00000000";
        ram_buffer(47190) := X"24040061";
        ram_buffer(47191) := X"1064000D";
        ram_buffer(47192) := X"00000000";
        ram_buffer(47193) := X"10000010";
        ram_buffer(47194) := X"00000000";
        ram_buffer(47195) := X"24110004";
        ram_buffer(47196) := X"00008021";
        ram_buffer(47197) := X"00009021";
        ram_buffer(47198) := X"10000011";
        ram_buffer(47199) := X"00000000";
        ram_buffer(47200) := X"24110008";
        ram_buffer(47201) := X"24100001";
        ram_buffer(47202) := X"24120600";
        ram_buffer(47203) := X"1000000C";
        ram_buffer(47204) := X"00000000";
        ram_buffer(47205) := X"24110108";
        ram_buffer(47206) := X"24100001";
        ram_buffer(47207) := X"24120208";
        ram_buffer(47208) := X"10000007";
        ram_buffer(47209) := X"00000000";
        ram_buffer(47210) := X"8FC20010";
        ram_buffer(47211) := X"24030016";
        ram_buffer(47212) := X"AC430000";
        ram_buffer(47213) := X"00001021";
        ram_buffer(47214) := X"10000023";
        ram_buffer(47215) := X"00000000";
        ram_buffer(47216) := X"10000017";
        ram_buffer(47217) := X"00000000";
        ram_buffer(47218) := X"80430000";
        ram_buffer(47219) := X"24040062";
        ram_buffer(47220) := X"10640013";
        ram_buffer(47221) := X"00000000";
        ram_buffer(47222) := X"24040078";
        ram_buffer(47223) := X"1064000C";
        ram_buffer(47224) := X"00000000";
        ram_buffer(47225) := X"2404002B";
        ram_buffer(47226) := X"1464000C";
        ram_buffer(47227) := X"00000000";
        ram_buffer(47228) := X"2403FFE3";
        ram_buffer(47229) := X"02231824";
        ram_buffer(47230) := X"34710010";
        ram_buffer(47231) := X"2403FFFC";
        ram_buffer(47232) := X"02031824";
        ram_buffer(47233) := X"34700002";
        ram_buffer(47234) := X"10000005";
        ram_buffer(47235) := X"00000000";
        ram_buffer(47236) := X"36100800";
        ram_buffer(47237) := X"10000002";
        ram_buffer(47238) := X"00000000";
        ram_buffer(47239) := X"00000000";
        ram_buffer(47240) := X"24420001";
        ram_buffer(47241) := X"80430000";
        ram_buffer(47242) := X"00000000";
        ram_buffer(47243) := X"1460FFE6";
        ram_buffer(47244) := X"00000000";
        ram_buffer(47245) := X"02121825";
        ram_buffer(47246) := X"8FC20018";
        ram_buffer(47247) := X"00000000";
        ram_buffer(47248) := X"AC430000";
        ram_buffer(47249) := X"02201021";
        ram_buffer(47250) := X"03C0E821";
        ram_buffer(47251) := X"8FBE000C";
        ram_buffer(47252) := X"8FB20008";
        ram_buffer(47253) := X"8FB10004";
        ram_buffer(47254) := X"8FB00000";
        ram_buffer(47255) := X"27BD0010";
        ram_buffer(47256) := X"03E00008";
        ram_buffer(47257) := X"00000000";
        ram_buffer(47258) := X"27BDFFB8";
        ram_buffer(47259) := X"AFBF0044";
        ram_buffer(47260) := X"AFBE0040";
        ram_buffer(47261) := X"AFB5003C";
        ram_buffer(47262) := X"AFB40038";
        ram_buffer(47263) := X"AFB30034";
        ram_buffer(47264) := X"AFB20030";
        ram_buffer(47265) := X"AFB1002C";
        ram_buffer(47266) := X"AFB00028";
        ram_buffer(47267) := X"03A0F021";
        ram_buffer(47268) := X"AFC40048";
        ram_buffer(47269) := X"00A08021";
        ram_buffer(47270) := X"00C0A821";
        ram_buffer(47271) := X"00009821";
        ram_buffer(47272) := X"8EB20008";
        ram_buffer(47273) := X"00000000";
        ram_buffer(47274) := X"16400004";
        ram_buffer(47275) := X"00000000";
        ram_buffer(47276) := X"00001021";
        ram_buffer(47277) := X"100001E2";
        ram_buffer(47278) := X"00000000";
        ram_buffer(47279) := X"8602000C";
        ram_buffer(47280) := X"00000000";
        ram_buffer(47281) := X"3042FFFF";
        ram_buffer(47282) := X"30420008";
        ram_buffer(47283) := X"10400005";
        ram_buffer(47284) := X"00000000";
        ram_buffer(47285) := X"8E020010";
        ram_buffer(47286) := X"00000000";
        ram_buffer(47287) := X"1440000A";
        ram_buffer(47288) := X"00000000";
        ram_buffer(47289) := X"02002821";
        ram_buffer(47290) := X"8FC40048";
        ram_buffer(47291) := X"0C02ACF1";
        ram_buffer(47292) := X"00000000";
        ram_buffer(47293) := X"10400004";
        ram_buffer(47294) := X"00000000";
        ram_buffer(47295) := X"2402FFFF";
        ram_buffer(47296) := X"100001CF";
        ram_buffer(47297) := X"00000000";
        ram_buffer(47298) := X"8EB40000";
        ram_buffer(47299) := X"00009021";
        ram_buffer(47300) := X"8602000C";
        ram_buffer(47301) := X"00000000";
        ram_buffer(47302) := X"3042FFFF";
        ram_buffer(47303) := X"30420002";
        ram_buffer(47304) := X"10400028";
        ram_buffer(47305) := X"00000000";
        ram_buffer(47306) := X"10000004";
        ram_buffer(47307) := X"00000000";
        ram_buffer(47308) := X"8E930000";
        ram_buffer(47309) := X"8E920004";
        ram_buffer(47310) := X"26940008";
        ram_buffer(47311) := X"1240FFFC";
        ram_buffer(47312) := X"00000000";
        ram_buffer(47313) := X"8E030024";
        ram_buffer(47314) := X"8E05001C";
        ram_buffer(47315) := X"02401021";
        ram_buffer(47316) := X"3C047FFF";
        ram_buffer(47317) := X"3484FC01";
        ram_buffer(47318) := X"0044202B";
        ram_buffer(47319) := X"14800003";
        ram_buffer(47320) := X"00000000";
        ram_buffer(47321) := X"3C027FFF";
        ram_buffer(47322) := X"3442FC00";
        ram_buffer(47323) := X"00403821";
        ram_buffer(47324) := X"02603021";
        ram_buffer(47325) := X"8FC40048";
        ram_buffer(47326) := X"0060F809";
        ram_buffer(47327) := X"00000000";
        ram_buffer(47328) := X"00408821";
        ram_buffer(47329) := X"1A2001A0";
        ram_buffer(47330) := X"00000000";
        ram_buffer(47331) := X"02201021";
        ram_buffer(47332) := X"02629821";
        ram_buffer(47333) := X"02201021";
        ram_buffer(47334) := X"02429023";
        ram_buffer(47335) := X"8EA20008";
        ram_buffer(47336) := X"02201821";
        ram_buffer(47337) := X"00431023";
        ram_buffer(47338) := X"AEA20008";
        ram_buffer(47339) := X"8EA20008";
        ram_buffer(47340) := X"00000000";
        ram_buffer(47341) := X"1440FFE1";
        ram_buffer(47342) := X"00000000";
        ram_buffer(47343) := X"1000018F";
        ram_buffer(47344) := X"00000000";
        ram_buffer(47345) := X"8602000C";
        ram_buffer(47346) := X"00000000";
        ram_buffer(47347) := X"3042FFFF";
        ram_buffer(47348) := X"30420001";
        ram_buffer(47349) := X"14400101";
        ram_buffer(47350) := X"00000000";
        ram_buffer(47351) := X"10000004";
        ram_buffer(47352) := X"00000000";
        ram_buffer(47353) := X"8E930000";
        ram_buffer(47354) := X"8E920004";
        ram_buffer(47355) := X"26940008";
        ram_buffer(47356) := X"1240FFFC";
        ram_buffer(47357) := X"00000000";
        ram_buffer(47358) := X"8E110008";
        ram_buffer(47359) := X"8602000C";
        ram_buffer(47360) := X"00000000";
        ram_buffer(47361) := X"3042FFFF";
        ram_buffer(47362) := X"30420200";
        ram_buffer(47363) := X"10400098";
        ram_buffer(47364) := X"00000000";
        ram_buffer(47365) := X"02201021";
        ram_buffer(47366) := X"0242102B";
        ram_buffer(47367) := X"1440007D";
        ram_buffer(47368) := X"00000000";
        ram_buffer(47369) := X"8602000C";
        ram_buffer(47370) := X"00000000";
        ram_buffer(47371) := X"3042FFFF";
        ram_buffer(47372) := X"30420480";
        ram_buffer(47373) := X"10400077";
        ram_buffer(47374) := X"00000000";
        ram_buffer(47375) := X"8E020000";
        ram_buffer(47376) := X"00000000";
        ram_buffer(47377) := X"00401821";
        ram_buffer(47378) := X"8E020010";
        ram_buffer(47379) := X"00000000";
        ram_buffer(47380) := X"00621023";
        ram_buffer(47381) := X"AFC20020";
        ram_buffer(47382) := X"8E030014";
        ram_buffer(47383) := X"00000000";
        ram_buffer(47384) := X"00601021";
        ram_buffer(47385) := X"00021040";
        ram_buffer(47386) := X"00431021";
        ram_buffer(47387) := X"00021FC2";
        ram_buffer(47388) := X"00621021";
        ram_buffer(47389) := X"00021043";
        ram_buffer(47390) := X"AFC2001C";
        ram_buffer(47391) := X"8FC20020";
        ram_buffer(47392) := X"00000000";
        ram_buffer(47393) := X"00521021";
        ram_buffer(47394) := X"24430001";
        ram_buffer(47395) := X"8FC2001C";
        ram_buffer(47396) := X"00000000";
        ram_buffer(47397) := X"0043102B";
        ram_buffer(47398) := X"10400006";
        ram_buffer(47399) := X"00000000";
        ram_buffer(47400) := X"8FC20020";
        ram_buffer(47401) := X"00000000";
        ram_buffer(47402) := X"00521021";
        ram_buffer(47403) := X"24420001";
        ram_buffer(47404) := X"AFC2001C";
        ram_buffer(47405) := X"8602000C";
        ram_buffer(47406) := X"00000000";
        ram_buffer(47407) := X"3042FFFF";
        ram_buffer(47408) := X"30420400";
        ram_buffer(47409) := X"10400024";
        ram_buffer(47410) := X"00000000";
        ram_buffer(47411) := X"8FC2001C";
        ram_buffer(47412) := X"00000000";
        ram_buffer(47413) := X"00402821";
        ram_buffer(47414) := X"8FC40048";
        ram_buffer(47415) := X"0C027B8F";
        ram_buffer(47416) := X"00000000";
        ram_buffer(47417) := X"AFC20018";
        ram_buffer(47418) := X"8FC20018";
        ram_buffer(47419) := X"00000000";
        ram_buffer(47420) := X"14400006";
        ram_buffer(47421) := X"00000000";
        ram_buffer(47422) := X"8FC20048";
        ram_buffer(47423) := X"2403000C";
        ram_buffer(47424) := X"AC430000";
        ram_buffer(47425) := X"10000147";
        ram_buffer(47426) := X"00000000";
        ram_buffer(47427) := X"8E020010";
        ram_buffer(47428) := X"8FC30020";
        ram_buffer(47429) := X"00000000";
        ram_buffer(47430) := X"00603021";
        ram_buffer(47431) := X"00402821";
        ram_buffer(47432) := X"8FC40018";
        ram_buffer(47433) := X"0C027F93";
        ram_buffer(47434) := X"00000000";
        ram_buffer(47435) := X"8603000C";
        ram_buffer(47436) := X"2402FB7F";
        ram_buffer(47437) := X"00621024";
        ram_buffer(47438) := X"00021400";
        ram_buffer(47439) := X"00021403";
        ram_buffer(47440) := X"34420080";
        ram_buffer(47441) := X"00021400";
        ram_buffer(47442) := X"00021403";
        ram_buffer(47443) := X"A602000C";
        ram_buffer(47444) := X"1000001F";
        ram_buffer(47445) := X"00000000";
        ram_buffer(47446) := X"8E020010";
        ram_buffer(47447) := X"8FC3001C";
        ram_buffer(47448) := X"00000000";
        ram_buffer(47449) := X"00603021";
        ram_buffer(47450) := X"00402821";
        ram_buffer(47451) := X"8FC40048";
        ram_buffer(47452) := X"0C02C6A7";
        ram_buffer(47453) := X"00000000";
        ram_buffer(47454) := X"AFC20018";
        ram_buffer(47455) := X"8FC20018";
        ram_buffer(47456) := X"00000000";
        ram_buffer(47457) := X"14400012";
        ram_buffer(47458) := X"00000000";
        ram_buffer(47459) := X"8E020010";
        ram_buffer(47460) := X"00000000";
        ram_buffer(47461) := X"00402821";
        ram_buffer(47462) := X"8FC40048";
        ram_buffer(47463) := X"0C027301";
        ram_buffer(47464) := X"00000000";
        ram_buffer(47465) := X"8603000C";
        ram_buffer(47466) := X"2402FF7F";
        ram_buffer(47467) := X"00621024";
        ram_buffer(47468) := X"00021400";
        ram_buffer(47469) := X"00021403";
        ram_buffer(47470) := X"A602000C";
        ram_buffer(47471) := X"8FC20048";
        ram_buffer(47472) := X"2403000C";
        ram_buffer(47473) := X"AC430000";
        ram_buffer(47474) := X"10000116";
        ram_buffer(47475) := X"00000000";
        ram_buffer(47476) := X"8FC20018";
        ram_buffer(47477) := X"00000000";
        ram_buffer(47478) := X"AE020010";
        ram_buffer(47479) := X"8FC20020";
        ram_buffer(47480) := X"8FC30018";
        ram_buffer(47481) := X"00000000";
        ram_buffer(47482) := X"00621021";
        ram_buffer(47483) := X"AE020000";
        ram_buffer(47484) := X"8FC2001C";
        ram_buffer(47485) := X"00000000";
        ram_buffer(47486) := X"AE020014";
        ram_buffer(47487) := X"02408821";
        ram_buffer(47488) := X"8FC3001C";
        ram_buffer(47489) := X"8FC20020";
        ram_buffer(47490) := X"00000000";
        ram_buffer(47491) := X"00621023";
        ram_buffer(47492) := X"AE020008";
        ram_buffer(47493) := X"02201021";
        ram_buffer(47494) := X"0242102B";
        ram_buffer(47495) := X"10400002";
        ram_buffer(47496) := X"00000000";
        ram_buffer(47497) := X"02408821";
        ram_buffer(47498) := X"8E020000";
        ram_buffer(47499) := X"02201821";
        ram_buffer(47500) := X"00603021";
        ram_buffer(47501) := X"02602821";
        ram_buffer(47502) := X"00402021";
        ram_buffer(47503) := X"0C02BCED";
        ram_buffer(47504) := X"00000000";
        ram_buffer(47505) := X"8E020008";
        ram_buffer(47506) := X"00000000";
        ram_buffer(47507) := X"00511023";
        ram_buffer(47508) := X"AE020008";
        ram_buffer(47509) := X"8E020000";
        ram_buffer(47510) := X"02201821";
        ram_buffer(47511) := X"00431021";
        ram_buffer(47512) := X"AE020000";
        ram_buffer(47513) := X"02408821";
        ram_buffer(47514) := X"1000004E";
        ram_buffer(47515) := X"00000000";
        ram_buffer(47516) := X"8E030000";
        ram_buffer(47517) := X"8E020010";
        ram_buffer(47518) := X"00000000";
        ram_buffer(47519) := X"0043102B";
        ram_buffer(47520) := X"14400006";
        ram_buffer(47521) := X"00000000";
        ram_buffer(47522) := X"8E020014";
        ram_buffer(47523) := X"00000000";
        ram_buffer(47524) := X"0242102B";
        ram_buffer(47525) := X"10400022";
        ram_buffer(47526) := X"00000000";
        ram_buffer(47527) := X"02201021";
        ram_buffer(47528) := X"0242182B";
        ram_buffer(47529) := X"10600002";
        ram_buffer(47530) := X"00000000";
        ram_buffer(47531) := X"02401021";
        ram_buffer(47532) := X"00408821";
        ram_buffer(47533) := X"8E020000";
        ram_buffer(47534) := X"02201821";
        ram_buffer(47535) := X"00603021";
        ram_buffer(47536) := X"02602821";
        ram_buffer(47537) := X"00402021";
        ram_buffer(47538) := X"0C02BCED";
        ram_buffer(47539) := X"00000000";
        ram_buffer(47540) := X"8E020008";
        ram_buffer(47541) := X"00000000";
        ram_buffer(47542) := X"00511023";
        ram_buffer(47543) := X"AE020008";
        ram_buffer(47544) := X"8E020000";
        ram_buffer(47545) := X"02201821";
        ram_buffer(47546) := X"00431021";
        ram_buffer(47547) := X"AE020000";
        ram_buffer(47548) := X"8E020008";
        ram_buffer(47549) := X"00000000";
        ram_buffer(47550) := X"14400029";
        ram_buffer(47551) := X"00000000";
        ram_buffer(47552) := X"02002821";
        ram_buffer(47553) := X"8FC40048";
        ram_buffer(47554) := X"0C026EE1";
        ram_buffer(47555) := X"00000000";
        ram_buffer(47556) := X"10400023";
        ram_buffer(47557) := X"00000000";
        ram_buffer(47558) := X"100000C2";
        ram_buffer(47559) := X"00000000";
        ram_buffer(47560) := X"02401021";
        ram_buffer(47561) := X"3C038000";
        ram_buffer(47562) := X"0043182B";
        ram_buffer(47563) := X"14600003";
        ram_buffer(47564) := X"00000000";
        ram_buffer(47565) := X"3C027FFF";
        ram_buffer(47566) := X"3442FFFF";
        ram_buffer(47567) := X"00401821";
        ram_buffer(47568) := X"8E020014";
        ram_buffer(47569) := X"00000000";
        ram_buffer(47570) := X"14400002";
        ram_buffer(47571) := X"0062001A";
        ram_buffer(47572) := X"0007000D";
        ram_buffer(47573) := X"00001010";
        ram_buffer(47574) := X"00001812";
        ram_buffer(47575) := X"8E020014";
        ram_buffer(47576) := X"00000000";
        ram_buffer(47577) := X"00620018";
        ram_buffer(47578) := X"00008812";
        ram_buffer(47579) := X"8E020024";
        ram_buffer(47580) := X"8E03001C";
        ram_buffer(47581) := X"02203821";
        ram_buffer(47582) := X"02603021";
        ram_buffer(47583) := X"00602821";
        ram_buffer(47584) := X"8FC40048";
        ram_buffer(47585) := X"0040F809";
        ram_buffer(47586) := X"00000000";
        ram_buffer(47587) := X"00408821";
        ram_buffer(47588) := X"1A2000A0";
        ram_buffer(47589) := X"00000000";
        ram_buffer(47590) := X"10000002";
        ram_buffer(47591) := X"00000000";
        ram_buffer(47592) := X"00000000";
        ram_buffer(47593) := X"02201021";
        ram_buffer(47594) := X"02629821";
        ram_buffer(47595) := X"02201021";
        ram_buffer(47596) := X"02429023";
        ram_buffer(47597) := X"8EA20008";
        ram_buffer(47598) := X"02201821";
        ram_buffer(47599) := X"00431023";
        ram_buffer(47600) := X"AEA20008";
        ram_buffer(47601) := X"8EA20008";
        ram_buffer(47602) := X"00000000";
        ram_buffer(47603) := X"1440FF08";
        ram_buffer(47604) := X"00000000";
        ram_buffer(47605) := X"10000089";
        ram_buffer(47606) := X"00000000";
        ram_buffer(47607) := X"AFC00010";
        ram_buffer(47608) := X"AFC00014";
        ram_buffer(47609) := X"10000005";
        ram_buffer(47610) := X"00000000";
        ram_buffer(47611) := X"AFC00010";
        ram_buffer(47612) := X"8E930000";
        ram_buffer(47613) := X"8E920004";
        ram_buffer(47614) := X"26940008";
        ram_buffer(47615) := X"1240FFFB";
        ram_buffer(47616) := X"00000000";
        ram_buffer(47617) := X"8FC20010";
        ram_buffer(47618) := X"00000000";
        ram_buffer(47619) := X"14400017";
        ram_buffer(47620) := X"00000000";
        ram_buffer(47621) := X"02403021";
        ram_buffer(47622) := X"2405000A";
        ram_buffer(47623) := X"02602021";
        ram_buffer(47624) := X"0C02BC51";
        ram_buffer(47625) := X"00000000";
        ram_buffer(47626) := X"AFC20024";
        ram_buffer(47627) := X"8FC20024";
        ram_buffer(47628) := X"00000000";
        ram_buffer(47629) := X"10400009";
        ram_buffer(47630) := X"00000000";
        ram_buffer(47631) := X"8FC20024";
        ram_buffer(47632) := X"00000000";
        ram_buffer(47633) := X"24420001";
        ram_buffer(47634) := X"00401821";
        ram_buffer(47635) := X"02601021";
        ram_buffer(47636) := X"00621023";
        ram_buffer(47637) := X"10000002";
        ram_buffer(47638) := X"00000000";
        ram_buffer(47639) := X"26420001";
        ram_buffer(47640) := X"AFC20014";
        ram_buffer(47641) := X"24020001";
        ram_buffer(47642) := X"AFC20010";
        ram_buffer(47643) := X"8FC20014";
        ram_buffer(47644) := X"00000000";
        ram_buffer(47645) := X"0242182B";
        ram_buffer(47646) := X"10600002";
        ram_buffer(47647) := X"00000000";
        ram_buffer(47648) := X"02401021";
        ram_buffer(47649) := X"0040F821";
        ram_buffer(47650) := X"8E030008";
        ram_buffer(47651) := X"8E020014";
        ram_buffer(47652) := X"00000000";
        ram_buffer(47653) := X"00628821";
        ram_buffer(47654) := X"8E030000";
        ram_buffer(47655) := X"8E020010";
        ram_buffer(47656) := X"00000000";
        ram_buffer(47657) := X"0043102B";
        ram_buffer(47658) := X"10400017";
        ram_buffer(47659) := X"00000000";
        ram_buffer(47660) := X"023F102A";
        ram_buffer(47661) := X"10400014";
        ram_buffer(47662) := X"00000000";
        ram_buffer(47663) := X"8E020000";
        ram_buffer(47664) := X"02201821";
        ram_buffer(47665) := X"00603021";
        ram_buffer(47666) := X"02602821";
        ram_buffer(47667) := X"00402021";
        ram_buffer(47668) := X"0C02BCED";
        ram_buffer(47669) := X"00000000";
        ram_buffer(47670) := X"8E020000";
        ram_buffer(47671) := X"02201821";
        ram_buffer(47672) := X"00431021";
        ram_buffer(47673) := X"AE020000";
        ram_buffer(47674) := X"02002821";
        ram_buffer(47675) := X"8FC40048";
        ram_buffer(47676) := X"0C026EE1";
        ram_buffer(47677) := X"00000000";
        ram_buffer(47678) := X"10400025";
        ram_buffer(47679) := X"00000000";
        ram_buffer(47680) := X"10000048";
        ram_buffer(47681) := X"00000000";
        ram_buffer(47682) := X"8E110014";
        ram_buffer(47683) := X"00000000";
        ram_buffer(47684) := X"03F1102A";
        ram_buffer(47685) := X"1440000E";
        ram_buffer(47686) := X"00000000";
        ram_buffer(47687) := X"8E020024";
        ram_buffer(47688) := X"8E03001C";
        ram_buffer(47689) := X"02203821";
        ram_buffer(47690) := X"02603021";
        ram_buffer(47691) := X"00602821";
        ram_buffer(47692) := X"8FC40048";
        ram_buffer(47693) := X"0040F809";
        ram_buffer(47694) := X"00000000";
        ram_buffer(47695) := X"00408821";
        ram_buffer(47696) := X"1E200013";
        ram_buffer(47697) := X"00000000";
        ram_buffer(47698) := X"10000036";
        ram_buffer(47699) := X"00000000";
        ram_buffer(47700) := X"03E08821";
        ram_buffer(47701) := X"8E020000";
        ram_buffer(47702) := X"02201821";
        ram_buffer(47703) := X"00603021";
        ram_buffer(47704) := X"02602821";
        ram_buffer(47705) := X"00402021";
        ram_buffer(47706) := X"0C02BCED";
        ram_buffer(47707) := X"00000000";
        ram_buffer(47708) := X"8E020008";
        ram_buffer(47709) := X"00000000";
        ram_buffer(47710) := X"00511023";
        ram_buffer(47711) := X"AE020008";
        ram_buffer(47712) := X"8E020000";
        ram_buffer(47713) := X"02201821";
        ram_buffer(47714) := X"00431021";
        ram_buffer(47715) := X"AE020000";
        ram_buffer(47716) := X"8FC20014";
        ram_buffer(47717) := X"00000000";
        ram_buffer(47718) := X"00511023";
        ram_buffer(47719) := X"AFC20014";
        ram_buffer(47720) := X"8FC20014";
        ram_buffer(47721) := X"00000000";
        ram_buffer(47722) := X"14400008";
        ram_buffer(47723) := X"00000000";
        ram_buffer(47724) := X"02002821";
        ram_buffer(47725) := X"8FC40048";
        ram_buffer(47726) := X"0C026EE1";
        ram_buffer(47727) := X"00000000";
        ram_buffer(47728) := X"14400017";
        ram_buffer(47729) := X"00000000";
        ram_buffer(47730) := X"AFC00010";
        ram_buffer(47731) := X"02201021";
        ram_buffer(47732) := X"02629821";
        ram_buffer(47733) := X"02201021";
        ram_buffer(47734) := X"02429023";
        ram_buffer(47735) := X"8EA20008";
        ram_buffer(47736) := X"02201821";
        ram_buffer(47737) := X"00431023";
        ram_buffer(47738) := X"AEA20008";
        ram_buffer(47739) := X"8EA20008";
        ram_buffer(47740) := X"00000000";
        ram_buffer(47741) := X"1440FF81";
        ram_buffer(47742) := X"00000000";
        ram_buffer(47743) := X"00001021";
        ram_buffer(47744) := X"1000000F";
        ram_buffer(47745) := X"00000000";
        ram_buffer(47746) := X"00000000";
        ram_buffer(47747) := X"10000005";
        ram_buffer(47748) := X"00000000";
        ram_buffer(47749) := X"00000000";
        ram_buffer(47750) := X"10000002";
        ram_buffer(47751) := X"00000000";
        ram_buffer(47752) := X"00000000";
        ram_buffer(47753) := X"8602000C";
        ram_buffer(47754) := X"00000000";
        ram_buffer(47755) := X"34420040";
        ram_buffer(47756) := X"00021400";
        ram_buffer(47757) := X"00021403";
        ram_buffer(47758) := X"A602000C";
        ram_buffer(47759) := X"2402FFFF";
        ram_buffer(47760) := X"03C0E821";
        ram_buffer(47761) := X"8FBF0044";
        ram_buffer(47762) := X"8FBE0040";
        ram_buffer(47763) := X"8FB5003C";
        ram_buffer(47764) := X"8FB40038";
        ram_buffer(47765) := X"8FB30034";
        ram_buffer(47766) := X"8FB20030";
        ram_buffer(47767) := X"8FB1002C";
        ram_buffer(47768) := X"8FB00028";
        ram_buffer(47769) := X"27BD0048";
        ram_buffer(47770) := X"03E00008";
        ram_buffer(47771) := X"00000000";
        ram_buffer(47772) := X"27BDFFE0";
        ram_buffer(47773) := X"AFBF001C";
        ram_buffer(47774) := X"AFBE0018";
        ram_buffer(47775) := X"03A0F021";
        ram_buffer(47776) := X"AFC40020";
        ram_buffer(47777) := X"AFC50024";
        ram_buffer(47778) := X"AF8081EC";
        ram_buffer(47779) := X"8FC40024";
        ram_buffer(47780) := X"0C02FBBB";
        ram_buffer(47781) := X"00000000";
        ram_buffer(47782) := X"AFC20010";
        ram_buffer(47783) := X"8FC30010";
        ram_buffer(47784) := X"2402FFFF";
        ram_buffer(47785) := X"14620009";
        ram_buffer(47786) := X"00000000";
        ram_buffer(47787) := X"8F8281EC";
        ram_buffer(47788) := X"00000000";
        ram_buffer(47789) := X"10400005";
        ram_buffer(47790) := X"00000000";
        ram_buffer(47791) := X"8F8381EC";
        ram_buffer(47792) := X"8FC20020";
        ram_buffer(47793) := X"00000000";
        ram_buffer(47794) := X"AC430000";
        ram_buffer(47795) := X"8FC20010";
        ram_buffer(47796) := X"03C0E821";
        ram_buffer(47797) := X"8FBF001C";
        ram_buffer(47798) := X"8FBE0018";
        ram_buffer(47799) := X"27BD0020";
        ram_buffer(47800) := X"03E00008";
        ram_buffer(47801) := X"00000000";
        ram_buffer(47802) := X"27BDFFF8";
        ram_buffer(47803) := X"AFBE0004";
        ram_buffer(47804) := X"03A0F021";
        ram_buffer(47805) := X"AFC40008";
        ram_buffer(47806) := X"8FC20008";
        ram_buffer(47807) := X"00000000";
        ram_buffer(47808) := X"2C420100";
        ram_buffer(47809) := X"1040000C";
        ram_buffer(47810) := X"00000000";
        ram_buffer(47811) := X"8F838090";
        ram_buffer(47812) := X"8FC20008";
        ram_buffer(47813) := X"00000000";
        ram_buffer(47814) := X"24420001";
        ram_buffer(47815) := X"00621021";
        ram_buffer(47816) := X"80420000";
        ram_buffer(47817) := X"00000000";
        ram_buffer(47818) := X"304200FF";
        ram_buffer(47819) := X"30420008";
        ram_buffer(47820) := X"10000002";
        ram_buffer(47821) := X"00000000";
        ram_buffer(47822) := X"00001021";
        ram_buffer(47823) := X"03C0E821";
        ram_buffer(47824) := X"8FBE0004";
        ram_buffer(47825) := X"27BD0008";
        ram_buffer(47826) := X"03E00008";
        ram_buffer(47827) := X"00000000";
        ram_buffer(47828) := X"27BDFFE8";
        ram_buffer(47829) := X"AFBF0014";
        ram_buffer(47830) := X"AFBE0010";
        ram_buffer(47831) := X"03A0F021";
        ram_buffer(47832) := X"AFC40018";
        ram_buffer(47833) := X"AFC5001C";
        ram_buffer(47834) := X"AFC60020";
        ram_buffer(47835) := X"8FC20020";
        ram_buffer(47836) := X"00000000";
        ram_buffer(47837) := X"10400019";
        ram_buffer(47838) := X"00000000";
        ram_buffer(47839) := X"3C02100D";
        ram_buffer(47840) := X"2445A924";
        ram_buffer(47841) := X"8FC40020";
        ram_buffer(47842) := X"0C02CC2F";
        ram_buffer(47843) := X"00000000";
        ram_buffer(47844) := X"10400012";
        ram_buffer(47845) := X"00000000";
        ram_buffer(47846) := X"3C02100D";
        ram_buffer(47847) := X"2445A92C";
        ram_buffer(47848) := X"8FC40020";
        ram_buffer(47849) := X"0C02CC2F";
        ram_buffer(47850) := X"00000000";
        ram_buffer(47851) := X"1040000B";
        ram_buffer(47852) := X"00000000";
        ram_buffer(47853) := X"3C02100D";
        ram_buffer(47854) := X"2445A920";
        ram_buffer(47855) := X"8FC40020";
        ram_buffer(47856) := X"0C02CC2F";
        ram_buffer(47857) := X"00000000";
        ram_buffer(47858) := X"10400004";
        ram_buffer(47859) := X"00000000";
        ram_buffer(47860) := X"00001021";
        ram_buffer(47861) := X"10000003";
        ram_buffer(47862) := X"00000000";
        ram_buffer(47863) := X"3C02100D";
        ram_buffer(47864) := X"2442A92C";
        ram_buffer(47865) := X"03C0E821";
        ram_buffer(47866) := X"8FBF0014";
        ram_buffer(47867) := X"8FBE0010";
        ram_buffer(47868) := X"27BD0018";
        ram_buffer(47869) := X"03E00008";
        ram_buffer(47870) := X"00000000";
        ram_buffer(47871) := X"27BDFFF8";
        ram_buffer(47872) := X"AFBE0004";
        ram_buffer(47873) := X"03A0F021";
        ram_buffer(47874) := X"3C02100D";
        ram_buffer(47875) := X"2442D020";
        ram_buffer(47876) := X"03C0E821";
        ram_buffer(47877) := X"8FBE0004";
        ram_buffer(47878) := X"27BD0008";
        ram_buffer(47879) := X"03E00008";
        ram_buffer(47880) := X"00000000";
        ram_buffer(47881) := X"27BDFFF8";
        ram_buffer(47882) := X"AFBE0004";
        ram_buffer(47883) := X"03A0F021";
        ram_buffer(47884) := X"8F828124";
        ram_buffer(47885) := X"03C0E821";
        ram_buffer(47886) := X"8FBE0004";
        ram_buffer(47887) := X"27BD0008";
        ram_buffer(47888) := X"03E00008";
        ram_buffer(47889) := X"00000000";
        ram_buffer(47890) := X"27BDFFF8";
        ram_buffer(47891) := X"AFBE0004";
        ram_buffer(47892) := X"03A0F021";
        ram_buffer(47893) := X"3C02100D";
        ram_buffer(47894) := X"2442D040";
        ram_buffer(47895) := X"03C0E821";
        ram_buffer(47896) := X"8FBE0004";
        ram_buffer(47897) := X"27BD0008";
        ram_buffer(47898) := X"03E00008";
        ram_buffer(47899) := X"00000000";
        ram_buffer(47900) := X"27BDFFF8";
        ram_buffer(47901) := X"AFBE0004";
        ram_buffer(47902) := X"03A0F021";
        ram_buffer(47903) := X"8F8281DC";
        ram_buffer(47904) := X"03C0E821";
        ram_buffer(47905) := X"8FBE0004";
        ram_buffer(47906) := X"27BD0008";
        ram_buffer(47907) := X"03E00008";
        ram_buffer(47908) := X"00000000";
        ram_buffer(47909) := X"27BDFFF8";
        ram_buffer(47910) := X"AFBE0004";
        ram_buffer(47911) := X"03A0F021";
        ram_buffer(47912) := X"AFC40008";
        ram_buffer(47913) := X"3C02100D";
        ram_buffer(47914) := X"2442CFE8";
        ram_buffer(47915) := X"03C0E821";
        ram_buffer(47916) := X"8FBE0004";
        ram_buffer(47917) := X"27BD0008";
        ram_buffer(47918) := X"03E00008";
        ram_buffer(47919) := X"00000000";
        ram_buffer(47920) := X"27BDFFE8";
        ram_buffer(47921) := X"AFBF0014";
        ram_buffer(47922) := X"AFBE0010";
        ram_buffer(47923) := X"03A0F021";
        ram_buffer(47924) := X"AFC40018";
        ram_buffer(47925) := X"AFC5001C";
        ram_buffer(47926) := X"8F828098";
        ram_buffer(47927) := X"8FC6001C";
        ram_buffer(47928) := X"8FC50018";
        ram_buffer(47929) := X"00402021";
        ram_buffer(47930) := X"0C02BAD4";
        ram_buffer(47931) := X"00000000";
        ram_buffer(47932) := X"03C0E821";
        ram_buffer(47933) := X"8FBF0014";
        ram_buffer(47934) := X"8FBE0010";
        ram_buffer(47935) := X"27BD0018";
        ram_buffer(47936) := X"03E00008";
        ram_buffer(47937) := X"00000000";
        ram_buffer(47938) := X"27BDFFE8";
        ram_buffer(47939) := X"AFBF0014";
        ram_buffer(47940) := X"AFBE0010";
        ram_buffer(47941) := X"03A0F021";
        ram_buffer(47942) := X"8F828098";
        ram_buffer(47943) := X"00000000";
        ram_buffer(47944) := X"00402021";
        ram_buffer(47945) := X"0C02BB25";
        ram_buffer(47946) := X"00000000";
        ram_buffer(47947) := X"03C0E821";
        ram_buffer(47948) := X"8FBF0014";
        ram_buffer(47949) := X"8FBE0010";
        ram_buffer(47950) := X"27BD0018";
        ram_buffer(47951) := X"03E00008";
        ram_buffer(47952) := X"00000000";
        ram_buffer(47953) := X"27BDFFE0";
        ram_buffer(47954) := X"AFBF001C";
        ram_buffer(47955) := X"AFBE0018";
        ram_buffer(47956) := X"03A0F021";
        ram_buffer(47957) := X"AFC40020";
        ram_buffer(47958) := X"AFC50024";
        ram_buffer(47959) := X"AFC60028";
        ram_buffer(47960) := X"AFC7002C";
        ram_buffer(47961) := X"AF8081EC";
        ram_buffer(47962) := X"8FC6002C";
        ram_buffer(47963) := X"8FC50028";
        ram_buffer(47964) := X"8FC40024";
        ram_buffer(47965) := X"0C02FBD9";
        ram_buffer(47966) := X"00000000";
        ram_buffer(47967) := X"AFC20010";
        ram_buffer(47968) := X"8FC30010";
        ram_buffer(47969) := X"2402FFFF";
        ram_buffer(47970) := X"14620009";
        ram_buffer(47971) := X"00000000";
        ram_buffer(47972) := X"8F8281EC";
        ram_buffer(47973) := X"00000000";
        ram_buffer(47974) := X"10400005";
        ram_buffer(47975) := X"00000000";
        ram_buffer(47976) := X"8F8381EC";
        ram_buffer(47977) := X"8FC20020";
        ram_buffer(47978) := X"00000000";
        ram_buffer(47979) := X"AC430000";
        ram_buffer(47980) := X"8FC20010";
        ram_buffer(47981) := X"03C0E821";
        ram_buffer(47982) := X"8FBF001C";
        ram_buffer(47983) := X"8FBE0018";
        ram_buffer(47984) := X"27BD0020";
        ram_buffer(47985) := X"03E00008";
        ram_buffer(47986) := X"00000000";
        ram_buffer(47987) := X"27BDFFD0";
        ram_buffer(47988) := X"AFBF002C";
        ram_buffer(47989) := X"AFBE0028";
        ram_buffer(47990) := X"AFB00024";
        ram_buffer(47991) := X"03A0F021";
        ram_buffer(47992) := X"AFC40030";
        ram_buffer(47993) := X"AFC50034";
        ram_buffer(47994) := X"AFC60038";
        ram_buffer(47995) := X"AFC7003C";
        ram_buffer(47996) := X"AFC00018";
        ram_buffer(47997) := X"8FC20038";
        ram_buffer(47998) := X"00000000";
        ram_buffer(47999) := X"14400013";
        ram_buffer(48000) := X"00000000";
        ram_buffer(48001) := X"8F908128";
        ram_buffer(48002) := X"0C02BAFF";
        ram_buffer(48003) := X"00000000";
        ram_buffer(48004) := X"00401821";
        ram_buffer(48005) := X"8FC20040";
        ram_buffer(48006) := X"00000000";
        ram_buffer(48007) := X"AFA20014";
        ram_buffer(48008) := X"AFA30010";
        ram_buffer(48009) := X"24070001";
        ram_buffer(48010) := X"3C02100D";
        ram_buffer(48011) := X"2446A930";
        ram_buffer(48012) := X"00002821";
        ram_buffer(48013) := X"8FC40030";
        ram_buffer(48014) := X"0200F809";
        ram_buffer(48015) := X"00000000";
        ram_buffer(48016) := X"AFC20018";
        ram_buffer(48017) := X"10000010";
        ram_buffer(48018) := X"00000000";
        ram_buffer(48019) := X"8F908128";
        ram_buffer(48020) := X"0C02BAFF";
        ram_buffer(48021) := X"00000000";
        ram_buffer(48022) := X"00401821";
        ram_buffer(48023) := X"8FC20040";
        ram_buffer(48024) := X"00000000";
        ram_buffer(48025) := X"AFA20014";
        ram_buffer(48026) := X"AFA30010";
        ram_buffer(48027) := X"8FC7003C";
        ram_buffer(48028) := X"8FC60038";
        ram_buffer(48029) := X"8FC50034";
        ram_buffer(48030) := X"8FC40030";
        ram_buffer(48031) := X"0200F809";
        ram_buffer(48032) := X"00000000";
        ram_buffer(48033) := X"AFC20018";
        ram_buffer(48034) := X"8FC30018";
        ram_buffer(48035) := X"2402FFFF";
        ram_buffer(48036) := X"1462000A";
        ram_buffer(48037) := X"00000000";
        ram_buffer(48038) := X"8FC20040";
        ram_buffer(48039) := X"00000000";
        ram_buffer(48040) := X"AC400000";
        ram_buffer(48041) := X"8FC20030";
        ram_buffer(48042) := X"2403008A";
        ram_buffer(48043) := X"AC430000";
        ram_buffer(48044) := X"2402FFFF";
        ram_buffer(48045) := X"10000002";
        ram_buffer(48046) := X"00000000";
        ram_buffer(48047) := X"8FC20018";
        ram_buffer(48048) := X"03C0E821";
        ram_buffer(48049) := X"8FBF002C";
        ram_buffer(48050) := X"8FBE0028";
        ram_buffer(48051) := X"8FB00024";
        ram_buffer(48052) := X"27BD0030";
        ram_buffer(48053) := X"03E00008";
        ram_buffer(48054) := X"00000000";
        ram_buffer(48055) := X"27BDFFD0";
        ram_buffer(48056) := X"AFBF002C";
        ram_buffer(48057) := X"AFBE0028";
        ram_buffer(48058) := X"AFB00024";
        ram_buffer(48059) := X"03A0F021";
        ram_buffer(48060) := X"AFC40030";
        ram_buffer(48061) := X"AFC50034";
        ram_buffer(48062) := X"AFC60038";
        ram_buffer(48063) := X"AFC7003C";
        ram_buffer(48064) := X"AFC00018";
        ram_buffer(48065) := X"8F828098";
        ram_buffer(48066) := X"00000000";
        ram_buffer(48067) := X"AFC2001C";
        ram_buffer(48068) := X"8FC20034";
        ram_buffer(48069) := X"00000000";
        ram_buffer(48070) := X"14400013";
        ram_buffer(48071) := X"00000000";
        ram_buffer(48072) := X"8F908128";
        ram_buffer(48073) := X"0C02BAFF";
        ram_buffer(48074) := X"00000000";
        ram_buffer(48075) := X"00401821";
        ram_buffer(48076) := X"8FC2003C";
        ram_buffer(48077) := X"00000000";
        ram_buffer(48078) := X"AFA20014";
        ram_buffer(48079) := X"AFA30010";
        ram_buffer(48080) := X"24070001";
        ram_buffer(48081) := X"3C02100D";
        ram_buffer(48082) := X"2446A930";
        ram_buffer(48083) := X"00002821";
        ram_buffer(48084) := X"8FC4001C";
        ram_buffer(48085) := X"0200F809";
        ram_buffer(48086) := X"00000000";
        ram_buffer(48087) := X"AFC20018";
        ram_buffer(48088) := X"10000010";
        ram_buffer(48089) := X"00000000";
        ram_buffer(48090) := X"8F908128";
        ram_buffer(48091) := X"0C02BAFF";
        ram_buffer(48092) := X"00000000";
        ram_buffer(48093) := X"00401821";
        ram_buffer(48094) := X"8FC2003C";
        ram_buffer(48095) := X"00000000";
        ram_buffer(48096) := X"AFA20014";
        ram_buffer(48097) := X"AFA30010";
        ram_buffer(48098) := X"8FC70038";
        ram_buffer(48099) := X"8FC60034";
        ram_buffer(48100) := X"8FC50030";
        ram_buffer(48101) := X"8FC4001C";
        ram_buffer(48102) := X"0200F809";
        ram_buffer(48103) := X"00000000";
        ram_buffer(48104) := X"AFC20018";
        ram_buffer(48105) := X"8FC30018";
        ram_buffer(48106) := X"2402FFFF";
        ram_buffer(48107) := X"1462000A";
        ram_buffer(48108) := X"00000000";
        ram_buffer(48109) := X"8FC2003C";
        ram_buffer(48110) := X"00000000";
        ram_buffer(48111) := X"AC400000";
        ram_buffer(48112) := X"8FC2001C";
        ram_buffer(48113) := X"2403008A";
        ram_buffer(48114) := X"AC430000";
        ram_buffer(48115) := X"2402FFFF";
        ram_buffer(48116) := X"10000002";
        ram_buffer(48117) := X"00000000";
        ram_buffer(48118) := X"8FC20018";
        ram_buffer(48119) := X"03C0E821";
        ram_buffer(48120) := X"8FBF002C";
        ram_buffer(48121) := X"8FBE0028";
        ram_buffer(48122) := X"8FB00024";
        ram_buffer(48123) := X"27BD0030";
        ram_buffer(48124) := X"03E00008";
        ram_buffer(48125) := X"00000000";
        ram_buffer(48126) := X"27BDFFD8";
        ram_buffer(48127) := X"AFBF0024";
        ram_buffer(48128) := X"AFBE0020";
        ram_buffer(48129) := X"AFB0001C";
        ram_buffer(48130) := X"03A0F021";
        ram_buffer(48131) := X"AFC40028";
        ram_buffer(48132) := X"AFC5002C";
        ram_buffer(48133) := X"AFC60030";
        ram_buffer(48134) := X"AFC70034";
        ram_buffer(48135) := X"8F908128";
        ram_buffer(48136) := X"0C02BAFF";
        ram_buffer(48137) := X"00000000";
        ram_buffer(48138) := X"00401821";
        ram_buffer(48139) := X"8FC20038";
        ram_buffer(48140) := X"00000000";
        ram_buffer(48141) := X"AFA20014";
        ram_buffer(48142) := X"AFA30010";
        ram_buffer(48143) := X"8FC70034";
        ram_buffer(48144) := X"8FC60030";
        ram_buffer(48145) := X"8FC5002C";
        ram_buffer(48146) := X"8FC40028";
        ram_buffer(48147) := X"0200F809";
        ram_buffer(48148) := X"00000000";
        ram_buffer(48149) := X"03C0E821";
        ram_buffer(48150) := X"8FBF0024";
        ram_buffer(48151) := X"8FBE0020";
        ram_buffer(48152) := X"8FB0001C";
        ram_buffer(48153) := X"27BD0028";
        ram_buffer(48154) := X"03E00008";
        ram_buffer(48155) := X"00000000";
        ram_buffer(48156) := X"27BDFFF0";
        ram_buffer(48157) := X"AFBE000C";
        ram_buffer(48158) := X"03A0F021";
        ram_buffer(48159) := X"AFC40010";
        ram_buffer(48160) := X"AFC50014";
        ram_buffer(48161) := X"AFC60018";
        ram_buffer(48162) := X"AFC7001C";
        ram_buffer(48163) := X"8FC20018";
        ram_buffer(48164) := X"00000000";
        ram_buffer(48165) := X"AFC20000";
        ram_buffer(48166) := X"8FC20014";
        ram_buffer(48167) := X"00000000";
        ram_buffer(48168) := X"14400003";
        ram_buffer(48169) := X"00000000";
        ram_buffer(48170) := X"27C20004";
        ram_buffer(48171) := X"AFC20014";
        ram_buffer(48172) := X"8FC20018";
        ram_buffer(48173) := X"00000000";
        ram_buffer(48174) := X"14400004";
        ram_buffer(48175) := X"00000000";
        ram_buffer(48176) := X"00001021";
        ram_buffer(48177) := X"1000001A";
        ram_buffer(48178) := X"00000000";
        ram_buffer(48179) := X"8FC2001C";
        ram_buffer(48180) := X"00000000";
        ram_buffer(48181) := X"14400004";
        ram_buffer(48182) := X"00000000";
        ram_buffer(48183) := X"2402FFFE";
        ram_buffer(48184) := X"10000013";
        ram_buffer(48185) := X"00000000";
        ram_buffer(48186) := X"8FC20000";
        ram_buffer(48187) := X"00000000";
        ram_buffer(48188) := X"90420000";
        ram_buffer(48189) := X"00000000";
        ram_buffer(48190) := X"00401821";
        ram_buffer(48191) := X"8FC20014";
        ram_buffer(48192) := X"00000000";
        ram_buffer(48193) := X"AC430000";
        ram_buffer(48194) := X"8FC20000";
        ram_buffer(48195) := X"00000000";
        ram_buffer(48196) := X"90420000";
        ram_buffer(48197) := X"00000000";
        ram_buffer(48198) := X"14400004";
        ram_buffer(48199) := X"00000000";
        ram_buffer(48200) := X"00001021";
        ram_buffer(48201) := X"10000002";
        ram_buffer(48202) := X"00000000";
        ram_buffer(48203) := X"24020001";
        ram_buffer(48204) := X"03C0E821";
        ram_buffer(48205) := X"8FBE000C";
        ram_buffer(48206) := X"27BD0010";
        ram_buffer(48207) := X"03E00008";
        ram_buffer(48208) := X"00000000";
        ram_buffer(48209) := X"27BDFFE0";
        ram_buffer(48210) := X"AFBE001C";
        ram_buffer(48211) := X"03A0F021";
        ram_buffer(48212) := X"AFC40020";
        ram_buffer(48213) := X"AFC50024";
        ram_buffer(48214) := X"AFC60028";
        ram_buffer(48215) := X"8FC20020";
        ram_buffer(48216) := X"00000000";
        ram_buffer(48217) := X"AFC20000";
        ram_buffer(48218) := X"8FC20024";
        ram_buffer(48219) := X"00000000";
        ram_buffer(48220) := X"A3C20010";
        ram_buffer(48221) := X"10000018";
        ram_buffer(48222) := X"00000000";
        ram_buffer(48223) := X"8FC20028";
        ram_buffer(48224) := X"00000000";
        ram_buffer(48225) := X"2443FFFF";
        ram_buffer(48226) := X"AFC30028";
        ram_buffer(48227) := X"14400004";
        ram_buffer(48228) := X"00000000";
        ram_buffer(48229) := X"00001021";
        ram_buffer(48230) := X"10000081";
        ram_buffer(48231) := X"00000000";
        ram_buffer(48232) := X"8FC20000";
        ram_buffer(48233) := X"00000000";
        ram_buffer(48234) := X"90420000";
        ram_buffer(48235) := X"93C30010";
        ram_buffer(48236) := X"00000000";
        ram_buffer(48237) := X"14620004";
        ram_buffer(48238) := X"00000000";
        ram_buffer(48239) := X"8FC20000";
        ram_buffer(48240) := X"10000077";
        ram_buffer(48241) := X"00000000";
        ram_buffer(48242) := X"8FC20000";
        ram_buffer(48243) := X"00000000";
        ram_buffer(48244) := X"24420001";
        ram_buffer(48245) := X"AFC20000";
        ram_buffer(48246) := X"8FC20000";
        ram_buffer(48247) := X"00000000";
        ram_buffer(48248) := X"30420003";
        ram_buffer(48249) := X"1440FFE5";
        ram_buffer(48250) := X"00000000";
        ram_buffer(48251) := X"8FC20028";
        ram_buffer(48252) := X"00000000";
        ram_buffer(48253) := X"2C420004";
        ram_buffer(48254) := X"14400062";
        ram_buffer(48255) := X"00000000";
        ram_buffer(48256) := X"8FC20000";
        ram_buffer(48257) := X"00000000";
        ram_buffer(48258) := X"AFC20004";
        ram_buffer(48259) := X"93C20010";
        ram_buffer(48260) := X"00000000";
        ram_buffer(48261) := X"00021A00";
        ram_buffer(48262) := X"93C20010";
        ram_buffer(48263) := X"00000000";
        ram_buffer(48264) := X"00621025";
        ram_buffer(48265) := X"AFC20008";
        ram_buffer(48266) := X"8FC20008";
        ram_buffer(48267) := X"00000000";
        ram_buffer(48268) := X"00021400";
        ram_buffer(48269) := X"8FC30008";
        ram_buffer(48270) := X"00000000";
        ram_buffer(48271) := X"00621025";
        ram_buffer(48272) := X"AFC20008";
        ram_buffer(48273) := X"24020020";
        ram_buffer(48274) := X"AFC2000C";
        ram_buffer(48275) := X"1000000D";
        ram_buffer(48276) := X"00000000";
        ram_buffer(48277) := X"8FC30008";
        ram_buffer(48278) := X"8FC2000C";
        ram_buffer(48279) := X"00000000";
        ram_buffer(48280) := X"00431004";
        ram_buffer(48281) := X"8FC30008";
        ram_buffer(48282) := X"00000000";
        ram_buffer(48283) := X"00621025";
        ram_buffer(48284) := X"AFC20008";
        ram_buffer(48285) := X"8FC2000C";
        ram_buffer(48286) := X"00000000";
        ram_buffer(48287) := X"00021040";
        ram_buffer(48288) := X"AFC2000C";
        ram_buffer(48289) := X"8FC2000C";
        ram_buffer(48290) := X"00000000";
        ram_buffer(48291) := X"2C420020";
        ram_buffer(48292) := X"1440FFF0";
        ram_buffer(48293) := X"00000000";
        ram_buffer(48294) := X"1000001F";
        ram_buffer(48295) := X"00000000";
        ram_buffer(48296) := X"8FC20004";
        ram_buffer(48297) := X"00000000";
        ram_buffer(48298) := X"8C430000";
        ram_buffer(48299) := X"8FC20008";
        ram_buffer(48300) := X"00000000";
        ram_buffer(48301) := X"00621826";
        ram_buffer(48302) := X"3C02FEFE";
        ram_buffer(48303) := X"3442FEFF";
        ram_buffer(48304) := X"00621821";
        ram_buffer(48305) := X"8FC20004";
        ram_buffer(48306) := X"00000000";
        ram_buffer(48307) := X"8C440000";
        ram_buffer(48308) := X"8FC20008";
        ram_buffer(48309) := X"00000000";
        ram_buffer(48310) := X"00821026";
        ram_buffer(48311) := X"00021027";
        ram_buffer(48312) := X"00621824";
        ram_buffer(48313) := X"3C028080";
        ram_buffer(48314) := X"34428080";
        ram_buffer(48315) := X"00621024";
        ram_buffer(48316) := X"14400010";
        ram_buffer(48317) := X"00000000";
        ram_buffer(48318) := X"8FC20028";
        ram_buffer(48319) := X"00000000";
        ram_buffer(48320) := X"2442FFFC";
        ram_buffer(48321) := X"AFC20028";
        ram_buffer(48322) := X"8FC20004";
        ram_buffer(48323) := X"00000000";
        ram_buffer(48324) := X"24420004";
        ram_buffer(48325) := X"AFC20004";
        ram_buffer(48326) := X"8FC20028";
        ram_buffer(48327) := X"00000000";
        ram_buffer(48328) := X"2C420004";
        ram_buffer(48329) := X"1040FFDE";
        ram_buffer(48330) := X"00000000";
        ram_buffer(48331) := X"10000002";
        ram_buffer(48332) := X"00000000";
        ram_buffer(48333) := X"00000000";
        ram_buffer(48334) := X"8FC20004";
        ram_buffer(48335) := X"00000000";
        ram_buffer(48336) := X"AFC20000";
        ram_buffer(48337) := X"1000000F";
        ram_buffer(48338) := X"00000000";
        ram_buffer(48339) := X"8FC20000";
        ram_buffer(48340) := X"00000000";
        ram_buffer(48341) := X"90420000";
        ram_buffer(48342) := X"93C30010";
        ram_buffer(48343) := X"00000000";
        ram_buffer(48344) := X"14620004";
        ram_buffer(48345) := X"00000000";
        ram_buffer(48346) := X"8FC20000";
        ram_buffer(48347) := X"1000000C";
        ram_buffer(48348) := X"00000000";
        ram_buffer(48349) := X"8FC20000";
        ram_buffer(48350) := X"00000000";
        ram_buffer(48351) := X"24420001";
        ram_buffer(48352) := X"AFC20000";
        ram_buffer(48353) := X"8FC20028";
        ram_buffer(48354) := X"00000000";
        ram_buffer(48355) := X"2443FFFF";
        ram_buffer(48356) := X"AFC30028";
        ram_buffer(48357) := X"1440FFED";
        ram_buffer(48358) := X"00000000";
        ram_buffer(48359) := X"00001021";
        ram_buffer(48360) := X"03C0E821";
        ram_buffer(48361) := X"8FBE001C";
        ram_buffer(48362) := X"27BD0020";
        ram_buffer(48363) := X"03E00008";
        ram_buffer(48364) := X"00000000";
        ram_buffer(48365) := X"27BDFFE8";
        ram_buffer(48366) := X"AFBE0014";
        ram_buffer(48367) := X"03A0F021";
        ram_buffer(48368) := X"AFC40018";
        ram_buffer(48369) := X"AFC5001C";
        ram_buffer(48370) := X"AFC60020";
        ram_buffer(48371) := X"8FC20018";
        ram_buffer(48372) := X"00000000";
        ram_buffer(48373) := X"AFC20000";
        ram_buffer(48374) := X"8FC2001C";
        ram_buffer(48375) := X"00000000";
        ram_buffer(48376) := X"AFC20004";
        ram_buffer(48377) := X"8FC30004";
        ram_buffer(48378) := X"8FC20000";
        ram_buffer(48379) := X"00000000";
        ram_buffer(48380) := X"0062102B";
        ram_buffer(48381) := X"1040002C";
        ram_buffer(48382) := X"00000000";
        ram_buffer(48383) := X"8FC30004";
        ram_buffer(48384) := X"8FC20020";
        ram_buffer(48385) := X"00000000";
        ram_buffer(48386) := X"00621821";
        ram_buffer(48387) := X"8FC20000";
        ram_buffer(48388) := X"00000000";
        ram_buffer(48389) := X"0043102B";
        ram_buffer(48390) := X"10400023";
        ram_buffer(48391) := X"00000000";
        ram_buffer(48392) := X"8FC30004";
        ram_buffer(48393) := X"8FC20020";
        ram_buffer(48394) := X"00000000";
        ram_buffer(48395) := X"00621021";
        ram_buffer(48396) := X"AFC20004";
        ram_buffer(48397) := X"8FC30000";
        ram_buffer(48398) := X"8FC20020";
        ram_buffer(48399) := X"00000000";
        ram_buffer(48400) := X"00621021";
        ram_buffer(48401) := X"AFC20000";
        ram_buffer(48402) := X"1000000F";
        ram_buffer(48403) := X"00000000";
        ram_buffer(48404) := X"8FC20000";
        ram_buffer(48405) := X"00000000";
        ram_buffer(48406) := X"2442FFFF";
        ram_buffer(48407) := X"AFC20000";
        ram_buffer(48408) := X"8FC20004";
        ram_buffer(48409) := X"00000000";
        ram_buffer(48410) := X"2442FFFF";
        ram_buffer(48411) := X"AFC20004";
        ram_buffer(48412) := X"8FC20004";
        ram_buffer(48413) := X"00000000";
        ram_buffer(48414) := X"80430000";
        ram_buffer(48415) := X"8FC20000";
        ram_buffer(48416) := X"00000000";
        ram_buffer(48417) := X"A0430000";
        ram_buffer(48418) := X"8FC20020";
        ram_buffer(48419) := X"00000000";
        ram_buffer(48420) := X"2443FFFF";
        ram_buffer(48421) := X"AFC30020";
        ram_buffer(48422) := X"1440FFED";
        ram_buffer(48423) := X"00000000";
        ram_buffer(48424) := X"10000079";
        ram_buffer(48425) := X"00000000";
        ram_buffer(48426) := X"8FC20020";
        ram_buffer(48427) := X"00000000";
        ram_buffer(48428) := X"2C420010";
        ram_buffer(48429) := X"1440006E";
        ram_buffer(48430) := X"00000000";
        ram_buffer(48431) := X"8FC30004";
        ram_buffer(48432) := X"8FC20000";
        ram_buffer(48433) := X"00000000";
        ram_buffer(48434) := X"00621025";
        ram_buffer(48435) := X"30420003";
        ram_buffer(48436) := X"14400067";
        ram_buffer(48437) := X"00000000";
        ram_buffer(48438) := X"8FC20000";
        ram_buffer(48439) := X"00000000";
        ram_buffer(48440) := X"AFC20008";
        ram_buffer(48441) := X"8FC20004";
        ram_buffer(48442) := X"00000000";
        ram_buffer(48443) := X"AFC2000C";
        ram_buffer(48444) := X"10000031";
        ram_buffer(48445) := X"00000000";
        ram_buffer(48446) := X"8FC20008";
        ram_buffer(48447) := X"00000000";
        ram_buffer(48448) := X"24430004";
        ram_buffer(48449) := X"AFC30008";
        ram_buffer(48450) := X"8FC3000C";
        ram_buffer(48451) := X"00000000";
        ram_buffer(48452) := X"24640004";
        ram_buffer(48453) := X"AFC4000C";
        ram_buffer(48454) := X"8C630000";
        ram_buffer(48455) := X"00000000";
        ram_buffer(48456) := X"AC430000";
        ram_buffer(48457) := X"8FC20008";
        ram_buffer(48458) := X"00000000";
        ram_buffer(48459) := X"24430004";
        ram_buffer(48460) := X"AFC30008";
        ram_buffer(48461) := X"8FC3000C";
        ram_buffer(48462) := X"00000000";
        ram_buffer(48463) := X"24640004";
        ram_buffer(48464) := X"AFC4000C";
        ram_buffer(48465) := X"8C630000";
        ram_buffer(48466) := X"00000000";
        ram_buffer(48467) := X"AC430000";
        ram_buffer(48468) := X"8FC20008";
        ram_buffer(48469) := X"00000000";
        ram_buffer(48470) := X"24430004";
        ram_buffer(48471) := X"AFC30008";
        ram_buffer(48472) := X"8FC3000C";
        ram_buffer(48473) := X"00000000";
        ram_buffer(48474) := X"24640004";
        ram_buffer(48475) := X"AFC4000C";
        ram_buffer(48476) := X"8C630000";
        ram_buffer(48477) := X"00000000";
        ram_buffer(48478) := X"AC430000";
        ram_buffer(48479) := X"8FC20008";
        ram_buffer(48480) := X"00000000";
        ram_buffer(48481) := X"24430004";
        ram_buffer(48482) := X"AFC30008";
        ram_buffer(48483) := X"8FC3000C";
        ram_buffer(48484) := X"00000000";
        ram_buffer(48485) := X"24640004";
        ram_buffer(48486) := X"AFC4000C";
        ram_buffer(48487) := X"8C630000";
        ram_buffer(48488) := X"00000000";
        ram_buffer(48489) := X"AC430000";
        ram_buffer(48490) := X"8FC20020";
        ram_buffer(48491) := X"00000000";
        ram_buffer(48492) := X"2442FFF0";
        ram_buffer(48493) := X"AFC20020";
        ram_buffer(48494) := X"8FC20020";
        ram_buffer(48495) := X"00000000";
        ram_buffer(48496) := X"2C420010";
        ram_buffer(48497) := X"1040FFCC";
        ram_buffer(48498) := X"00000000";
        ram_buffer(48499) := X"10000010";
        ram_buffer(48500) := X"00000000";
        ram_buffer(48501) := X"8FC20008";
        ram_buffer(48502) := X"00000000";
        ram_buffer(48503) := X"24430004";
        ram_buffer(48504) := X"AFC30008";
        ram_buffer(48505) := X"8FC3000C";
        ram_buffer(48506) := X"00000000";
        ram_buffer(48507) := X"24640004";
        ram_buffer(48508) := X"AFC4000C";
        ram_buffer(48509) := X"8C630000";
        ram_buffer(48510) := X"00000000";
        ram_buffer(48511) := X"AC430000";
        ram_buffer(48512) := X"8FC20020";
        ram_buffer(48513) := X"00000000";
        ram_buffer(48514) := X"2442FFFC";
        ram_buffer(48515) := X"AFC20020";
        ram_buffer(48516) := X"8FC20020";
        ram_buffer(48517) := X"00000000";
        ram_buffer(48518) := X"2C420004";
        ram_buffer(48519) := X"1040FFED";
        ram_buffer(48520) := X"00000000";
        ram_buffer(48521) := X"8FC20008";
        ram_buffer(48522) := X"00000000";
        ram_buffer(48523) := X"AFC20000";
        ram_buffer(48524) := X"8FC2000C";
        ram_buffer(48525) := X"00000000";
        ram_buffer(48526) := X"AFC20004";
        ram_buffer(48527) := X"1000000C";
        ram_buffer(48528) := X"00000000";
        ram_buffer(48529) := X"8FC20000";
        ram_buffer(48530) := X"00000000";
        ram_buffer(48531) := X"24430001";
        ram_buffer(48532) := X"AFC30000";
        ram_buffer(48533) := X"8FC30004";
        ram_buffer(48534) := X"00000000";
        ram_buffer(48535) := X"24640001";
        ram_buffer(48536) := X"AFC40004";
        ram_buffer(48537) := X"80630000";
        ram_buffer(48538) := X"00000000";
        ram_buffer(48539) := X"A0430000";
        ram_buffer(48540) := X"8FC20020";
        ram_buffer(48541) := X"00000000";
        ram_buffer(48542) := X"2443FFFF";
        ram_buffer(48543) := X"AFC30020";
        ram_buffer(48544) := X"1440FFF0";
        ram_buffer(48545) := X"00000000";
        ram_buffer(48546) := X"8FC20018";
        ram_buffer(48547) := X"03C0E821";
        ram_buffer(48548) := X"8FBE0014";
        ram_buffer(48549) := X"27BD0018";
        ram_buffer(48550) := X"03E00008";
        ram_buffer(48551) := X"00000000";
        ram_buffer(48552) := X"27BDFFE0";
        ram_buffer(48553) := X"AFBF001C";
        ram_buffer(48554) := X"AFBE0018";
        ram_buffer(48555) := X"03A0F021";
        ram_buffer(48556) := X"AFC40020";
        ram_buffer(48557) := X"AFC50024";
        ram_buffer(48558) := X"8FC20020";
        ram_buffer(48559) := X"00000000";
        ram_buffer(48560) := X"8C42004C";
        ram_buffer(48561) := X"00000000";
        ram_buffer(48562) := X"14400013";
        ram_buffer(48563) := X"00000000";
        ram_buffer(48564) := X"24060021";
        ram_buffer(48565) := X"24050004";
        ram_buffer(48566) := X"8FC40020";
        ram_buffer(48567) := X"0C02F251";
        ram_buffer(48568) := X"00000000";
        ram_buffer(48569) := X"00401821";
        ram_buffer(48570) := X"8FC20020";
        ram_buffer(48571) := X"00000000";
        ram_buffer(48572) := X"AC43004C";
        ram_buffer(48573) := X"8FC20020";
        ram_buffer(48574) := X"00000000";
        ram_buffer(48575) := X"8C42004C";
        ram_buffer(48576) := X"00000000";
        ram_buffer(48577) := X"14400004";
        ram_buffer(48578) := X"00000000";
        ram_buffer(48579) := X"00001021";
        ram_buffer(48580) := X"10000045";
        ram_buffer(48581) := X"00000000";
        ram_buffer(48582) := X"8FC20020";
        ram_buffer(48583) := X"00000000";
        ram_buffer(48584) := X"8C43004C";
        ram_buffer(48585) := X"8FC20024";
        ram_buffer(48586) := X"00000000";
        ram_buffer(48587) := X"00021080";
        ram_buffer(48588) := X"00621021";
        ram_buffer(48589) := X"8C420000";
        ram_buffer(48590) := X"00000000";
        ram_buffer(48591) := X"AFC20010";
        ram_buffer(48592) := X"8FC20010";
        ram_buffer(48593) := X"00000000";
        ram_buffer(48594) := X"1040000F";
        ram_buffer(48595) := X"00000000";
        ram_buffer(48596) := X"8FC20020";
        ram_buffer(48597) := X"00000000";
        ram_buffer(48598) := X"8C43004C";
        ram_buffer(48599) := X"8FC20024";
        ram_buffer(48600) := X"00000000";
        ram_buffer(48601) := X"00021080";
        ram_buffer(48602) := X"00621021";
        ram_buffer(48603) := X"8FC30010";
        ram_buffer(48604) := X"00000000";
        ram_buffer(48605) := X"8C630000";
        ram_buffer(48606) := X"00000000";
        ram_buffer(48607) := X"AC430000";
        ram_buffer(48608) := X"1000001F";
        ram_buffer(48609) := X"00000000";
        ram_buffer(48610) := X"24030001";
        ram_buffer(48611) := X"8FC20024";
        ram_buffer(48612) := X"00000000";
        ram_buffer(48613) := X"00431004";
        ram_buffer(48614) := X"AFC20014";
        ram_buffer(48615) := X"8FC20014";
        ram_buffer(48616) := X"00000000";
        ram_buffer(48617) := X"24420005";
        ram_buffer(48618) := X"00021080";
        ram_buffer(48619) := X"00403021";
        ram_buffer(48620) := X"24050001";
        ram_buffer(48621) := X"8FC40020";
        ram_buffer(48622) := X"0C02F251";
        ram_buffer(48623) := X"00000000";
        ram_buffer(48624) := X"AFC20010";
        ram_buffer(48625) := X"8FC20010";
        ram_buffer(48626) := X"00000000";
        ram_buffer(48627) := X"14400004";
        ram_buffer(48628) := X"00000000";
        ram_buffer(48629) := X"00001021";
        ram_buffer(48630) := X"10000013";
        ram_buffer(48631) := X"00000000";
        ram_buffer(48632) := X"8FC20010";
        ram_buffer(48633) := X"8FC30024";
        ram_buffer(48634) := X"00000000";
        ram_buffer(48635) := X"AC430004";
        ram_buffer(48636) := X"8FC20010";
        ram_buffer(48637) := X"8FC30014";
        ram_buffer(48638) := X"00000000";
        ram_buffer(48639) := X"AC430008";
        ram_buffer(48640) := X"8FC20010";
        ram_buffer(48641) := X"00000000";
        ram_buffer(48642) := X"AC400010";
        ram_buffer(48643) := X"8FC20010";
        ram_buffer(48644) := X"00000000";
        ram_buffer(48645) := X"8C430010";
        ram_buffer(48646) := X"8FC20010";
        ram_buffer(48647) := X"00000000";
        ram_buffer(48648) := X"AC43000C";
        ram_buffer(48649) := X"8FC20010";
        ram_buffer(48650) := X"03C0E821";
        ram_buffer(48651) := X"8FBF001C";
        ram_buffer(48652) := X"8FBE0018";
        ram_buffer(48653) := X"27BD0020";
        ram_buffer(48654) := X"03E00008";
        ram_buffer(48655) := X"00000000";
        ram_buffer(48656) := X"27BDFFF8";
        ram_buffer(48657) := X"AFBE0004";
        ram_buffer(48658) := X"03A0F021";
        ram_buffer(48659) := X"AFC40008";
        ram_buffer(48660) := X"AFC5000C";
        ram_buffer(48661) := X"8FC2000C";
        ram_buffer(48662) := X"00000000";
        ram_buffer(48663) := X"1040001A";
        ram_buffer(48664) := X"00000000";
        ram_buffer(48665) := X"8FC20008";
        ram_buffer(48666) := X"00000000";
        ram_buffer(48667) := X"8C43004C";
        ram_buffer(48668) := X"8FC2000C";
        ram_buffer(48669) := X"00000000";
        ram_buffer(48670) := X"8C420004";
        ram_buffer(48671) := X"00000000";
        ram_buffer(48672) := X"00021080";
        ram_buffer(48673) := X"00621021";
        ram_buffer(48674) := X"8C430000";
        ram_buffer(48675) := X"8FC2000C";
        ram_buffer(48676) := X"00000000";
        ram_buffer(48677) := X"AC430000";
        ram_buffer(48678) := X"8FC20008";
        ram_buffer(48679) := X"00000000";
        ram_buffer(48680) := X"8C43004C";
        ram_buffer(48681) := X"8FC2000C";
        ram_buffer(48682) := X"00000000";
        ram_buffer(48683) := X"8C420004";
        ram_buffer(48684) := X"00000000";
        ram_buffer(48685) := X"00021080";
        ram_buffer(48686) := X"00621021";
        ram_buffer(48687) := X"8FC3000C";
        ram_buffer(48688) := X"00000000";
        ram_buffer(48689) := X"AC430000";
        ram_buffer(48690) := X"00000000";
        ram_buffer(48691) := X"03C0E821";
        ram_buffer(48692) := X"8FBE0004";
        ram_buffer(48693) := X"27BD0008";
        ram_buffer(48694) := X"03E00008";
        ram_buffer(48695) := X"00000000";
        ram_buffer(48696) := X"27BDFFC8";
        ram_buffer(48697) := X"AFBF0034";
        ram_buffer(48698) := X"AFBE0030";
        ram_buffer(48699) := X"03A0F021";
        ram_buffer(48700) := X"AFC40038";
        ram_buffer(48701) := X"AFC5003C";
        ram_buffer(48702) := X"AFC60040";
        ram_buffer(48703) := X"AFC70044";
        ram_buffer(48704) := X"8FC2003C";
        ram_buffer(48705) := X"00000000";
        ram_buffer(48706) := X"8C420010";
        ram_buffer(48707) := X"00000000";
        ram_buffer(48708) := X"AFC20018";
        ram_buffer(48709) := X"8FC2003C";
        ram_buffer(48710) := X"00000000";
        ram_buffer(48711) := X"24420014";
        ram_buffer(48712) := X"AFC20014";
        ram_buffer(48713) := X"AFC00010";
        ram_buffer(48714) := X"8FC20014";
        ram_buffer(48715) := X"00000000";
        ram_buffer(48716) := X"8C420000";
        ram_buffer(48717) := X"00000000";
        ram_buffer(48718) := X"AFC2001C";
        ram_buffer(48719) := X"8FC2001C";
        ram_buffer(48720) := X"00000000";
        ram_buffer(48721) := X"3043FFFF";
        ram_buffer(48722) := X"8FC20040";
        ram_buffer(48723) := X"00000000";
        ram_buffer(48724) := X"00620018";
        ram_buffer(48725) := X"8FC20044";
        ram_buffer(48726) := X"00001812";
        ram_buffer(48727) := X"00621021";
        ram_buffer(48728) := X"AFC20020";
        ram_buffer(48729) := X"8FC2001C";
        ram_buffer(48730) := X"00000000";
        ram_buffer(48731) := X"00021C02";
        ram_buffer(48732) := X"8FC20040";
        ram_buffer(48733) := X"00000000";
        ram_buffer(48734) := X"00620018";
        ram_buffer(48735) := X"8FC20020";
        ram_buffer(48736) := X"00000000";
        ram_buffer(48737) := X"00021402";
        ram_buffer(48738) := X"00001812";
        ram_buffer(48739) := X"00621021";
        ram_buffer(48740) := X"AFC20024";
        ram_buffer(48741) := X"8FC20024";
        ram_buffer(48742) := X"00000000";
        ram_buffer(48743) := X"00021402";
        ram_buffer(48744) := X"AFC20044";
        ram_buffer(48745) := X"8FC20014";
        ram_buffer(48746) := X"00000000";
        ram_buffer(48747) := X"24430004";
        ram_buffer(48748) := X"AFC30014";
        ram_buffer(48749) := X"8FC30024";
        ram_buffer(48750) := X"00000000";
        ram_buffer(48751) := X"00032400";
        ram_buffer(48752) := X"8FC30020";
        ram_buffer(48753) := X"00000000";
        ram_buffer(48754) := X"3063FFFF";
        ram_buffer(48755) := X"00831821";
        ram_buffer(48756) := X"AC430000";
        ram_buffer(48757) := X"8FC20010";
        ram_buffer(48758) := X"00000000";
        ram_buffer(48759) := X"24420001";
        ram_buffer(48760) := X"AFC20010";
        ram_buffer(48761) := X"8FC30010";
        ram_buffer(48762) := X"8FC20018";
        ram_buffer(48763) := X"00000000";
        ram_buffer(48764) := X"0062102A";
        ram_buffer(48765) := X"1440FFCC";
        ram_buffer(48766) := X"00000000";
        ram_buffer(48767) := X"8FC20044";
        ram_buffer(48768) := X"00000000";
        ram_buffer(48769) := X"10400039";
        ram_buffer(48770) := X"00000000";
        ram_buffer(48771) := X"8FC2003C";
        ram_buffer(48772) := X"00000000";
        ram_buffer(48773) := X"8C430008";
        ram_buffer(48774) := X"8FC20018";
        ram_buffer(48775) := X"00000000";
        ram_buffer(48776) := X"0043102A";
        ram_buffer(48777) := X"14400023";
        ram_buffer(48778) := X"00000000";
        ram_buffer(48779) := X"8FC2003C";
        ram_buffer(48780) := X"00000000";
        ram_buffer(48781) := X"8C420004";
        ram_buffer(48782) := X"00000000";
        ram_buffer(48783) := X"24420001";
        ram_buffer(48784) := X"00402821";
        ram_buffer(48785) := X"8FC40038";
        ram_buffer(48786) := X"0C02BDA8";
        ram_buffer(48787) := X"00000000";
        ram_buffer(48788) := X"AFC20028";
        ram_buffer(48789) := X"8FC20028";
        ram_buffer(48790) := X"00000000";
        ram_buffer(48791) := X"2443000C";
        ram_buffer(48792) := X"8FC2003C";
        ram_buffer(48793) := X"00000000";
        ram_buffer(48794) := X"2444000C";
        ram_buffer(48795) := X"8FC2003C";
        ram_buffer(48796) := X"00000000";
        ram_buffer(48797) := X"8C420010";
        ram_buffer(48798) := X"00000000";
        ram_buffer(48799) := X"24420002";
        ram_buffer(48800) := X"00021080";
        ram_buffer(48801) := X"00403021";
        ram_buffer(48802) := X"00802821";
        ram_buffer(48803) := X"00602021";
        ram_buffer(48804) := X"0C027F93";
        ram_buffer(48805) := X"00000000";
        ram_buffer(48806) := X"8FC5003C";
        ram_buffer(48807) := X"8FC40038";
        ram_buffer(48808) := X"0C02BE10";
        ram_buffer(48809) := X"00000000";
        ram_buffer(48810) := X"8FC20028";
        ram_buffer(48811) := X"00000000";
        ram_buffer(48812) := X"AFC2003C";
        ram_buffer(48813) := X"8FC20018";
        ram_buffer(48814) := X"00000000";
        ram_buffer(48815) := X"24430001";
        ram_buffer(48816) := X"AFC30018";
        ram_buffer(48817) := X"8FC30044";
        ram_buffer(48818) := X"8FC4003C";
        ram_buffer(48819) := X"24420004";
        ram_buffer(48820) := X"00021080";
        ram_buffer(48821) := X"00821021";
        ram_buffer(48822) := X"AC430004";
        ram_buffer(48823) := X"8FC2003C";
        ram_buffer(48824) := X"8FC30018";
        ram_buffer(48825) := X"00000000";
        ram_buffer(48826) := X"AC430010";
        ram_buffer(48827) := X"8FC2003C";
        ram_buffer(48828) := X"03C0E821";
        ram_buffer(48829) := X"8FBF0034";
        ram_buffer(48830) := X"8FBE0030";
        ram_buffer(48831) := X"27BD0038";
        ram_buffer(48832) := X"03E00008";
        ram_buffer(48833) := X"00000000";
        ram_buffer(48834) := X"27BDFFD0";
        ram_buffer(48835) := X"AFBF002C";
        ram_buffer(48836) := X"AFBE0028";
        ram_buffer(48837) := X"03A0F021";
        ram_buffer(48838) := X"AFC40030";
        ram_buffer(48839) := X"AFC50034";
        ram_buffer(48840) := X"AFC60038";
        ram_buffer(48841) := X"AFC7003C";
        ram_buffer(48842) := X"8FC2003C";
        ram_buffer(48843) := X"00000000";
        ram_buffer(48844) := X"24430008";
        ram_buffer(48845) := X"24020009";
        ram_buffer(48846) := X"14400002";
        ram_buffer(48847) := X"0062001A";
        ram_buffer(48848) := X"0007000D";
        ram_buffer(48849) := X"00001010";
        ram_buffer(48850) := X"00001012";
        ram_buffer(48851) := X"AFC20020";
        ram_buffer(48852) := X"AFC00018";
        ram_buffer(48853) := X"24020001";
        ram_buffer(48854) := X"AFC2001C";
        ram_buffer(48855) := X"10000009";
        ram_buffer(48856) := X"00000000";
        ram_buffer(48857) := X"8FC2001C";
        ram_buffer(48858) := X"00000000";
        ram_buffer(48859) := X"00021040";
        ram_buffer(48860) := X"AFC2001C";
        ram_buffer(48861) := X"8FC20018";
        ram_buffer(48862) := X"00000000";
        ram_buffer(48863) := X"24420001";
        ram_buffer(48864) := X"AFC20018";
        ram_buffer(48865) := X"8FC30020";
        ram_buffer(48866) := X"8FC2001C";
        ram_buffer(48867) := X"00000000";
        ram_buffer(48868) := X"0043102A";
        ram_buffer(48869) := X"1440FFF3";
        ram_buffer(48870) := X"00000000";
        ram_buffer(48871) := X"8FC50018";
        ram_buffer(48872) := X"8FC40030";
        ram_buffer(48873) := X"0C02BDA8";
        ram_buffer(48874) := X"00000000";
        ram_buffer(48875) := X"AFC20010";
        ram_buffer(48876) := X"8FC20010";
        ram_buffer(48877) := X"8FC30040";
        ram_buffer(48878) := X"00000000";
        ram_buffer(48879) := X"AC430014";
        ram_buffer(48880) := X"8FC20010";
        ram_buffer(48881) := X"24030001";
        ram_buffer(48882) := X"AC430010";
        ram_buffer(48883) := X"24020009";
        ram_buffer(48884) := X"AFC20014";
        ram_buffer(48885) := X"8FC20038";
        ram_buffer(48886) := X"00000000";
        ram_buffer(48887) := X"2842000A";
        ram_buffer(48888) := X"14400023";
        ram_buffer(48889) := X"00000000";
        ram_buffer(48890) := X"8FC20034";
        ram_buffer(48891) := X"00000000";
        ram_buffer(48892) := X"24420009";
        ram_buffer(48893) := X"AFC20034";
        ram_buffer(48894) := X"8FC20034";
        ram_buffer(48895) := X"00000000";
        ram_buffer(48896) := X"24430001";
        ram_buffer(48897) := X"AFC30034";
        ram_buffer(48898) := X"80420000";
        ram_buffer(48899) := X"00000000";
        ram_buffer(48900) := X"2442FFD0";
        ram_buffer(48901) := X"00403821";
        ram_buffer(48902) := X"2406000A";
        ram_buffer(48903) := X"8FC50010";
        ram_buffer(48904) := X"8FC40030";
        ram_buffer(48905) := X"0C02BE38";
        ram_buffer(48906) := X"00000000";
        ram_buffer(48907) := X"AFC20010";
        ram_buffer(48908) := X"8FC20014";
        ram_buffer(48909) := X"00000000";
        ram_buffer(48910) := X"24420001";
        ram_buffer(48911) := X"AFC20014";
        ram_buffer(48912) := X"8FC30014";
        ram_buffer(48913) := X"8FC20038";
        ram_buffer(48914) := X"00000000";
        ram_buffer(48915) := X"0062102A";
        ram_buffer(48916) := X"1440FFE9";
        ram_buffer(48917) := X"00000000";
        ram_buffer(48918) := X"8FC20034";
        ram_buffer(48919) := X"00000000";
        ram_buffer(48920) := X"24420001";
        ram_buffer(48921) := X"AFC20034";
        ram_buffer(48922) := X"10000019";
        ram_buffer(48923) := X"00000000";
        ram_buffer(48924) := X"8FC20034";
        ram_buffer(48925) := X"00000000";
        ram_buffer(48926) := X"2442000A";
        ram_buffer(48927) := X"AFC20034";
        ram_buffer(48928) := X"10000013";
        ram_buffer(48929) := X"00000000";
        ram_buffer(48930) := X"8FC20034";
        ram_buffer(48931) := X"00000000";
        ram_buffer(48932) := X"24430001";
        ram_buffer(48933) := X"AFC30034";
        ram_buffer(48934) := X"80420000";
        ram_buffer(48935) := X"00000000";
        ram_buffer(48936) := X"2442FFD0";
        ram_buffer(48937) := X"00403821";
        ram_buffer(48938) := X"2406000A";
        ram_buffer(48939) := X"8FC50010";
        ram_buffer(48940) := X"8FC40030";
        ram_buffer(48941) := X"0C02BE38";
        ram_buffer(48942) := X"00000000";
        ram_buffer(48943) := X"AFC20010";
        ram_buffer(48944) := X"8FC20014";
        ram_buffer(48945) := X"00000000";
        ram_buffer(48946) := X"24420001";
        ram_buffer(48947) := X"AFC20014";
        ram_buffer(48948) := X"8FC30014";
        ram_buffer(48949) := X"8FC2003C";
        ram_buffer(48950) := X"00000000";
        ram_buffer(48951) := X"0062102A";
        ram_buffer(48952) := X"1440FFE9";
        ram_buffer(48953) := X"00000000";
        ram_buffer(48954) := X"8FC20010";
        ram_buffer(48955) := X"03C0E821";
        ram_buffer(48956) := X"8FBF002C";
        ram_buffer(48957) := X"8FBE0028";
        ram_buffer(48958) := X"27BD0030";
        ram_buffer(48959) := X"03E00008";
        ram_buffer(48960) := X"00000000";
        ram_buffer(48961) := X"27BDFFF8";
        ram_buffer(48962) := X"AFBE0004";
        ram_buffer(48963) := X"AFB00000";
        ram_buffer(48964) := X"03A0F021";
        ram_buffer(48965) := X"00801021";
        ram_buffer(48966) := X"00008021";
        ram_buffer(48967) := X"3C03FFFF";
        ram_buffer(48968) := X"00431824";
        ram_buffer(48969) := X"14600003";
        ram_buffer(48970) := X"00000000";
        ram_buffer(48971) := X"24100010";
        ram_buffer(48972) := X"00021400";
        ram_buffer(48973) := X"3C03FF00";
        ram_buffer(48974) := X"00431824";
        ram_buffer(48975) := X"14600003";
        ram_buffer(48976) := X"00000000";
        ram_buffer(48977) := X"26100008";
        ram_buffer(48978) := X"00021200";
        ram_buffer(48979) := X"3C03F000";
        ram_buffer(48980) := X"00431824";
        ram_buffer(48981) := X"14600003";
        ram_buffer(48982) := X"00000000";
        ram_buffer(48983) := X"26100004";
        ram_buffer(48984) := X"00021100";
        ram_buffer(48985) := X"3C03C000";
        ram_buffer(48986) := X"00431824";
        ram_buffer(48987) := X"14600003";
        ram_buffer(48988) := X"00000000";
        ram_buffer(48989) := X"26100002";
        ram_buffer(48990) := X"00021080";
        ram_buffer(48991) := X"00401821";
        ram_buffer(48992) := X"04600009";
        ram_buffer(48993) := X"00000000";
        ram_buffer(48994) := X"26100001";
        ram_buffer(48995) := X"3C034000";
        ram_buffer(48996) := X"00431024";
        ram_buffer(48997) := X"14400004";
        ram_buffer(48998) := X"00000000";
        ram_buffer(48999) := X"24020020";
        ram_buffer(49000) := X"10000002";
        ram_buffer(49001) := X"00000000";
        ram_buffer(49002) := X"02001021";
        ram_buffer(49003) := X"03C0E821";
        ram_buffer(49004) := X"8FBE0004";
        ram_buffer(49005) := X"8FB00000";
        ram_buffer(49006) := X"27BD0008";
        ram_buffer(49007) := X"03E00008";
        ram_buffer(49008) := X"00000000";
        ram_buffer(49009) := X"27BDFFF0";
        ram_buffer(49010) := X"AFBE000C";
        ram_buffer(49011) := X"AFB10008";
        ram_buffer(49012) := X"AFB00004";
        ram_buffer(49013) := X"03A0F021";
        ram_buffer(49014) := X"AFC40010";
        ram_buffer(49015) := X"8FC20010";
        ram_buffer(49016) := X"00000000";
        ram_buffer(49017) := X"8C500000";
        ram_buffer(49018) := X"00000000";
        ram_buffer(49019) := X"32020007";
        ram_buffer(49020) := X"10400018";
        ram_buffer(49021) := X"00000000";
        ram_buffer(49022) := X"32020001";
        ram_buffer(49023) := X"10400004";
        ram_buffer(49024) := X"00000000";
        ram_buffer(49025) := X"00001021";
        ram_buffer(49026) := X"10000035";
        ram_buffer(49027) := X"00000000";
        ram_buffer(49028) := X"32020002";
        ram_buffer(49029) := X"10400008";
        ram_buffer(49030) := X"00000000";
        ram_buffer(49031) := X"00101842";
        ram_buffer(49032) := X"8FC20010";
        ram_buffer(49033) := X"00000000";
        ram_buffer(49034) := X"AC430000";
        ram_buffer(49035) := X"24020001";
        ram_buffer(49036) := X"1000002B";
        ram_buffer(49037) := X"00000000";
        ram_buffer(49038) := X"00101882";
        ram_buffer(49039) := X"8FC20010";
        ram_buffer(49040) := X"00000000";
        ram_buffer(49041) := X"AC430000";
        ram_buffer(49042) := X"24020002";
        ram_buffer(49043) := X"10000024";
        ram_buffer(49044) := X"00000000";
        ram_buffer(49045) := X"00008821";
        ram_buffer(49046) := X"3202FFFF";
        ram_buffer(49047) := X"14400003";
        ram_buffer(49048) := X"00000000";
        ram_buffer(49049) := X"24110010";
        ram_buffer(49050) := X"00108402";
        ram_buffer(49051) := X"320200FF";
        ram_buffer(49052) := X"14400003";
        ram_buffer(49053) := X"00000000";
        ram_buffer(49054) := X"26310008";
        ram_buffer(49055) := X"00108202";
        ram_buffer(49056) := X"3202000F";
        ram_buffer(49057) := X"14400003";
        ram_buffer(49058) := X"00000000";
        ram_buffer(49059) := X"26310004";
        ram_buffer(49060) := X"00108102";
        ram_buffer(49061) := X"32020003";
        ram_buffer(49062) := X"14400003";
        ram_buffer(49063) := X"00000000";
        ram_buffer(49064) := X"26310002";
        ram_buffer(49065) := X"00108082";
        ram_buffer(49066) := X"32020001";
        ram_buffer(49067) := X"14400008";
        ram_buffer(49068) := X"00000000";
        ram_buffer(49069) := X"26310001";
        ram_buffer(49070) := X"00108042";
        ram_buffer(49071) := X"16000004";
        ram_buffer(49072) := X"00000000";
        ram_buffer(49073) := X"24020020";
        ram_buffer(49074) := X"10000005";
        ram_buffer(49075) := X"00000000";
        ram_buffer(49076) := X"8FC20010";
        ram_buffer(49077) := X"00000000";
        ram_buffer(49078) := X"AC500000";
        ram_buffer(49079) := X"02201021";
        ram_buffer(49080) := X"03C0E821";
        ram_buffer(49081) := X"8FBE000C";
        ram_buffer(49082) := X"8FB10008";
        ram_buffer(49083) := X"8FB00004";
        ram_buffer(49084) := X"27BD0010";
        ram_buffer(49085) := X"03E00008";
        ram_buffer(49086) := X"00000000";
        ram_buffer(49087) := X"27BDFFE0";
        ram_buffer(49088) := X"AFBF001C";
        ram_buffer(49089) := X"AFBE0018";
        ram_buffer(49090) := X"03A0F021";
        ram_buffer(49091) := X"AFC40020";
        ram_buffer(49092) := X"AFC50024";
        ram_buffer(49093) := X"24050001";
        ram_buffer(49094) := X"8FC40020";
        ram_buffer(49095) := X"0C02BDA8";
        ram_buffer(49096) := X"00000000";
        ram_buffer(49097) := X"AFC20010";
        ram_buffer(49098) := X"8FC30024";
        ram_buffer(49099) := X"8FC20010";
        ram_buffer(49100) := X"00000000";
        ram_buffer(49101) := X"AC430014";
        ram_buffer(49102) := X"8FC20010";
        ram_buffer(49103) := X"24030001";
        ram_buffer(49104) := X"AC430010";
        ram_buffer(49105) := X"8FC20010";
        ram_buffer(49106) := X"03C0E821";
        ram_buffer(49107) := X"8FBF001C";
        ram_buffer(49108) := X"8FBE0018";
        ram_buffer(49109) := X"27BD0020";
        ram_buffer(49110) := X"03E00008";
        ram_buffer(49111) := X"00000000";
        ram_buffer(49112) := X"27BDFFA8";
        ram_buffer(49113) := X"AFBF0054";
        ram_buffer(49114) := X"AFBE0050";
        ram_buffer(49115) := X"03A0F021";
        ram_buffer(49116) := X"AFC40058";
        ram_buffer(49117) := X"AFC5005C";
        ram_buffer(49118) := X"AFC60060";
        ram_buffer(49119) := X"8FC2005C";
        ram_buffer(49120) := X"00000000";
        ram_buffer(49121) := X"8C430010";
        ram_buffer(49122) := X"8FC20060";
        ram_buffer(49123) := X"00000000";
        ram_buffer(49124) := X"8C420010";
        ram_buffer(49125) := X"00000000";
        ram_buffer(49126) := X"0062102A";
        ram_buffer(49127) := X"1040000A";
        ram_buffer(49128) := X"00000000";
        ram_buffer(49129) := X"8FC2005C";
        ram_buffer(49130) := X"00000000";
        ram_buffer(49131) := X"AFC20030";
        ram_buffer(49132) := X"8FC20060";
        ram_buffer(49133) := X"00000000";
        ram_buffer(49134) := X"AFC2005C";
        ram_buffer(49135) := X"8FC20030";
        ram_buffer(49136) := X"00000000";
        ram_buffer(49137) := X"AFC20060";
        ram_buffer(49138) := X"8FC2005C";
        ram_buffer(49139) := X"00000000";
        ram_buffer(49140) := X"8C420004";
        ram_buffer(49141) := X"00000000";
        ram_buffer(49142) := X"AFC20010";
        ram_buffer(49143) := X"8FC2005C";
        ram_buffer(49144) := X"00000000";
        ram_buffer(49145) := X"8C420010";
        ram_buffer(49146) := X"00000000";
        ram_buffer(49147) := X"AFC20034";
        ram_buffer(49148) := X"8FC20060";
        ram_buffer(49149) := X"00000000";
        ram_buffer(49150) := X"8C420010";
        ram_buffer(49151) := X"00000000";
        ram_buffer(49152) := X"AFC20038";
        ram_buffer(49153) := X"8FC30034";
        ram_buffer(49154) := X"8FC20038";
        ram_buffer(49155) := X"00000000";
        ram_buffer(49156) := X"00621021";
        ram_buffer(49157) := X"AFC20014";
        ram_buffer(49158) := X"8FC2005C";
        ram_buffer(49159) := X"00000000";
        ram_buffer(49160) := X"8C430008";
        ram_buffer(49161) := X"8FC20014";
        ram_buffer(49162) := X"00000000";
        ram_buffer(49163) := X"0062102A";
        ram_buffer(49164) := X"10400005";
        ram_buffer(49165) := X"00000000";
        ram_buffer(49166) := X"8FC20010";
        ram_buffer(49167) := X"00000000";
        ram_buffer(49168) := X"24420001";
        ram_buffer(49169) := X"AFC20010";
        ram_buffer(49170) := X"8FC50010";
        ram_buffer(49171) := X"8FC40058";
        ram_buffer(49172) := X"0C02BDA8";
        ram_buffer(49173) := X"00000000";
        ram_buffer(49174) := X"AFC20030";
        ram_buffer(49175) := X"8FC20030";
        ram_buffer(49176) := X"00000000";
        ram_buffer(49177) := X"24420014";
        ram_buffer(49178) := X"AFC2001C";
        ram_buffer(49179) := X"8FC20014";
        ram_buffer(49180) := X"00000000";
        ram_buffer(49181) := X"00021080";
        ram_buffer(49182) := X"8FC3001C";
        ram_buffer(49183) := X"00000000";
        ram_buffer(49184) := X"00621021";
        ram_buffer(49185) := X"AFC2003C";
        ram_buffer(49186) := X"10000008";
        ram_buffer(49187) := X"00000000";
        ram_buffer(49188) := X"8FC2001C";
        ram_buffer(49189) := X"00000000";
        ram_buffer(49190) := X"AC400000";
        ram_buffer(49191) := X"8FC2001C";
        ram_buffer(49192) := X"00000000";
        ram_buffer(49193) := X"24420004";
        ram_buffer(49194) := X"AFC2001C";
        ram_buffer(49195) := X"8FC3001C";
        ram_buffer(49196) := X"8FC2003C";
        ram_buffer(49197) := X"00000000";
        ram_buffer(49198) := X"0062102B";
        ram_buffer(49199) := X"1440FFF4";
        ram_buffer(49200) := X"00000000";
        ram_buffer(49201) := X"8FC2005C";
        ram_buffer(49202) := X"00000000";
        ram_buffer(49203) := X"24420014";
        ram_buffer(49204) := X"AFC2003C";
        ram_buffer(49205) := X"8FC20034";
        ram_buffer(49206) := X"00000000";
        ram_buffer(49207) := X"00021080";
        ram_buffer(49208) := X"8FC3003C";
        ram_buffer(49209) := X"00000000";
        ram_buffer(49210) := X"00621021";
        ram_buffer(49211) := X"AFC20040";
        ram_buffer(49212) := X"8FC20060";
        ram_buffer(49213) := X"00000000";
        ram_buffer(49214) := X"24420014";
        ram_buffer(49215) := X"AFC20020";
        ram_buffer(49216) := X"8FC20038";
        ram_buffer(49217) := X"00000000";
        ram_buffer(49218) := X"00021080";
        ram_buffer(49219) := X"8FC30020";
        ram_buffer(49220) := X"00000000";
        ram_buffer(49221) := X"00621021";
        ram_buffer(49222) := X"AFC20044";
        ram_buffer(49223) := X"8FC20030";
        ram_buffer(49224) := X"00000000";
        ram_buffer(49225) := X"24420014";
        ram_buffer(49226) := X"AFC20028";
        ram_buffer(49227) := X"100000BC";
        ram_buffer(49228) := X"00000000";
        ram_buffer(49229) := X"8FC20020";
        ram_buffer(49230) := X"00000000";
        ram_buffer(49231) := X"8C420000";
        ram_buffer(49232) := X"00000000";
        ram_buffer(49233) := X"3042FFFF";
        ram_buffer(49234) := X"AFC20048";
        ram_buffer(49235) := X"8FC20048";
        ram_buffer(49236) := X"00000000";
        ram_buffer(49237) := X"1040004E";
        ram_buffer(49238) := X"00000000";
        ram_buffer(49239) := X"8FC2003C";
        ram_buffer(49240) := X"00000000";
        ram_buffer(49241) := X"AFC2001C";
        ram_buffer(49242) := X"8FC20028";
        ram_buffer(49243) := X"00000000";
        ram_buffer(49244) := X"AFC20024";
        ram_buffer(49245) := X"AFC00018";
        ram_buffer(49246) := X"8FC2001C";
        ram_buffer(49247) := X"00000000";
        ram_buffer(49248) := X"8C420000";
        ram_buffer(49249) := X"00000000";
        ram_buffer(49250) := X"3043FFFF";
        ram_buffer(49251) := X"8FC20048";
        ram_buffer(49252) := X"00000000";
        ram_buffer(49253) := X"00620018";
        ram_buffer(49254) := X"8FC20024";
        ram_buffer(49255) := X"00000000";
        ram_buffer(49256) := X"8C420000";
        ram_buffer(49257) := X"00000000";
        ram_buffer(49258) := X"3042FFFF";
        ram_buffer(49259) := X"00001812";
        ram_buffer(49260) := X"00621821";
        ram_buffer(49261) := X"8FC20018";
        ram_buffer(49262) := X"00000000";
        ram_buffer(49263) := X"00621021";
        ram_buffer(49264) := X"AFC2004C";
        ram_buffer(49265) := X"8FC2004C";
        ram_buffer(49266) := X"00000000";
        ram_buffer(49267) := X"00021402";
        ram_buffer(49268) := X"AFC20018";
        ram_buffer(49269) := X"8FC2001C";
        ram_buffer(49270) := X"00000000";
        ram_buffer(49271) := X"24430004";
        ram_buffer(49272) := X"AFC3001C";
        ram_buffer(49273) := X"8C420000";
        ram_buffer(49274) := X"00000000";
        ram_buffer(49275) := X"00021C02";
        ram_buffer(49276) := X"8FC20048";
        ram_buffer(49277) := X"00000000";
        ram_buffer(49278) := X"00620018";
        ram_buffer(49279) := X"8FC20024";
        ram_buffer(49280) := X"00000000";
        ram_buffer(49281) := X"8C420000";
        ram_buffer(49282) := X"00000000";
        ram_buffer(49283) := X"00021402";
        ram_buffer(49284) := X"00001812";
        ram_buffer(49285) := X"00621821";
        ram_buffer(49286) := X"8FC20018";
        ram_buffer(49287) := X"00000000";
        ram_buffer(49288) := X"00621021";
        ram_buffer(49289) := X"AFC2002C";
        ram_buffer(49290) := X"8FC2002C";
        ram_buffer(49291) := X"00000000";
        ram_buffer(49292) := X"00021402";
        ram_buffer(49293) := X"AFC20018";
        ram_buffer(49294) := X"8FC20024";
        ram_buffer(49295) := X"00000000";
        ram_buffer(49296) := X"24430004";
        ram_buffer(49297) := X"AFC30024";
        ram_buffer(49298) := X"8FC3002C";
        ram_buffer(49299) := X"00000000";
        ram_buffer(49300) := X"00032400";
        ram_buffer(49301) := X"8FC3004C";
        ram_buffer(49302) := X"00000000";
        ram_buffer(49303) := X"3063FFFF";
        ram_buffer(49304) := X"00831825";
        ram_buffer(49305) := X"AC430000";
        ram_buffer(49306) := X"8FC3001C";
        ram_buffer(49307) := X"8FC20040";
        ram_buffer(49308) := X"00000000";
        ram_buffer(49309) := X"0062102B";
        ram_buffer(49310) := X"1440FFBF";
        ram_buffer(49311) := X"00000000";
        ram_buffer(49312) := X"8FC20024";
        ram_buffer(49313) := X"8FC30018";
        ram_buffer(49314) := X"00000000";
        ram_buffer(49315) := X"AC430000";
        ram_buffer(49316) := X"8FC20020";
        ram_buffer(49317) := X"00000000";
        ram_buffer(49318) := X"8C420000";
        ram_buffer(49319) := X"00000000";
        ram_buffer(49320) := X"00021402";
        ram_buffer(49321) := X"AFC20048";
        ram_buffer(49322) := X"8FC20048";
        ram_buffer(49323) := X"00000000";
        ram_buffer(49324) := X"10400053";
        ram_buffer(49325) := X"00000000";
        ram_buffer(49326) := X"8FC2003C";
        ram_buffer(49327) := X"00000000";
        ram_buffer(49328) := X"AFC2001C";
        ram_buffer(49329) := X"8FC20028";
        ram_buffer(49330) := X"00000000";
        ram_buffer(49331) := X"AFC20024";
        ram_buffer(49332) := X"AFC00018";
        ram_buffer(49333) := X"8FC20024";
        ram_buffer(49334) := X"00000000";
        ram_buffer(49335) := X"8C420000";
        ram_buffer(49336) := X"00000000";
        ram_buffer(49337) := X"AFC2002C";
        ram_buffer(49338) := X"8FC2001C";
        ram_buffer(49339) := X"00000000";
        ram_buffer(49340) := X"8C420000";
        ram_buffer(49341) := X"00000000";
        ram_buffer(49342) := X"3043FFFF";
        ram_buffer(49343) := X"8FC20048";
        ram_buffer(49344) := X"00000000";
        ram_buffer(49345) := X"00620018";
        ram_buffer(49346) := X"8FC20024";
        ram_buffer(49347) := X"00000000";
        ram_buffer(49348) := X"8C420000";
        ram_buffer(49349) := X"00000000";
        ram_buffer(49350) := X"00021402";
        ram_buffer(49351) := X"00001812";
        ram_buffer(49352) := X"00621821";
        ram_buffer(49353) := X"8FC20018";
        ram_buffer(49354) := X"00000000";
        ram_buffer(49355) := X"00621021";
        ram_buffer(49356) := X"AFC2004C";
        ram_buffer(49357) := X"8FC2004C";
        ram_buffer(49358) := X"00000000";
        ram_buffer(49359) := X"00021402";
        ram_buffer(49360) := X"AFC20018";
        ram_buffer(49361) := X"8FC20024";
        ram_buffer(49362) := X"00000000";
        ram_buffer(49363) := X"24430004";
        ram_buffer(49364) := X"AFC30024";
        ram_buffer(49365) := X"8FC3004C";
        ram_buffer(49366) := X"00000000";
        ram_buffer(49367) := X"00032400";
        ram_buffer(49368) := X"8FC3002C";
        ram_buffer(49369) := X"00000000";
        ram_buffer(49370) := X"3063FFFF";
        ram_buffer(49371) := X"00831825";
        ram_buffer(49372) := X"AC430000";
        ram_buffer(49373) := X"8FC2001C";
        ram_buffer(49374) := X"00000000";
        ram_buffer(49375) := X"24430004";
        ram_buffer(49376) := X"AFC3001C";
        ram_buffer(49377) := X"8C420000";
        ram_buffer(49378) := X"00000000";
        ram_buffer(49379) := X"00021C02";
        ram_buffer(49380) := X"8FC20048";
        ram_buffer(49381) := X"00000000";
        ram_buffer(49382) := X"00620018";
        ram_buffer(49383) := X"8FC20024";
        ram_buffer(49384) := X"00000000";
        ram_buffer(49385) := X"8C420000";
        ram_buffer(49386) := X"00000000";
        ram_buffer(49387) := X"3042FFFF";
        ram_buffer(49388) := X"00001812";
        ram_buffer(49389) := X"00621821";
        ram_buffer(49390) := X"8FC20018";
        ram_buffer(49391) := X"00000000";
        ram_buffer(49392) := X"00621021";
        ram_buffer(49393) := X"AFC2002C";
        ram_buffer(49394) := X"8FC2002C";
        ram_buffer(49395) := X"00000000";
        ram_buffer(49396) := X"00021402";
        ram_buffer(49397) := X"AFC20018";
        ram_buffer(49398) := X"8FC3001C";
        ram_buffer(49399) := X"8FC20040";
        ram_buffer(49400) := X"00000000";
        ram_buffer(49401) := X"0062102B";
        ram_buffer(49402) := X"1440FFBF";
        ram_buffer(49403) := X"00000000";
        ram_buffer(49404) := X"8FC20024";
        ram_buffer(49405) := X"8FC3002C";
        ram_buffer(49406) := X"00000000";
        ram_buffer(49407) := X"AC430000";
        ram_buffer(49408) := X"8FC20020";
        ram_buffer(49409) := X"00000000";
        ram_buffer(49410) := X"24420004";
        ram_buffer(49411) := X"AFC20020";
        ram_buffer(49412) := X"8FC20028";
        ram_buffer(49413) := X"00000000";
        ram_buffer(49414) := X"24420004";
        ram_buffer(49415) := X"AFC20028";
        ram_buffer(49416) := X"8FC30020";
        ram_buffer(49417) := X"8FC20044";
        ram_buffer(49418) := X"00000000";
        ram_buffer(49419) := X"0062102B";
        ram_buffer(49420) := X"1440FF40";
        ram_buffer(49421) := X"00000000";
        ram_buffer(49422) := X"8FC20030";
        ram_buffer(49423) := X"00000000";
        ram_buffer(49424) := X"24420014";
        ram_buffer(49425) := X"AFC20028";
        ram_buffer(49426) := X"8FC20014";
        ram_buffer(49427) := X"00000000";
        ram_buffer(49428) := X"00021080";
        ram_buffer(49429) := X"8FC30028";
        ram_buffer(49430) := X"00000000";
        ram_buffer(49431) := X"00621021";
        ram_buffer(49432) := X"AFC20024";
        ram_buffer(49433) := X"10000005";
        ram_buffer(49434) := X"00000000";
        ram_buffer(49435) := X"8FC20014";
        ram_buffer(49436) := X"00000000";
        ram_buffer(49437) := X"2442FFFF";
        ram_buffer(49438) := X"AFC20014";
        ram_buffer(49439) := X"8FC20014";
        ram_buffer(49440) := X"00000000";
        ram_buffer(49441) := X"1840000B";
        ram_buffer(49442) := X"00000000";
        ram_buffer(49443) := X"8FC20024";
        ram_buffer(49444) := X"00000000";
        ram_buffer(49445) := X"2442FFFC";
        ram_buffer(49446) := X"AFC20024";
        ram_buffer(49447) := X"8FC20024";
        ram_buffer(49448) := X"00000000";
        ram_buffer(49449) := X"8C420000";
        ram_buffer(49450) := X"00000000";
        ram_buffer(49451) := X"1040FFEF";
        ram_buffer(49452) := X"00000000";
        ram_buffer(49453) := X"8FC20030";
        ram_buffer(49454) := X"8FC30014";
        ram_buffer(49455) := X"00000000";
        ram_buffer(49456) := X"AC430010";
        ram_buffer(49457) := X"8FC20030";
        ram_buffer(49458) := X"03C0E821";
        ram_buffer(49459) := X"8FBF0054";
        ram_buffer(49460) := X"8FBE0050";
        ram_buffer(49461) := X"27BD0058";
        ram_buffer(49462) := X"03E00008";
        ram_buffer(49463) := X"00000000";
        ram_buffer(49464) := X"27BDFFD8";
        ram_buffer(49465) := X"AFBF0024";
        ram_buffer(49466) := X"AFBE0020";
        ram_buffer(49467) := X"03A0F021";
        ram_buffer(49468) := X"AFC40028";
        ram_buffer(49469) := X"AFC5002C";
        ram_buffer(49470) := X"AFC60030";
        ram_buffer(49471) := X"8FC20030";
        ram_buffer(49472) := X"00000000";
        ram_buffer(49473) := X"30420003";
        ram_buffer(49474) := X"AFC20018";
        ram_buffer(49475) := X"8FC20018";
        ram_buffer(49476) := X"00000000";
        ram_buffer(49477) := X"10400010";
        ram_buffer(49478) := X"00000000";
        ram_buffer(49479) := X"8FC20018";
        ram_buffer(49480) := X"00000000";
        ram_buffer(49481) := X"2443FFFF";
        ram_buffer(49482) := X"3C02100D";
        ram_buffer(49483) := X"00031880";
        ram_buffer(49484) := X"2442AA50";
        ram_buffer(49485) := X"00621021";
        ram_buffer(49486) := X"8C420000";
        ram_buffer(49487) := X"00003821";
        ram_buffer(49488) := X"00403021";
        ram_buffer(49489) := X"8FC5002C";
        ram_buffer(49490) := X"8FC40028";
        ram_buffer(49491) := X"0C02BE38";
        ram_buffer(49492) := X"00000000";
        ram_buffer(49493) := X"AFC2002C";
        ram_buffer(49494) := X"8FC20030";
        ram_buffer(49495) := X"00000000";
        ram_buffer(49496) := X"00021083";
        ram_buffer(49497) := X"AFC20030";
        ram_buffer(49498) := X"8FC20030";
        ram_buffer(49499) := X"00000000";
        ram_buffer(49500) := X"14400004";
        ram_buffer(49501) := X"00000000";
        ram_buffer(49502) := X"8FC2002C";
        ram_buffer(49503) := X"10000055";
        ram_buffer(49504) := X"00000000";
        ram_buffer(49505) := X"8FC20028";
        ram_buffer(49506) := X"00000000";
        ram_buffer(49507) := X"8C420048";
        ram_buffer(49508) := X"00000000";
        ram_buffer(49509) := X"AFC20010";
        ram_buffer(49510) := X"8FC20010";
        ram_buffer(49511) := X"00000000";
        ram_buffer(49512) := X"14400011";
        ram_buffer(49513) := X"00000000";
        ram_buffer(49514) := X"24050271";
        ram_buffer(49515) := X"8FC40028";
        ram_buffer(49516) := X"0C02BFBF";
        ram_buffer(49517) := X"00000000";
        ram_buffer(49518) := X"00401821";
        ram_buffer(49519) := X"8FC20028";
        ram_buffer(49520) := X"00000000";
        ram_buffer(49521) := X"AC430048";
        ram_buffer(49522) := X"8FC20028";
        ram_buffer(49523) := X"00000000";
        ram_buffer(49524) := X"8C420048";
        ram_buffer(49525) := X"00000000";
        ram_buffer(49526) := X"AFC20010";
        ram_buffer(49527) := X"8FC20010";
        ram_buffer(49528) := X"00000000";
        ram_buffer(49529) := X"AC400000";
        ram_buffer(49530) := X"8FC20030";
        ram_buffer(49531) := X"00000000";
        ram_buffer(49532) := X"30420001";
        ram_buffer(49533) := X"1040000E";
        ram_buffer(49534) := X"00000000";
        ram_buffer(49535) := X"8FC60010";
        ram_buffer(49536) := X"8FC5002C";
        ram_buffer(49537) := X"8FC40028";
        ram_buffer(49538) := X"0C02BFD8";
        ram_buffer(49539) := X"00000000";
        ram_buffer(49540) := X"AFC2001C";
        ram_buffer(49541) := X"8FC5002C";
        ram_buffer(49542) := X"8FC40028";
        ram_buffer(49543) := X"0C02BE10";
        ram_buffer(49544) := X"00000000";
        ram_buffer(49545) := X"8FC2001C";
        ram_buffer(49546) := X"00000000";
        ram_buffer(49547) := X"AFC2002C";
        ram_buffer(49548) := X"8FC20030";
        ram_buffer(49549) := X"00000000";
        ram_buffer(49550) := X"00021043";
        ram_buffer(49551) := X"AFC20030";
        ram_buffer(49552) := X"8FC20030";
        ram_buffer(49553) := X"00000000";
        ram_buffer(49554) := X"10400020";
        ram_buffer(49555) := X"00000000";
        ram_buffer(49556) := X"8FC20010";
        ram_buffer(49557) := X"00000000";
        ram_buffer(49558) := X"8C420000";
        ram_buffer(49559) := X"00000000";
        ram_buffer(49560) := X"AFC20014";
        ram_buffer(49561) := X"8FC20014";
        ram_buffer(49562) := X"00000000";
        ram_buffer(49563) := X"14400012";
        ram_buffer(49564) := X"00000000";
        ram_buffer(49565) := X"8FC60010";
        ram_buffer(49566) := X"8FC50010";
        ram_buffer(49567) := X"8FC40028";
        ram_buffer(49568) := X"0C02BFD8";
        ram_buffer(49569) := X"00000000";
        ram_buffer(49570) := X"00401821";
        ram_buffer(49571) := X"8FC20010";
        ram_buffer(49572) := X"00000000";
        ram_buffer(49573) := X"AC430000";
        ram_buffer(49574) := X"8FC20010";
        ram_buffer(49575) := X"00000000";
        ram_buffer(49576) := X"8C420000";
        ram_buffer(49577) := X"00000000";
        ram_buffer(49578) := X"AFC20014";
        ram_buffer(49579) := X"8FC20014";
        ram_buffer(49580) := X"00000000";
        ram_buffer(49581) := X"AC400000";
        ram_buffer(49582) := X"8FC20014";
        ram_buffer(49583) := X"00000000";
        ram_buffer(49584) := X"AFC20010";
        ram_buffer(49585) := X"1000FFC8";
        ram_buffer(49586) := X"00000000";
        ram_buffer(49587) := X"00000000";
        ram_buffer(49588) := X"8FC2002C";
        ram_buffer(49589) := X"03C0E821";
        ram_buffer(49590) := X"8FBF0024";
        ram_buffer(49591) := X"8FBE0020";
        ram_buffer(49592) := X"27BD0028";
        ram_buffer(49593) := X"03E00008";
        ram_buffer(49594) := X"00000000";
        ram_buffer(49595) := X"27BDFFC0";
        ram_buffer(49596) := X"AFBF003C";
        ram_buffer(49597) := X"AFBE0038";
        ram_buffer(49598) := X"03A0F021";
        ram_buffer(49599) := X"AFC40040";
        ram_buffer(49600) := X"AFC50044";
        ram_buffer(49601) := X"AFC60048";
        ram_buffer(49602) := X"8FC20048";
        ram_buffer(49603) := X"00000000";
        ram_buffer(49604) := X"00021143";
        ram_buffer(49605) := X"AFC20028";
        ram_buffer(49606) := X"8FC20044";
        ram_buffer(49607) := X"00000000";
        ram_buffer(49608) := X"8C420004";
        ram_buffer(49609) := X"00000000";
        ram_buffer(49610) := X"AFC20014";
        ram_buffer(49611) := X"8FC20044";
        ram_buffer(49612) := X"00000000";
        ram_buffer(49613) := X"8C430010";
        ram_buffer(49614) := X"8FC20028";
        ram_buffer(49615) := X"00000000";
        ram_buffer(49616) := X"00621021";
        ram_buffer(49617) := X"24420001";
        ram_buffer(49618) := X"AFC20018";
        ram_buffer(49619) := X"8FC20044";
        ram_buffer(49620) := X"00000000";
        ram_buffer(49621) := X"8C420008";
        ram_buffer(49622) := X"00000000";
        ram_buffer(49623) := X"AFC20010";
        ram_buffer(49624) := X"10000009";
        ram_buffer(49625) := X"00000000";
        ram_buffer(49626) := X"8FC20014";
        ram_buffer(49627) := X"00000000";
        ram_buffer(49628) := X"24420001";
        ram_buffer(49629) := X"AFC20014";
        ram_buffer(49630) := X"8FC20010";
        ram_buffer(49631) := X"00000000";
        ram_buffer(49632) := X"00021040";
        ram_buffer(49633) := X"AFC20010";
        ram_buffer(49634) := X"8FC30018";
        ram_buffer(49635) := X"8FC20010";
        ram_buffer(49636) := X"00000000";
        ram_buffer(49637) := X"0043102A";
        ram_buffer(49638) := X"1440FFF3";
        ram_buffer(49639) := X"00000000";
        ram_buffer(49640) := X"8FC50014";
        ram_buffer(49641) := X"8FC40040";
        ram_buffer(49642) := X"0C02BDA8";
        ram_buffer(49643) := X"00000000";
        ram_buffer(49644) := X"AFC2002C";
        ram_buffer(49645) := X"8FC2002C";
        ram_buffer(49646) := X"00000000";
        ram_buffer(49647) := X"24420014";
        ram_buffer(49648) := X"AFC20020";
        ram_buffer(49649) := X"AFC00010";
        ram_buffer(49650) := X"1000000A";
        ram_buffer(49651) := X"00000000";
        ram_buffer(49652) := X"8FC20020";
        ram_buffer(49653) := X"00000000";
        ram_buffer(49654) := X"24430004";
        ram_buffer(49655) := X"AFC30020";
        ram_buffer(49656) := X"AC400000";
        ram_buffer(49657) := X"8FC20010";
        ram_buffer(49658) := X"00000000";
        ram_buffer(49659) := X"24420001";
        ram_buffer(49660) := X"AFC20010";
        ram_buffer(49661) := X"8FC30010";
        ram_buffer(49662) := X"8FC20028";
        ram_buffer(49663) := X"00000000";
        ram_buffer(49664) := X"0062102A";
        ram_buffer(49665) := X"1440FFF2";
        ram_buffer(49666) := X"00000000";
        ram_buffer(49667) := X"8FC20044";
        ram_buffer(49668) := X"00000000";
        ram_buffer(49669) := X"24420014";
        ram_buffer(49670) := X"AFC2001C";
        ram_buffer(49671) := X"8FC20044";
        ram_buffer(49672) := X"00000000";
        ram_buffer(49673) := X"8C420010";
        ram_buffer(49674) := X"00000000";
        ram_buffer(49675) := X"00021080";
        ram_buffer(49676) := X"8FC3001C";
        ram_buffer(49677) := X"00000000";
        ram_buffer(49678) := X"00621021";
        ram_buffer(49679) := X"AFC20030";
        ram_buffer(49680) := X"8FC20048";
        ram_buffer(49681) := X"00000000";
        ram_buffer(49682) := X"3042001F";
        ram_buffer(49683) := X"AFC20048";
        ram_buffer(49684) := X"8FC20048";
        ram_buffer(49685) := X"00000000";
        ram_buffer(49686) := X"10400034";
        ram_buffer(49687) := X"00000000";
        ram_buffer(49688) := X"24030020";
        ram_buffer(49689) := X"8FC20048";
        ram_buffer(49690) := X"00000000";
        ram_buffer(49691) := X"00621023";
        ram_buffer(49692) := X"AFC20014";
        ram_buffer(49693) := X"AFC00024";
        ram_buffer(49694) := X"8FC20020";
        ram_buffer(49695) := X"00000000";
        ram_buffer(49696) := X"24430004";
        ram_buffer(49697) := X"AFC30020";
        ram_buffer(49698) := X"8FC3001C";
        ram_buffer(49699) := X"00000000";
        ram_buffer(49700) := X"8C640000";
        ram_buffer(49701) := X"8FC30048";
        ram_buffer(49702) := X"00000000";
        ram_buffer(49703) := X"00642004";
        ram_buffer(49704) := X"8FC30024";
        ram_buffer(49705) := X"00000000";
        ram_buffer(49706) := X"00831825";
        ram_buffer(49707) := X"AC430000";
        ram_buffer(49708) := X"8FC2001C";
        ram_buffer(49709) := X"00000000";
        ram_buffer(49710) := X"24430004";
        ram_buffer(49711) := X"AFC3001C";
        ram_buffer(49712) := X"8C430000";
        ram_buffer(49713) := X"8FC20014";
        ram_buffer(49714) := X"00000000";
        ram_buffer(49715) := X"00431006";
        ram_buffer(49716) := X"AFC20024";
        ram_buffer(49717) := X"8FC3001C";
        ram_buffer(49718) := X"8FC20030";
        ram_buffer(49719) := X"00000000";
        ram_buffer(49720) := X"0062102B";
        ram_buffer(49721) := X"1440FFE4";
        ram_buffer(49722) := X"00000000";
        ram_buffer(49723) := X"8FC20020";
        ram_buffer(49724) := X"8FC30024";
        ram_buffer(49725) := X"00000000";
        ram_buffer(49726) := X"AC430000";
        ram_buffer(49727) := X"8FC20020";
        ram_buffer(49728) := X"00000000";
        ram_buffer(49729) := X"8C420000";
        ram_buffer(49730) := X"00000000";
        ram_buffer(49731) := X"10400018";
        ram_buffer(49732) := X"00000000";
        ram_buffer(49733) := X"8FC20018";
        ram_buffer(49734) := X"00000000";
        ram_buffer(49735) := X"24420001";
        ram_buffer(49736) := X"AFC20018";
        ram_buffer(49737) := X"10000012";
        ram_buffer(49738) := X"00000000";
        ram_buffer(49739) := X"8FC20020";
        ram_buffer(49740) := X"00000000";
        ram_buffer(49741) := X"24430004";
        ram_buffer(49742) := X"AFC30020";
        ram_buffer(49743) := X"8FC3001C";
        ram_buffer(49744) := X"00000000";
        ram_buffer(49745) := X"24640004";
        ram_buffer(49746) := X"AFC4001C";
        ram_buffer(49747) := X"8C630000";
        ram_buffer(49748) := X"00000000";
        ram_buffer(49749) := X"AC430000";
        ram_buffer(49750) := X"8FC3001C";
        ram_buffer(49751) := X"8FC20030";
        ram_buffer(49752) := X"00000000";
        ram_buffer(49753) := X"0062102B";
        ram_buffer(49754) := X"1440FFF0";
        ram_buffer(49755) := X"00000000";
        ram_buffer(49756) := X"8FC20018";
        ram_buffer(49757) := X"00000000";
        ram_buffer(49758) := X"2443FFFF";
        ram_buffer(49759) := X"8FC2002C";
        ram_buffer(49760) := X"00000000";
        ram_buffer(49761) := X"AC430010";
        ram_buffer(49762) := X"8FC50044";
        ram_buffer(49763) := X"8FC40040";
        ram_buffer(49764) := X"0C02BE10";
        ram_buffer(49765) := X"00000000";
        ram_buffer(49766) := X"8FC2002C";
        ram_buffer(49767) := X"03C0E821";
        ram_buffer(49768) := X"8FBF003C";
        ram_buffer(49769) := X"8FBE0038";
        ram_buffer(49770) := X"27BD0040";
        ram_buffer(49771) := X"03E00008";
        ram_buffer(49772) := X"00000000";
        ram_buffer(49773) := X"27BDFFE0";
        ram_buffer(49774) := X"AFBE001C";
        ram_buffer(49775) := X"03A0F021";
        ram_buffer(49776) := X"AFC40020";
        ram_buffer(49777) := X"AFC50024";
        ram_buffer(49778) := X"8FC20020";
        ram_buffer(49779) := X"00000000";
        ram_buffer(49780) := X"8C420010";
        ram_buffer(49781) := X"00000000";
        ram_buffer(49782) := X"AFC20008";
        ram_buffer(49783) := X"8FC20024";
        ram_buffer(49784) := X"00000000";
        ram_buffer(49785) := X"8C420010";
        ram_buffer(49786) := X"00000000";
        ram_buffer(49787) := X"AFC2000C";
        ram_buffer(49788) := X"8FC30008";
        ram_buffer(49789) := X"8FC2000C";
        ram_buffer(49790) := X"00000000";
        ram_buffer(49791) := X"00621023";
        ram_buffer(49792) := X"AFC20008";
        ram_buffer(49793) := X"8FC20008";
        ram_buffer(49794) := X"00000000";
        ram_buffer(49795) := X"10400004";
        ram_buffer(49796) := X"00000000";
        ram_buffer(49797) := X"8FC20008";
        ram_buffer(49798) := X"10000042";
        ram_buffer(49799) := X"00000000";
        ram_buffer(49800) := X"8FC20020";
        ram_buffer(49801) := X"00000000";
        ram_buffer(49802) := X"24420014";
        ram_buffer(49803) := X"AFC20010";
        ram_buffer(49804) := X"8FC2000C";
        ram_buffer(49805) := X"00000000";
        ram_buffer(49806) := X"00021080";
        ram_buffer(49807) := X"8FC30010";
        ram_buffer(49808) := X"00000000";
        ram_buffer(49809) := X"00621021";
        ram_buffer(49810) := X"AFC20000";
        ram_buffer(49811) := X"8FC20024";
        ram_buffer(49812) := X"00000000";
        ram_buffer(49813) := X"24420014";
        ram_buffer(49814) := X"AFC20014";
        ram_buffer(49815) := X"8FC2000C";
        ram_buffer(49816) := X"00000000";
        ram_buffer(49817) := X"00021080";
        ram_buffer(49818) := X"8FC30014";
        ram_buffer(49819) := X"00000000";
        ram_buffer(49820) := X"00621021";
        ram_buffer(49821) := X"AFC20004";
        ram_buffer(49822) := X"8FC20000";
        ram_buffer(49823) := X"00000000";
        ram_buffer(49824) := X"2442FFFC";
        ram_buffer(49825) := X"AFC20000";
        ram_buffer(49826) := X"8FC20000";
        ram_buffer(49827) := X"00000000";
        ram_buffer(49828) := X"8C430000";
        ram_buffer(49829) := X"8FC20004";
        ram_buffer(49830) := X"00000000";
        ram_buffer(49831) := X"2442FFFC";
        ram_buffer(49832) := X"AFC20004";
        ram_buffer(49833) := X"8FC20004";
        ram_buffer(49834) := X"00000000";
        ram_buffer(49835) := X"8C420000";
        ram_buffer(49836) := X"00000000";
        ram_buffer(49837) := X"10620011";
        ram_buffer(49838) := X"00000000";
        ram_buffer(49839) := X"8FC20000";
        ram_buffer(49840) := X"00000000";
        ram_buffer(49841) := X"8C430000";
        ram_buffer(49842) := X"8FC20004";
        ram_buffer(49843) := X"00000000";
        ram_buffer(49844) := X"8C420000";
        ram_buffer(49845) := X"00000000";
        ram_buffer(49846) := X"0062102B";
        ram_buffer(49847) := X"10400004";
        ram_buffer(49848) := X"00000000";
        ram_buffer(49849) := X"2402FFFF";
        ram_buffer(49850) := X"1000000E";
        ram_buffer(49851) := X"00000000";
        ram_buffer(49852) := X"24020001";
        ram_buffer(49853) := X"1000000B";
        ram_buffer(49854) := X"00000000";
        ram_buffer(49855) := X"8FC30000";
        ram_buffer(49856) := X"8FC20010";
        ram_buffer(49857) := X"00000000";
        ram_buffer(49858) := X"0043102B";
        ram_buffer(49859) := X"10400003";
        ram_buffer(49860) := X"00000000";
        ram_buffer(49861) := X"1000FFD8";
        ram_buffer(49862) := X"00000000";
        ram_buffer(49863) := X"00000000";
        ram_buffer(49864) := X"00001021";
        ram_buffer(49865) := X"03C0E821";
        ram_buffer(49866) := X"8FBE001C";
        ram_buffer(49867) := X"27BD0020";
        ram_buffer(49868) := X"03E00008";
        ram_buffer(49869) := X"00000000";
        ram_buffer(49870) := X"27BDFFB8";
        ram_buffer(49871) := X"AFBF0044";
        ram_buffer(49872) := X"AFBE0040";
        ram_buffer(49873) := X"03A0F021";
        ram_buffer(49874) := X"AFC40048";
        ram_buffer(49875) := X"AFC5004C";
        ram_buffer(49876) := X"AFC60050";
        ram_buffer(49877) := X"8FC50050";
        ram_buffer(49878) := X"8FC4004C";
        ram_buffer(49879) := X"0C02C26D";
        ram_buffer(49880) := X"00000000";
        ram_buffer(49881) := X"AFC20010";
        ram_buffer(49882) := X"8FC20010";
        ram_buffer(49883) := X"00000000";
        ram_buffer(49884) := X"1440000F";
        ram_buffer(49885) := X"00000000";
        ram_buffer(49886) := X"00002821";
        ram_buffer(49887) := X"8FC40048";
        ram_buffer(49888) := X"0C02BDA8";
        ram_buffer(49889) := X"00000000";
        ram_buffer(49890) := X"AFC20028";
        ram_buffer(49891) := X"8FC20028";
        ram_buffer(49892) := X"24030001";
        ram_buffer(49893) := X"AC430010";
        ram_buffer(49894) := X"8FC20028";
        ram_buffer(49895) := X"00000000";
        ram_buffer(49896) := X"AC400014";
        ram_buffer(49897) := X"8FC20028";
        ram_buffer(49898) := X"100000C6";
        ram_buffer(49899) := X"00000000";
        ram_buffer(49900) := X"8FC20010";
        ram_buffer(49901) := X"00000000";
        ram_buffer(49902) := X"0441000E";
        ram_buffer(49903) := X"00000000";
        ram_buffer(49904) := X"8FC2004C";
        ram_buffer(49905) := X"00000000";
        ram_buffer(49906) := X"AFC20028";
        ram_buffer(49907) := X"8FC20050";
        ram_buffer(49908) := X"00000000";
        ram_buffer(49909) := X"AFC2004C";
        ram_buffer(49910) := X"8FC20028";
        ram_buffer(49911) := X"00000000";
        ram_buffer(49912) := X"AFC20050";
        ram_buffer(49913) := X"24020001";
        ram_buffer(49914) := X"AFC20010";
        ram_buffer(49915) := X"10000002";
        ram_buffer(49916) := X"00000000";
        ram_buffer(49917) := X"AFC00010";
        ram_buffer(49918) := X"8FC2004C";
        ram_buffer(49919) := X"00000000";
        ram_buffer(49920) := X"8C420004";
        ram_buffer(49921) := X"00000000";
        ram_buffer(49922) := X"00402821";
        ram_buffer(49923) := X"8FC40048";
        ram_buffer(49924) := X"0C02BDA8";
        ram_buffer(49925) := X"00000000";
        ram_buffer(49926) := X"AFC20028";
        ram_buffer(49927) := X"8FC20028";
        ram_buffer(49928) := X"8FC30010";
        ram_buffer(49929) := X"00000000";
        ram_buffer(49930) := X"AC43000C";
        ram_buffer(49931) := X"8FC2004C";
        ram_buffer(49932) := X"00000000";
        ram_buffer(49933) := X"8C420010";
        ram_buffer(49934) := X"00000000";
        ram_buffer(49935) := X"AFC20014";
        ram_buffer(49936) := X"8FC2004C";
        ram_buffer(49937) := X"00000000";
        ram_buffer(49938) := X"24420014";
        ram_buffer(49939) := X"AFC2001C";
        ram_buffer(49940) := X"8FC20014";
        ram_buffer(49941) := X"00000000";
        ram_buffer(49942) := X"00021080";
        ram_buffer(49943) := X"8FC3001C";
        ram_buffer(49944) := X"00000000";
        ram_buffer(49945) := X"00621021";
        ram_buffer(49946) := X"AFC2002C";
        ram_buffer(49947) := X"8FC20050";
        ram_buffer(49948) := X"00000000";
        ram_buffer(49949) := X"8C420010";
        ram_buffer(49950) := X"00000000";
        ram_buffer(49951) := X"AFC20030";
        ram_buffer(49952) := X"8FC20050";
        ram_buffer(49953) := X"00000000";
        ram_buffer(49954) := X"24420014";
        ram_buffer(49955) := X"AFC20020";
        ram_buffer(49956) := X"8FC20030";
        ram_buffer(49957) := X"00000000";
        ram_buffer(49958) := X"00021080";
        ram_buffer(49959) := X"8FC30020";
        ram_buffer(49960) := X"00000000";
        ram_buffer(49961) := X"00621021";
        ram_buffer(49962) := X"AFC20034";
        ram_buffer(49963) := X"8FC20028";
        ram_buffer(49964) := X"00000000";
        ram_buffer(49965) := X"24420014";
        ram_buffer(49966) := X"AFC20024";
        ram_buffer(49967) := X"AFC00018";
        ram_buffer(49968) := X"8FC2001C";
        ram_buffer(49969) := X"00000000";
        ram_buffer(49970) := X"8C420000";
        ram_buffer(49971) := X"00000000";
        ram_buffer(49972) := X"3043FFFF";
        ram_buffer(49973) := X"8FC20020";
        ram_buffer(49974) := X"00000000";
        ram_buffer(49975) := X"8C420000";
        ram_buffer(49976) := X"00000000";
        ram_buffer(49977) := X"3042FFFF";
        ram_buffer(49978) := X"00621823";
        ram_buffer(49979) := X"8FC20018";
        ram_buffer(49980) := X"00000000";
        ram_buffer(49981) := X"00621021";
        ram_buffer(49982) := X"AFC20038";
        ram_buffer(49983) := X"8FC20038";
        ram_buffer(49984) := X"00000000";
        ram_buffer(49985) := X"00021403";
        ram_buffer(49986) := X"AFC20018";
        ram_buffer(49987) := X"8FC2001C";
        ram_buffer(49988) := X"00000000";
        ram_buffer(49989) := X"24430004";
        ram_buffer(49990) := X"AFC3001C";
        ram_buffer(49991) := X"8C420000";
        ram_buffer(49992) := X"00000000";
        ram_buffer(49993) := X"00021C02";
        ram_buffer(49994) := X"8FC20020";
        ram_buffer(49995) := X"00000000";
        ram_buffer(49996) := X"24440004";
        ram_buffer(49997) := X"AFC40020";
        ram_buffer(49998) := X"8C420000";
        ram_buffer(49999) := X"00000000";
        ram_buffer(50000) := X"00021402";
        ram_buffer(50001) := X"00621823";
        ram_buffer(50002) := X"8FC20018";
        ram_buffer(50003) := X"00000000";
        ram_buffer(50004) := X"00621021";
        ram_buffer(50005) := X"AFC2003C";
        ram_buffer(50006) := X"8FC2003C";
        ram_buffer(50007) := X"00000000";
        ram_buffer(50008) := X"00021403";
        ram_buffer(50009) := X"AFC20018";
        ram_buffer(50010) := X"8FC20024";
        ram_buffer(50011) := X"00000000";
        ram_buffer(50012) := X"24430004";
        ram_buffer(50013) := X"AFC30024";
        ram_buffer(50014) := X"8FC3003C";
        ram_buffer(50015) := X"00000000";
        ram_buffer(50016) := X"00032400";
        ram_buffer(50017) := X"8FC30038";
        ram_buffer(50018) := X"00000000";
        ram_buffer(50019) := X"3063FFFF";
        ram_buffer(50020) := X"00831825";
        ram_buffer(50021) := X"AC430000";
        ram_buffer(50022) := X"8FC30020";
        ram_buffer(50023) := X"8FC20034";
        ram_buffer(50024) := X"00000000";
        ram_buffer(50025) := X"0062102B";
        ram_buffer(50026) := X"1440FFC5";
        ram_buffer(50027) := X"00000000";
        ram_buffer(50028) := X"10000029";
        ram_buffer(50029) := X"00000000";
        ram_buffer(50030) := X"8FC2001C";
        ram_buffer(50031) := X"00000000";
        ram_buffer(50032) := X"8C420000";
        ram_buffer(50033) := X"00000000";
        ram_buffer(50034) := X"3043FFFF";
        ram_buffer(50035) := X"8FC20018";
        ram_buffer(50036) := X"00000000";
        ram_buffer(50037) := X"00621021";
        ram_buffer(50038) := X"AFC20038";
        ram_buffer(50039) := X"8FC20038";
        ram_buffer(50040) := X"00000000";
        ram_buffer(50041) := X"00021403";
        ram_buffer(50042) := X"AFC20018";
        ram_buffer(50043) := X"8FC2001C";
        ram_buffer(50044) := X"00000000";
        ram_buffer(50045) := X"24430004";
        ram_buffer(50046) := X"AFC3001C";
        ram_buffer(50047) := X"8C420000";
        ram_buffer(50048) := X"00000000";
        ram_buffer(50049) := X"00021C02";
        ram_buffer(50050) := X"8FC20018";
        ram_buffer(50051) := X"00000000";
        ram_buffer(50052) := X"00621021";
        ram_buffer(50053) := X"AFC2003C";
        ram_buffer(50054) := X"8FC2003C";
        ram_buffer(50055) := X"00000000";
        ram_buffer(50056) := X"00021403";
        ram_buffer(50057) := X"AFC20018";
        ram_buffer(50058) := X"8FC20024";
        ram_buffer(50059) := X"00000000";
        ram_buffer(50060) := X"24430004";
        ram_buffer(50061) := X"AFC30024";
        ram_buffer(50062) := X"8FC3003C";
        ram_buffer(50063) := X"00000000";
        ram_buffer(50064) := X"00032400";
        ram_buffer(50065) := X"8FC30038";
        ram_buffer(50066) := X"00000000";
        ram_buffer(50067) := X"3063FFFF";
        ram_buffer(50068) := X"00831825";
        ram_buffer(50069) := X"AC430000";
        ram_buffer(50070) := X"8FC3001C";
        ram_buffer(50071) := X"8FC2002C";
        ram_buffer(50072) := X"00000000";
        ram_buffer(50073) := X"0062102B";
        ram_buffer(50074) := X"1440FFD3";
        ram_buffer(50075) := X"00000000";
        ram_buffer(50076) := X"10000005";
        ram_buffer(50077) := X"00000000";
        ram_buffer(50078) := X"8FC20014";
        ram_buffer(50079) := X"00000000";
        ram_buffer(50080) := X"2442FFFF";
        ram_buffer(50081) := X"AFC20014";
        ram_buffer(50082) := X"8FC20024";
        ram_buffer(50083) := X"00000000";
        ram_buffer(50084) := X"2442FFFC";
        ram_buffer(50085) := X"AFC20024";
        ram_buffer(50086) := X"8FC20024";
        ram_buffer(50087) := X"00000000";
        ram_buffer(50088) := X"8C420000";
        ram_buffer(50089) := X"00000000";
        ram_buffer(50090) := X"1040FFF3";
        ram_buffer(50091) := X"00000000";
        ram_buffer(50092) := X"8FC20028";
        ram_buffer(50093) := X"8FC30014";
        ram_buffer(50094) := X"00000000";
        ram_buffer(50095) := X"AC430010";
        ram_buffer(50096) := X"8FC20028";
        ram_buffer(50097) := X"03C0E821";
        ram_buffer(50098) := X"8FBF0044";
        ram_buffer(50099) := X"8FBE0040";
        ram_buffer(50100) := X"27BD0048";
        ram_buffer(50101) := X"03E00008";
        ram_buffer(50102) := X"00000000";
        ram_buffer(50103) := X"27BDFFE8";
        ram_buffer(50104) := X"AFBE0014";
        ram_buffer(50105) := X"AFB00010";
        ram_buffer(50106) := X"03A0F021";
        ram_buffer(50107) := X"AFC5001C";
        ram_buffer(50108) := X"AFC40018";
        ram_buffer(50109) := X"8FC3001C";
        ram_buffer(50110) := X"8FC20018";
        ram_buffer(50111) := X"AFC30004";
        ram_buffer(50112) := X"AFC20000";
        ram_buffer(50113) := X"8FC30000";
        ram_buffer(50114) := X"3C027FF0";
        ram_buffer(50115) := X"00621824";
        ram_buffer(50116) := X"3C02FCC0";
        ram_buffer(50117) := X"00621021";
        ram_buffer(50118) := X"00408021";
        ram_buffer(50119) := X"1A000006";
        ram_buffer(50120) := X"00000000";
        ram_buffer(50121) := X"02001021";
        ram_buffer(50122) := X"AFC20008";
        ram_buffer(50123) := X"AFC0000C";
        ram_buffer(50124) := X"10000019";
        ram_buffer(50125) := X"00000000";
        ram_buffer(50126) := X"00101023";
        ram_buffer(50127) := X"00028503";
        ram_buffer(50128) := X"2A020014";
        ram_buffer(50129) := X"10400007";
        ram_buffer(50130) := X"00000000";
        ram_buffer(50131) := X"3C020008";
        ram_buffer(50132) := X"02021007";
        ram_buffer(50133) := X"AFC20008";
        ram_buffer(50134) := X"AFC0000C";
        ram_buffer(50135) := X"1000000E";
        ram_buffer(50136) := X"00000000";
        ram_buffer(50137) := X"AFC00008";
        ram_buffer(50138) := X"2610FFEC";
        ram_buffer(50139) := X"2A02001F";
        ram_buffer(50140) := X"10400007";
        ram_buffer(50141) := X"00000000";
        ram_buffer(50142) := X"2402001F";
        ram_buffer(50143) := X"00501023";
        ram_buffer(50144) := X"24030001";
        ram_buffer(50145) := X"00431004";
        ram_buffer(50146) := X"10000002";
        ram_buffer(50147) := X"00000000";
        ram_buffer(50148) := X"24020001";
        ram_buffer(50149) := X"AFC2000C";
        ram_buffer(50150) := X"8FC3000C";
        ram_buffer(50151) := X"8FC20008";
        ram_buffer(50152) := X"03C0E821";
        ram_buffer(50153) := X"8FBE0014";
        ram_buffer(50154) := X"8FB00010";
        ram_buffer(50155) := X"27BD0018";
        ram_buffer(50156) := X"03E00008";
        ram_buffer(50157) := X"00000000";
        ram_buffer(50158) := X"27BDFFC8";
        ram_buffer(50159) := X"AFBF0034";
        ram_buffer(50160) := X"AFBE0030";
        ram_buffer(50161) := X"03A0F021";
        ram_buffer(50162) := X"AFC40038";
        ram_buffer(50163) := X"AFC5003C";
        ram_buffer(50164) := X"8FC20038";
        ram_buffer(50165) := X"00000000";
        ram_buffer(50166) := X"24420014";
        ram_buffer(50167) := X"AFC20014";
        ram_buffer(50168) := X"8FC20038";
        ram_buffer(50169) := X"00000000";
        ram_buffer(50170) := X"8C420010";
        ram_buffer(50171) := X"00000000";
        ram_buffer(50172) := X"00021080";
        ram_buffer(50173) := X"8FC30014";
        ram_buffer(50174) := X"00000000";
        ram_buffer(50175) := X"00621021";
        ram_buffer(50176) := X"AFC20010";
        ram_buffer(50177) := X"8FC20010";
        ram_buffer(50178) := X"00000000";
        ram_buffer(50179) := X"2442FFFC";
        ram_buffer(50180) := X"AFC20010";
        ram_buffer(50181) := X"8FC20010";
        ram_buffer(50182) := X"00000000";
        ram_buffer(50183) := X"8C420000";
        ram_buffer(50184) := X"00000000";
        ram_buffer(50185) := X"AFC20018";
        ram_buffer(50186) := X"8FC40018";
        ram_buffer(50187) := X"0C02BF41";
        ram_buffer(50188) := X"00000000";
        ram_buffer(50189) := X"AFC2001C";
        ram_buffer(50190) := X"24030020";
        ram_buffer(50191) := X"8FC2001C";
        ram_buffer(50192) := X"00000000";
        ram_buffer(50193) := X"00621823";
        ram_buffer(50194) := X"8FC2003C";
        ram_buffer(50195) := X"00000000";
        ram_buffer(50196) := X"AC430000";
        ram_buffer(50197) := X"8FC2001C";
        ram_buffer(50198) := X"00000000";
        ram_buffer(50199) := X"2842000B";
        ram_buffer(50200) := X"1040002D";
        ram_buffer(50201) := X"00000000";
        ram_buffer(50202) := X"2403000B";
        ram_buffer(50203) := X"8FC2001C";
        ram_buffer(50204) := X"00000000";
        ram_buffer(50205) := X"00621023";
        ram_buffer(50206) := X"8FC30018";
        ram_buffer(50207) := X"00000000";
        ram_buffer(50208) := X"00431806";
        ram_buffer(50209) := X"3C023FF0";
        ram_buffer(50210) := X"00621025";
        ram_buffer(50211) := X"AFC20028";
        ram_buffer(50212) := X"8FC30010";
        ram_buffer(50213) := X"8FC20014";
        ram_buffer(50214) := X"00000000";
        ram_buffer(50215) := X"0043102B";
        ram_buffer(50216) := X"1040000A";
        ram_buffer(50217) := X"00000000";
        ram_buffer(50218) := X"8FC20010";
        ram_buffer(50219) := X"00000000";
        ram_buffer(50220) := X"2442FFFC";
        ram_buffer(50221) := X"AFC20010";
        ram_buffer(50222) := X"8FC20010";
        ram_buffer(50223) := X"00000000";
        ram_buffer(50224) := X"8C420000";
        ram_buffer(50225) := X"10000002";
        ram_buffer(50226) := X"00000000";
        ram_buffer(50227) := X"00001021";
        ram_buffer(50228) := X"AFC20020";
        ram_buffer(50229) := X"8FC2001C";
        ram_buffer(50230) := X"00000000";
        ram_buffer(50231) := X"24420015";
        ram_buffer(50232) := X"8FC30018";
        ram_buffer(50233) := X"00000000";
        ram_buffer(50234) := X"00431804";
        ram_buffer(50235) := X"2404000B";
        ram_buffer(50236) := X"8FC2001C";
        ram_buffer(50237) := X"00000000";
        ram_buffer(50238) := X"00821023";
        ram_buffer(50239) := X"8FC40020";
        ram_buffer(50240) := X"00000000";
        ram_buffer(50241) := X"00441006";
        ram_buffer(50242) := X"00621025";
        ram_buffer(50243) := X"AFC2002C";
        ram_buffer(50244) := X"10000050";
        ram_buffer(50245) := X"00000000";
        ram_buffer(50246) := X"8FC30010";
        ram_buffer(50247) := X"8FC20014";
        ram_buffer(50248) := X"00000000";
        ram_buffer(50249) := X"0043102B";
        ram_buffer(50250) := X"1040000A";
        ram_buffer(50251) := X"00000000";
        ram_buffer(50252) := X"8FC20010";
        ram_buffer(50253) := X"00000000";
        ram_buffer(50254) := X"2442FFFC";
        ram_buffer(50255) := X"AFC20010";
        ram_buffer(50256) := X"8FC20010";
        ram_buffer(50257) := X"00000000";
        ram_buffer(50258) := X"8C420000";
        ram_buffer(50259) := X"10000002";
        ram_buffer(50260) := X"00000000";
        ram_buffer(50261) := X"00001021";
        ram_buffer(50262) := X"AFC20024";
        ram_buffer(50263) := X"8FC2001C";
        ram_buffer(50264) := X"00000000";
        ram_buffer(50265) := X"2442FFF5";
        ram_buffer(50266) := X"AFC2001C";
        ram_buffer(50267) := X"8FC2001C";
        ram_buffer(50268) := X"00000000";
        ram_buffer(50269) := X"10400030";
        ram_buffer(50270) := X"00000000";
        ram_buffer(50271) := X"8FC30018";
        ram_buffer(50272) := X"8FC2001C";
        ram_buffer(50273) := X"00000000";
        ram_buffer(50274) := X"00431804";
        ram_buffer(50275) := X"24040020";
        ram_buffer(50276) := X"8FC2001C";
        ram_buffer(50277) := X"00000000";
        ram_buffer(50278) := X"00821023";
        ram_buffer(50279) := X"8FC40024";
        ram_buffer(50280) := X"00000000";
        ram_buffer(50281) := X"00441006";
        ram_buffer(50282) := X"00621825";
        ram_buffer(50283) := X"3C023FF0";
        ram_buffer(50284) := X"00621025";
        ram_buffer(50285) := X"AFC20028";
        ram_buffer(50286) := X"8FC30010";
        ram_buffer(50287) := X"8FC20014";
        ram_buffer(50288) := X"00000000";
        ram_buffer(50289) := X"0043102B";
        ram_buffer(50290) := X"1040000A";
        ram_buffer(50291) := X"00000000";
        ram_buffer(50292) := X"8FC20010";
        ram_buffer(50293) := X"00000000";
        ram_buffer(50294) := X"2442FFFC";
        ram_buffer(50295) := X"AFC20010";
        ram_buffer(50296) := X"8FC20010";
        ram_buffer(50297) := X"00000000";
        ram_buffer(50298) := X"8C420000";
        ram_buffer(50299) := X"10000002";
        ram_buffer(50300) := X"00000000";
        ram_buffer(50301) := X"00001021";
        ram_buffer(50302) := X"AFC20018";
        ram_buffer(50303) := X"8FC30024";
        ram_buffer(50304) := X"8FC2001C";
        ram_buffer(50305) := X"00000000";
        ram_buffer(50306) := X"00431804";
        ram_buffer(50307) := X"24040020";
        ram_buffer(50308) := X"8FC2001C";
        ram_buffer(50309) := X"00000000";
        ram_buffer(50310) := X"00821023";
        ram_buffer(50311) := X"8FC40018";
        ram_buffer(50312) := X"00000000";
        ram_buffer(50313) := X"00441006";
        ram_buffer(50314) := X"00621025";
        ram_buffer(50315) := X"AFC2002C";
        ram_buffer(50316) := X"10000008";
        ram_buffer(50317) := X"00000000";
        ram_buffer(50318) := X"8FC30018";
        ram_buffer(50319) := X"3C023FF0";
        ram_buffer(50320) := X"00621025";
        ram_buffer(50321) := X"AFC20028";
        ram_buffer(50322) := X"8FC20024";
        ram_buffer(50323) := X"00000000";
        ram_buffer(50324) := X"AFC2002C";
        ram_buffer(50325) := X"8FC3002C";
        ram_buffer(50326) := X"8FC20028";
        ram_buffer(50327) := X"03C0E821";
        ram_buffer(50328) := X"8FBF0034";
        ram_buffer(50329) := X"8FBE0030";
        ram_buffer(50330) := X"27BD0038";
        ram_buffer(50331) := X"03E00008";
        ram_buffer(50332) := X"00000000";
        ram_buffer(50333) := X"27BDFFB8";
        ram_buffer(50334) := X"AFBF0044";
        ram_buffer(50335) := X"AFBE0040";
        ram_buffer(50336) := X"AFB0003C";
        ram_buffer(50337) := X"03A0F021";
        ram_buffer(50338) := X"AFC40048";
        ram_buffer(50339) := X"AFC70054";
        ram_buffer(50340) := X"AFC60050";
        ram_buffer(50341) := X"8FC30054";
        ram_buffer(50342) := X"8FC20050";
        ram_buffer(50343) := X"AFC3002C";
        ram_buffer(50344) := X"AFC20028";
        ram_buffer(50345) := X"8FC30054";
        ram_buffer(50346) := X"8FC20050";
        ram_buffer(50347) := X"AFC3002C";
        ram_buffer(50348) := X"AFC20028";
        ram_buffer(50349) := X"24050001";
        ram_buffer(50350) := X"8FC40048";
        ram_buffer(50351) := X"0C02BDA8";
        ram_buffer(50352) := X"00000000";
        ram_buffer(50353) := X"AFC20018";
        ram_buffer(50354) := X"8FC20018";
        ram_buffer(50355) := X"00000000";
        ram_buffer(50356) := X"24420014";
        ram_buffer(50357) := X"AFC2001C";
        ram_buffer(50358) := X"8FC30028";
        ram_buffer(50359) := X"3C02000F";
        ram_buffer(50360) := X"3442FFFF";
        ram_buffer(50361) := X"00621024";
        ram_buffer(50362) := X"AFC20034";
        ram_buffer(50363) := X"8FC30028";
        ram_buffer(50364) := X"3C027FFF";
        ram_buffer(50365) := X"3442FFFF";
        ram_buffer(50366) := X"00621024";
        ram_buffer(50367) := X"AFC20028";
        ram_buffer(50368) := X"8FC20028";
        ram_buffer(50369) := X"00000000";
        ram_buffer(50370) := X"00021502";
        ram_buffer(50371) := X"AFC20020";
        ram_buffer(50372) := X"8FC20020";
        ram_buffer(50373) := X"00000000";
        ram_buffer(50374) := X"10400005";
        ram_buffer(50375) := X"00000000";
        ram_buffer(50376) := X"8FC30034";
        ram_buffer(50377) := X"3C020010";
        ram_buffer(50378) := X"00621025";
        ram_buffer(50379) := X"AFC20034";
        ram_buffer(50380) := X"8FC2002C";
        ram_buffer(50381) := X"00000000";
        ram_buffer(50382) := X"1040003C";
        ram_buffer(50383) := X"00000000";
        ram_buffer(50384) := X"8FC2002C";
        ram_buffer(50385) := X"00000000";
        ram_buffer(50386) := X"AFC20030";
        ram_buffer(50387) := X"27C20030";
        ram_buffer(50388) := X"00402021";
        ram_buffer(50389) := X"0C02BF71";
        ram_buffer(50390) := X"00000000";
        ram_buffer(50391) := X"AFC20014";
        ram_buffer(50392) := X"8FC20014";
        ram_buffer(50393) := X"00000000";
        ram_buffer(50394) := X"10400014";
        ram_buffer(50395) := X"00000000";
        ram_buffer(50396) := X"8FC30034";
        ram_buffer(50397) := X"24040020";
        ram_buffer(50398) := X"8FC20014";
        ram_buffer(50399) := X"00000000";
        ram_buffer(50400) := X"00821023";
        ram_buffer(50401) := X"00431804";
        ram_buffer(50402) := X"8FC20030";
        ram_buffer(50403) := X"00000000";
        ram_buffer(50404) := X"00621825";
        ram_buffer(50405) := X"8FC2001C";
        ram_buffer(50406) := X"00000000";
        ram_buffer(50407) := X"AC430000";
        ram_buffer(50408) := X"8FC30034";
        ram_buffer(50409) := X"8FC20014";
        ram_buffer(50410) := X"00000000";
        ram_buffer(50411) := X"00431006";
        ram_buffer(50412) := X"AFC20034";
        ram_buffer(50413) := X"10000005";
        ram_buffer(50414) := X"00000000";
        ram_buffer(50415) := X"8FC30030";
        ram_buffer(50416) := X"8FC2001C";
        ram_buffer(50417) := X"00000000";
        ram_buffer(50418) := X"AC430000";
        ram_buffer(50419) := X"8FC2001C";
        ram_buffer(50420) := X"00000000";
        ram_buffer(50421) := X"24420004";
        ram_buffer(50422) := X"8FC30034";
        ram_buffer(50423) := X"00000000";
        ram_buffer(50424) := X"AC430000";
        ram_buffer(50425) := X"8C420000";
        ram_buffer(50426) := X"00000000";
        ram_buffer(50427) := X"10400004";
        ram_buffer(50428) := X"00000000";
        ram_buffer(50429) := X"24020002";
        ram_buffer(50430) := X"10000002";
        ram_buffer(50431) := X"00000000";
        ram_buffer(50432) := X"24020001";
        ram_buffer(50433) := X"8FC30018";
        ram_buffer(50434) := X"00000000";
        ram_buffer(50435) := X"AC620010";
        ram_buffer(50436) := X"8FC20018";
        ram_buffer(50437) := X"00000000";
        ram_buffer(50438) := X"8C420010";
        ram_buffer(50439) := X"00000000";
        ram_buffer(50440) := X"AFC20010";
        ram_buffer(50441) := X"10000016";
        ram_buffer(50442) := X"00000000";
        ram_buffer(50443) := X"27C20034";
        ram_buffer(50444) := X"00402021";
        ram_buffer(50445) := X"0C02BF71";
        ram_buffer(50446) := X"00000000";
        ram_buffer(50447) := X"AFC20014";
        ram_buffer(50448) := X"8FC30034";
        ram_buffer(50449) := X"8FC2001C";
        ram_buffer(50450) := X"00000000";
        ram_buffer(50451) := X"AC430000";
        ram_buffer(50452) := X"8FC20018";
        ram_buffer(50453) := X"24030001";
        ram_buffer(50454) := X"AC430010";
        ram_buffer(50455) := X"8FC20018";
        ram_buffer(50456) := X"00000000";
        ram_buffer(50457) := X"8C420010";
        ram_buffer(50458) := X"00000000";
        ram_buffer(50459) := X"AFC20010";
        ram_buffer(50460) := X"8FC20014";
        ram_buffer(50461) := X"00000000";
        ram_buffer(50462) := X"24420020";
        ram_buffer(50463) := X"AFC20014";
        ram_buffer(50464) := X"8FC20020";
        ram_buffer(50465) := X"00000000";
        ram_buffer(50466) := X"10400013";
        ram_buffer(50467) := X"00000000";
        ram_buffer(50468) := X"8FC20020";
        ram_buffer(50469) := X"00000000";
        ram_buffer(50470) := X"2443FBCD";
        ram_buffer(50471) := X"8FC20014";
        ram_buffer(50472) := X"00000000";
        ram_buffer(50473) := X"00621821";
        ram_buffer(50474) := X"8FC20058";
        ram_buffer(50475) := X"00000000";
        ram_buffer(50476) := X"AC430000";
        ram_buffer(50477) := X"24030035";
        ram_buffer(50478) := X"8FC20014";
        ram_buffer(50479) := X"00000000";
        ram_buffer(50480) := X"00621823";
        ram_buffer(50481) := X"8FC2005C";
        ram_buffer(50482) := X"00000000";
        ram_buffer(50483) := X"AC430000";
        ram_buffer(50484) := X"1000001E";
        ram_buffer(50485) := X"00000000";
        ram_buffer(50486) := X"8FC20020";
        ram_buffer(50487) := X"00000000";
        ram_buffer(50488) := X"2443FBCE";
        ram_buffer(50489) := X"8FC20014";
        ram_buffer(50490) := X"00000000";
        ram_buffer(50491) := X"00621821";
        ram_buffer(50492) := X"8FC20058";
        ram_buffer(50493) := X"00000000";
        ram_buffer(50494) := X"AC430000";
        ram_buffer(50495) := X"8FC20010";
        ram_buffer(50496) := X"00000000";
        ram_buffer(50497) := X"00028140";
        ram_buffer(50498) := X"8FC30010";
        ram_buffer(50499) := X"3C023FFF";
        ram_buffer(50500) := X"3442FFFF";
        ram_buffer(50501) := X"00621021";
        ram_buffer(50502) := X"00021080";
        ram_buffer(50503) := X"8FC3001C";
        ram_buffer(50504) := X"00000000";
        ram_buffer(50505) := X"00621021";
        ram_buffer(50506) := X"8C420000";
        ram_buffer(50507) := X"00000000";
        ram_buffer(50508) := X"00402021";
        ram_buffer(50509) := X"0C02BF41";
        ram_buffer(50510) := X"00000000";
        ram_buffer(50511) := X"02021823";
        ram_buffer(50512) := X"8FC2005C";
        ram_buffer(50513) := X"00000000";
        ram_buffer(50514) := X"AC430000";
        ram_buffer(50515) := X"8FC20018";
        ram_buffer(50516) := X"03C0E821";
        ram_buffer(50517) := X"8FBF0044";
        ram_buffer(50518) := X"8FBE0040";
        ram_buffer(50519) := X"8FB0003C";
        ram_buffer(50520) := X"27BD0048";
        ram_buffer(50521) := X"03E00008";
        ram_buffer(50522) := X"00000000";
        ram_buffer(50523) := X"27BDFFC8";
        ram_buffer(50524) := X"AFBF0034";
        ram_buffer(50525) := X"AFBE0030";
        ram_buffer(50526) := X"03A0F021";
        ram_buffer(50527) := X"AFC40038";
        ram_buffer(50528) := X"AFC5003C";
        ram_buffer(50529) := X"27C20028";
        ram_buffer(50530) := X"00402821";
        ram_buffer(50531) := X"8FC40038";
        ram_buffer(50532) := X"0C02C3EE";
        ram_buffer(50533) := X"00000000";
        ram_buffer(50534) := X"AFC3001C";
        ram_buffer(50535) := X"AFC20018";
        ram_buffer(50536) := X"27C2002C";
        ram_buffer(50537) := X"00402821";
        ram_buffer(50538) := X"8FC4003C";
        ram_buffer(50539) := X"0C02C3EE";
        ram_buffer(50540) := X"00000000";
        ram_buffer(50541) := X"AFC30024";
        ram_buffer(50542) := X"AFC20020";
        ram_buffer(50543) := X"8FC30028";
        ram_buffer(50544) := X"8FC2002C";
        ram_buffer(50545) := X"00000000";
        ram_buffer(50546) := X"00621823";
        ram_buffer(50547) := X"8FC20038";
        ram_buffer(50548) := X"00000000";
        ram_buffer(50549) := X"8C440010";
        ram_buffer(50550) := X"8FC2003C";
        ram_buffer(50551) := X"00000000";
        ram_buffer(50552) := X"8C420010";
        ram_buffer(50553) := X"00000000";
        ram_buffer(50554) := X"00821023";
        ram_buffer(50555) := X"00021140";
        ram_buffer(50556) := X"00621021";
        ram_buffer(50557) := X"AFC20010";
        ram_buffer(50558) := X"8FC20010";
        ram_buffer(50559) := X"00000000";
        ram_buffer(50560) := X"18400009";
        ram_buffer(50561) := X"00000000";
        ram_buffer(50562) := X"8FC30018";
        ram_buffer(50563) := X"8FC20010";
        ram_buffer(50564) := X"00000000";
        ram_buffer(50565) := X"00021500";
        ram_buffer(50566) := X"00621021";
        ram_buffer(50567) := X"AFC20018";
        ram_buffer(50568) := X"1000000B";
        ram_buffer(50569) := X"00000000";
        ram_buffer(50570) := X"8FC20010";
        ram_buffer(50571) := X"00000000";
        ram_buffer(50572) := X"00021023";
        ram_buffer(50573) := X"AFC20010";
        ram_buffer(50574) := X"8FC30020";
        ram_buffer(50575) := X"8FC20010";
        ram_buffer(50576) := X"00000000";
        ram_buffer(50577) := X"00021500";
        ram_buffer(50578) := X"00621021";
        ram_buffer(50579) := X"AFC20020";
        ram_buffer(50580) := X"8FC3001C";
        ram_buffer(50581) := X"8FC20018";
        ram_buffer(50582) := X"8FC50024";
        ram_buffer(50583) := X"8FC40020";
        ram_buffer(50584) := X"00A03821";
        ram_buffer(50585) := X"00803021";
        ram_buffer(50586) := X"00602821";
        ram_buffer(50587) := X"00402021";
        ram_buffer(50588) := X"0C03144F";
        ram_buffer(50589) := X"00000000";
        ram_buffer(50590) := X"03C0E821";
        ram_buffer(50591) := X"8FBF0034";
        ram_buffer(50592) := X"8FBE0030";
        ram_buffer(50593) := X"27BD0038";
        ram_buffer(50594) := X"03E00008";
        ram_buffer(50595) := X"00000000";
        ram_buffer(50596) := X"27BDFFE0";
        ram_buffer(50597) := X"AFBF001C";
        ram_buffer(50598) := X"AFBE0018";
        ram_buffer(50599) := X"03A0F021";
        ram_buffer(50600) := X"AFC40020";
        ram_buffer(50601) := X"8F838134";
        ram_buffer(50602) := X"8F828130";
        ram_buffer(50603) := X"AFC30014";
        ram_buffer(50604) := X"AFC20010";
        ram_buffer(50605) := X"8FC20020";
        ram_buffer(50606) := X"00000000";
        ram_buffer(50607) := X"28420018";
        ram_buffer(50608) := X"10400017";
        ram_buffer(50609) := X"00000000";
        ram_buffer(50610) := X"3C02100D";
        ram_buffer(50611) := X"8FC30020";
        ram_buffer(50612) := X"00000000";
        ram_buffer(50613) := X"000318C0";
        ram_buffer(50614) := X"2442A938";
        ram_buffer(50615) := X"00621021";
        ram_buffer(50616) := X"8C430004";
        ram_buffer(50617) := X"8C420000";
        ram_buffer(50618) := X"10000013";
        ram_buffer(50619) := X"00000000";
        ram_buffer(50620) := X"8F87813C";
        ram_buffer(50621) := X"8F868138";
        ram_buffer(50622) := X"8FC50014";
        ram_buffer(50623) := X"8FC40010";
        ram_buffer(50624) := X"0C03174A";
        ram_buffer(50625) := X"00000000";
        ram_buffer(50626) := X"AFC30014";
        ram_buffer(50627) := X"AFC20010";
        ram_buffer(50628) := X"8FC20020";
        ram_buffer(50629) := X"00000000";
        ram_buffer(50630) := X"2442FFFF";
        ram_buffer(50631) := X"AFC20020";
        ram_buffer(50632) := X"8FC20020";
        ram_buffer(50633) := X"00000000";
        ram_buffer(50634) := X"1C40FFF1";
        ram_buffer(50635) := X"00000000";
        ram_buffer(50636) := X"8FC30014";
        ram_buffer(50637) := X"8FC20010";
        ram_buffer(50638) := X"03C0E821";
        ram_buffer(50639) := X"8FBF001C";
        ram_buffer(50640) := X"8FBE0018";
        ram_buffer(50641) := X"27BD0020";
        ram_buffer(50642) := X"03E00008";
        ram_buffer(50643) := X"00000000";
        ram_buffer(50644) := X"27BDFFE8";
        ram_buffer(50645) := X"AFBE0014";
        ram_buffer(50646) := X"03A0F021";
        ram_buffer(50647) := X"AFC40018";
        ram_buffer(50648) := X"AFC5001C";
        ram_buffer(50649) := X"AFC60020";
        ram_buffer(50650) := X"8FC2001C";
        ram_buffer(50651) := X"00000000";
        ram_buffer(50652) := X"2442FFFF";
        ram_buffer(50653) := X"00021143";
        ram_buffer(50654) := X"24420001";
        ram_buffer(50655) := X"00021080";
        ram_buffer(50656) := X"8FC30018";
        ram_buffer(50657) := X"00000000";
        ram_buffer(50658) := X"00621021";
        ram_buffer(50659) := X"AFC20004";
        ram_buffer(50660) := X"8FC20020";
        ram_buffer(50661) := X"00000000";
        ram_buffer(50662) := X"24420014";
        ram_buffer(50663) := X"AFC20000";
        ram_buffer(50664) := X"8FC20020";
        ram_buffer(50665) := X"00000000";
        ram_buffer(50666) := X"8C420010";
        ram_buffer(50667) := X"00000000";
        ram_buffer(50668) := X"00021080";
        ram_buffer(50669) := X"8FC30000";
        ram_buffer(50670) := X"00000000";
        ram_buffer(50671) := X"00621021";
        ram_buffer(50672) := X"AFC20008";
        ram_buffer(50673) := X"1000000C";
        ram_buffer(50674) := X"00000000";
        ram_buffer(50675) := X"8FC20018";
        ram_buffer(50676) := X"00000000";
        ram_buffer(50677) := X"24430004";
        ram_buffer(50678) := X"AFC30018";
        ram_buffer(50679) := X"8FC30000";
        ram_buffer(50680) := X"00000000";
        ram_buffer(50681) := X"24640004";
        ram_buffer(50682) := X"AFC40000";
        ram_buffer(50683) := X"8C630000";
        ram_buffer(50684) := X"00000000";
        ram_buffer(50685) := X"AC430000";
        ram_buffer(50686) := X"8FC30000";
        ram_buffer(50687) := X"8FC20008";
        ram_buffer(50688) := X"00000000";
        ram_buffer(50689) := X"0062102B";
        ram_buffer(50690) := X"1440FFF0";
        ram_buffer(50691) := X"00000000";
        ram_buffer(50692) := X"10000006";
        ram_buffer(50693) := X"00000000";
        ram_buffer(50694) := X"8FC20018";
        ram_buffer(50695) := X"00000000";
        ram_buffer(50696) := X"24430004";
        ram_buffer(50697) := X"AFC30018";
        ram_buffer(50698) := X"AC400000";
        ram_buffer(50699) := X"8FC30018";
        ram_buffer(50700) := X"8FC20004";
        ram_buffer(50701) := X"00000000";
        ram_buffer(50702) := X"0062102B";
        ram_buffer(50703) := X"1440FFF6";
        ram_buffer(50704) := X"00000000";
        ram_buffer(50705) := X"00000000";
        ram_buffer(50706) := X"03C0E821";
        ram_buffer(50707) := X"8FBE0014";
        ram_buffer(50708) := X"27BD0018";
        ram_buffer(50709) := X"03E00008";
        ram_buffer(50710) := X"00000000";
        ram_buffer(50711) := X"27BDFFE0";
        ram_buffer(50712) := X"AFBE001C";
        ram_buffer(50713) := X"03A0F021";
        ram_buffer(50714) := X"AFC40020";
        ram_buffer(50715) := X"AFC50024";
        ram_buffer(50716) := X"8FC20020";
        ram_buffer(50717) := X"00000000";
        ram_buffer(50718) := X"24420014";
        ram_buffer(50719) := X"AFC20004";
        ram_buffer(50720) := X"8FC20020";
        ram_buffer(50721) := X"00000000";
        ram_buffer(50722) := X"8C420010";
        ram_buffer(50723) := X"00000000";
        ram_buffer(50724) := X"AFC20008";
        ram_buffer(50725) := X"8FC20024";
        ram_buffer(50726) := X"00000000";
        ram_buffer(50727) := X"00021143";
        ram_buffer(50728) := X"AFC20000";
        ram_buffer(50729) := X"8FC30000";
        ram_buffer(50730) := X"8FC20008";
        ram_buffer(50731) := X"00000000";
        ram_buffer(50732) := X"0043102A";
        ram_buffer(50733) := X"10400006";
        ram_buffer(50734) := X"00000000";
        ram_buffer(50735) := X"8FC20008";
        ram_buffer(50736) := X"00000000";
        ram_buffer(50737) := X"AFC20000";
        ram_buffer(50738) := X"1000002D";
        ram_buffer(50739) := X"00000000";
        ram_buffer(50740) := X"8FC30000";
        ram_buffer(50741) := X"8FC20008";
        ram_buffer(50742) := X"00000000";
        ram_buffer(50743) := X"0062102A";
        ram_buffer(50744) := X"10400027";
        ram_buffer(50745) := X"00000000";
        ram_buffer(50746) := X"8FC20024";
        ram_buffer(50747) := X"00000000";
        ram_buffer(50748) := X"3042001F";
        ram_buffer(50749) := X"AFC20024";
        ram_buffer(50750) := X"8FC20024";
        ram_buffer(50751) := X"00000000";
        ram_buffer(50752) := X"1040001F";
        ram_buffer(50753) := X"00000000";
        ram_buffer(50754) := X"8FC20000";
        ram_buffer(50755) := X"00000000";
        ram_buffer(50756) := X"00021080";
        ram_buffer(50757) := X"8FC30004";
        ram_buffer(50758) := X"00000000";
        ram_buffer(50759) := X"00621021";
        ram_buffer(50760) := X"8C420000";
        ram_buffer(50761) := X"00000000";
        ram_buffer(50762) := X"AFC2000C";
        ram_buffer(50763) := X"8FC2000C";
        ram_buffer(50764) := X"00000000";
        ram_buffer(50765) := X"AFC20010";
        ram_buffer(50766) := X"8FC30010";
        ram_buffer(50767) := X"8FC20024";
        ram_buffer(50768) := X"00000000";
        ram_buffer(50769) := X"00431006";
        ram_buffer(50770) := X"AFC20010";
        ram_buffer(50771) := X"8FC30010";
        ram_buffer(50772) := X"8FC20024";
        ram_buffer(50773) := X"00000000";
        ram_buffer(50774) := X"00431004";
        ram_buffer(50775) := X"AFC20010";
        ram_buffer(50776) := X"8FC30010";
        ram_buffer(50777) := X"8FC2000C";
        ram_buffer(50778) := X"00000000";
        ram_buffer(50779) := X"10620004";
        ram_buffer(50780) := X"00000000";
        ram_buffer(50781) := X"24020001";
        ram_buffer(50782) := X"10000021";
        ram_buffer(50783) := X"00000000";
        ram_buffer(50784) := X"8FC20004";
        ram_buffer(50785) := X"00000000";
        ram_buffer(50786) := X"AFC20014";
        ram_buffer(50787) := X"8FC20000";
        ram_buffer(50788) := X"00000000";
        ram_buffer(50789) := X"00021080";
        ram_buffer(50790) := X"8FC30004";
        ram_buffer(50791) := X"00000000";
        ram_buffer(50792) := X"00621021";
        ram_buffer(50793) := X"AFC20004";
        ram_buffer(50794) := X"1000000E";
        ram_buffer(50795) := X"00000000";
        ram_buffer(50796) := X"8FC20004";
        ram_buffer(50797) := X"00000000";
        ram_buffer(50798) := X"2442FFFC";
        ram_buffer(50799) := X"AFC20004";
        ram_buffer(50800) := X"8FC20004";
        ram_buffer(50801) := X"00000000";
        ram_buffer(50802) := X"8C420000";
        ram_buffer(50803) := X"00000000";
        ram_buffer(50804) := X"10400004";
        ram_buffer(50805) := X"00000000";
        ram_buffer(50806) := X"24020001";
        ram_buffer(50807) := X"10000008";
        ram_buffer(50808) := X"00000000";
        ram_buffer(50809) := X"8FC30004";
        ram_buffer(50810) := X"8FC20014";
        ram_buffer(50811) := X"00000000";
        ram_buffer(50812) := X"0043102B";
        ram_buffer(50813) := X"1440FFEE";
        ram_buffer(50814) := X"00000000";
        ram_buffer(50815) := X"00001021";
        ram_buffer(50816) := X"03C0E821";
        ram_buffer(50817) := X"8FBE001C";
        ram_buffer(50818) := X"27BD0020";
        ram_buffer(50819) := X"03E00008";
        ram_buffer(50820) := X"00000000";
        ram_buffer(50821) := X"27BDFFE0";
        ram_buffer(50822) := X"AFBF001C";
        ram_buffer(50823) := X"AFBE0018";
        ram_buffer(50824) := X"03A0F021";
        ram_buffer(50825) := X"AFC40020";
        ram_buffer(50826) := X"AFC50024";
        ram_buffer(50827) := X"AFC60028";
        ram_buffer(50828) := X"AFC7002C";
        ram_buffer(50829) := X"AF8081EC";
        ram_buffer(50830) := X"8FC6002C";
        ram_buffer(50831) := X"8FC50028";
        ram_buffer(50832) := X"8FC40024";
        ram_buffer(50833) := X"0C02FC2E";
        ram_buffer(50834) := X"00000000";
        ram_buffer(50835) := X"AFC20010";
        ram_buffer(50836) := X"8FC30010";
        ram_buffer(50837) := X"2402FFFF";
        ram_buffer(50838) := X"14620009";
        ram_buffer(50839) := X"00000000";
        ram_buffer(50840) := X"8F8281EC";
        ram_buffer(50841) := X"00000000";
        ram_buffer(50842) := X"10400005";
        ram_buffer(50843) := X"00000000";
        ram_buffer(50844) := X"8F8381EC";
        ram_buffer(50845) := X"8FC20020";
        ram_buffer(50846) := X"00000000";
        ram_buffer(50847) := X"AC430000";
        ram_buffer(50848) := X"8FC20010";
        ram_buffer(50849) := X"03C0E821";
        ram_buffer(50850) := X"8FBF001C";
        ram_buffer(50851) := X"8FBE0018";
        ram_buffer(50852) := X"27BD0020";
        ram_buffer(50853) := X"03E00008";
        ram_buffer(50854) := X"00000000";
        ram_buffer(50855) := X"27BDFF80";
        ram_buffer(50856) := X"AFBF007C";
        ram_buffer(50857) := X"AFBE0078";
        ram_buffer(50858) := X"03A0F021";
        ram_buffer(50859) := X"AFC40080";
        ram_buffer(50860) := X"AFC50084";
        ram_buffer(50861) := X"AFC60088";
        ram_buffer(50862) := X"8FC20084";
        ram_buffer(50863) := X"00000000";
        ram_buffer(50864) := X"14400007";
        ram_buffer(50865) := X"00000000";
        ram_buffer(50866) := X"8FC50088";
        ram_buffer(50867) := X"8FC40080";
        ram_buffer(50868) := X"0C027B8F";
        ram_buffer(50869) := X"00000000";
        ram_buffer(50870) := X"10000430";
        ram_buffer(50871) := X"00000000";
        ram_buffer(50872) := X"8FC40080";
        ram_buffer(50873) := X"0C0280C3";
        ram_buffer(50874) := X"00000000";
        ram_buffer(50875) := X"8FC20084";
        ram_buffer(50876) := X"00000000";
        ram_buffer(50877) := X"2442FFF8";
        ram_buffer(50878) := X"AFC20040";
        ram_buffer(50879) := X"8FC20040";
        ram_buffer(50880) := X"00000000";
        ram_buffer(50881) := X"AFC20010";
        ram_buffer(50882) := X"8FC20040";
        ram_buffer(50883) := X"00000000";
        ram_buffer(50884) := X"8C430004";
        ram_buffer(50885) := X"2402FFFC";
        ram_buffer(50886) := X"00621024";
        ram_buffer(50887) := X"AFC20044";
        ram_buffer(50888) := X"8FC20044";
        ram_buffer(50889) := X"00000000";
        ram_buffer(50890) := X"AFC20014";
        ram_buffer(50891) := X"8FC20088";
        ram_buffer(50892) := X"00000000";
        ram_buffer(50893) := X"2442000B";
        ram_buffer(50894) := X"2C420017";
        ram_buffer(50895) := X"14400008";
        ram_buffer(50896) := X"00000000";
        ram_buffer(50897) := X"8FC20088";
        ram_buffer(50898) := X"00000000";
        ram_buffer(50899) := X"2443000B";
        ram_buffer(50900) := X"2402FFF8";
        ram_buffer(50901) := X"00621024";
        ram_buffer(50902) := X"10000002";
        ram_buffer(50903) := X"00000000";
        ram_buffer(50904) := X"24020010";
        ram_buffer(50905) := X"AFC20048";
        ram_buffer(50906) := X"8FC20048";
        ram_buffer(50907) := X"00000000";
        ram_buffer(50908) := X"04400007";
        ram_buffer(50909) := X"00000000";
        ram_buffer(50910) := X"8FC30048";
        ram_buffer(50911) := X"8FC20088";
        ram_buffer(50912) := X"00000000";
        ram_buffer(50913) := X"0062102B";
        ram_buffer(50914) := X"10400007";
        ram_buffer(50915) := X"00000000";
        ram_buffer(50916) := X"8FC20080";
        ram_buffer(50917) := X"2403000C";
        ram_buffer(50918) := X"AC430000";
        ram_buffer(50919) := X"00001021";
        ram_buffer(50920) := X"100003FE";
        ram_buffer(50921) := X"00000000";
        ram_buffer(50922) := X"8FC30044";
        ram_buffer(50923) := X"8FC20048";
        ram_buffer(50924) := X"00000000";
        ram_buffer(50925) := X"0062102A";
        ram_buffer(50926) := X"104003A6";
        ram_buffer(50927) := X"00000000";
        ram_buffer(50928) := X"8FC30040";
        ram_buffer(50929) := X"8FC20044";
        ram_buffer(50930) := X"00000000";
        ram_buffer(50931) := X"00621021";
        ram_buffer(50932) := X"AFC20018";
        ram_buffer(50933) := X"3C02100D";
        ram_buffer(50934) := X"2442CBE0";
        ram_buffer(50935) := X"8C430008";
        ram_buffer(50936) := X"8FC20018";
        ram_buffer(50937) := X"00000000";
        ram_buffer(50938) := X"1062000E";
        ram_buffer(50939) := X"00000000";
        ram_buffer(50940) := X"8FC20018";
        ram_buffer(50941) := X"00000000";
        ram_buffer(50942) := X"8C430004";
        ram_buffer(50943) := X"2402FFFE";
        ram_buffer(50944) := X"00621024";
        ram_buffer(50945) := X"8FC30018";
        ram_buffer(50946) := X"00000000";
        ram_buffer(50947) := X"00621021";
        ram_buffer(50948) := X"8C420004";
        ram_buffer(50949) := X"00000000";
        ram_buffer(50950) := X"30420001";
        ram_buffer(50951) := X"14400064";
        ram_buffer(50952) := X"00000000";
        ram_buffer(50953) := X"8FC20018";
        ram_buffer(50954) := X"00000000";
        ram_buffer(50955) := X"8C430004";
        ram_buffer(50956) := X"2402FFFC";
        ram_buffer(50957) := X"00621024";
        ram_buffer(50958) := X"AFC2001C";
        ram_buffer(50959) := X"3C02100D";
        ram_buffer(50960) := X"2442CBE0";
        ram_buffer(50961) := X"8C430008";
        ram_buffer(50962) := X"8FC20018";
        ram_buffer(50963) := X"00000000";
        ram_buffer(50964) := X"14620034";
        ram_buffer(50965) := X"00000000";
        ram_buffer(50966) := X"8FC3001C";
        ram_buffer(50967) := X"8FC20014";
        ram_buffer(50968) := X"00000000";
        ram_buffer(50969) := X"00621021";
        ram_buffer(50970) := X"00401821";
        ram_buffer(50971) := X"8FC20048";
        ram_buffer(50972) := X"00000000";
        ram_buffer(50973) := X"24420010";
        ram_buffer(50974) := X"0062102A";
        ram_buffer(50975) := X"14400050";
        ram_buffer(50976) := X"00000000";
        ram_buffer(50977) := X"8FC30014";
        ram_buffer(50978) := X"8FC2001C";
        ram_buffer(50979) := X"00000000";
        ram_buffer(50980) := X"00621021";
        ram_buffer(50981) := X"AFC20014";
        ram_buffer(50982) := X"3C02100D";
        ram_buffer(50983) := X"2442CBE0";
        ram_buffer(50984) := X"8FC40040";
        ram_buffer(50985) := X"8FC30048";
        ram_buffer(50986) := X"00000000";
        ram_buffer(50987) := X"00831821";
        ram_buffer(50988) := X"AC430008";
        ram_buffer(50989) := X"3C02100D";
        ram_buffer(50990) := X"2442CBE0";
        ram_buffer(50991) := X"8C420008";
        ram_buffer(50992) := X"8FC40014";
        ram_buffer(50993) := X"8FC30048";
        ram_buffer(50994) := X"00000000";
        ram_buffer(50995) := X"00831823";
        ram_buffer(50996) := X"34630001";
        ram_buffer(50997) := X"AC430004";
        ram_buffer(50998) := X"8FC20040";
        ram_buffer(50999) := X"00000000";
        ram_buffer(51000) := X"8C420004";
        ram_buffer(51001) := X"00000000";
        ram_buffer(51002) := X"30430001";
        ram_buffer(51003) := X"8FC20048";
        ram_buffer(51004) := X"00000000";
        ram_buffer(51005) := X"00621825";
        ram_buffer(51006) := X"8FC20040";
        ram_buffer(51007) := X"00000000";
        ram_buffer(51008) := X"AC430004";
        ram_buffer(51009) := X"8FC40080";
        ram_buffer(51010) := X"0C0280CD";
        ram_buffer(51011) := X"00000000";
        ram_buffer(51012) := X"8FC20040";
        ram_buffer(51013) := X"00000000";
        ram_buffer(51014) := X"24420008";
        ram_buffer(51015) := X"1000039F";
        ram_buffer(51016) := X"00000000";
        ram_buffer(51017) := X"8FC3001C";
        ram_buffer(51018) := X"8FC20014";
        ram_buffer(51019) := X"00000000";
        ram_buffer(51020) := X"00621021";
        ram_buffer(51021) := X"00401821";
        ram_buffer(51022) := X"8FC20048";
        ram_buffer(51023) := X"00000000";
        ram_buffer(51024) := X"0062102A";
        ram_buffer(51025) := X"1440001E";
        ram_buffer(51026) := X"00000000";
        ram_buffer(51027) := X"8FC20018";
        ram_buffer(51028) := X"00000000";
        ram_buffer(51029) := X"8C42000C";
        ram_buffer(51030) := X"00000000";
        ram_buffer(51031) := X"AFC2004C";
        ram_buffer(51032) := X"8FC20018";
        ram_buffer(51033) := X"00000000";
        ram_buffer(51034) := X"8C420008";
        ram_buffer(51035) := X"00000000";
        ram_buffer(51036) := X"AFC20050";
        ram_buffer(51037) := X"8FC20050";
        ram_buffer(51038) := X"8FC3004C";
        ram_buffer(51039) := X"00000000";
        ram_buffer(51040) := X"AC43000C";
        ram_buffer(51041) := X"8FC2004C";
        ram_buffer(51042) := X"8FC30050";
        ram_buffer(51043) := X"00000000";
        ram_buffer(51044) := X"AC430008";
        ram_buffer(51045) := X"8FC30014";
        ram_buffer(51046) := X"8FC2001C";
        ram_buffer(51047) := X"00000000";
        ram_buffer(51048) := X"00621021";
        ram_buffer(51049) := X"AFC20014";
        ram_buffer(51050) := X"1000032A";
        ram_buffer(51051) := X"00000000";
        ram_buffer(51052) := X"AFC00018";
        ram_buffer(51053) := X"AFC0001C";
        ram_buffer(51054) := X"10000002";
        ram_buffer(51055) := X"00000000";
        ram_buffer(51056) := X"00000000";
        ram_buffer(51057) := X"8FC20040";
        ram_buffer(51058) := X"00000000";
        ram_buffer(51059) := X"8C420004";
        ram_buffer(51060) := X"00000000";
        ram_buffer(51061) := X"30420001";
        ram_buffer(51062) := X"14400264";
        ram_buffer(51063) := X"00000000";
        ram_buffer(51064) := X"8FC20040";
        ram_buffer(51065) := X"00000000";
        ram_buffer(51066) := X"8C420000";
        ram_buffer(51067) := X"00000000";
        ram_buffer(51068) := X"00021023";
        ram_buffer(51069) := X"8FC30040";
        ram_buffer(51070) := X"00000000";
        ram_buffer(51071) := X"00621021";
        ram_buffer(51072) := X"AFC20054";
        ram_buffer(51073) := X"8FC20054";
        ram_buffer(51074) := X"00000000";
        ram_buffer(51075) := X"8C430004";
        ram_buffer(51076) := X"2402FFFC";
        ram_buffer(51077) := X"00621024";
        ram_buffer(51078) := X"AFC20058";
        ram_buffer(51079) := X"8FC20018";
        ram_buffer(51080) := X"00000000";
        ram_buffer(51081) := X"104001A0";
        ram_buffer(51082) := X"00000000";
        ram_buffer(51083) := X"3C02100D";
        ram_buffer(51084) := X"2442CBE0";
        ram_buffer(51085) := X"8C430008";
        ram_buffer(51086) := X"8FC20018";
        ram_buffer(51087) := X"00000000";
        ram_buffer(51088) := X"146200D4";
        ram_buffer(51089) := X"00000000";
        ram_buffer(51090) := X"8FC3001C";
        ram_buffer(51091) := X"8FC20058";
        ram_buffer(51092) := X"00000000";
        ram_buffer(51093) := X"00621821";
        ram_buffer(51094) := X"8FC20014";
        ram_buffer(51095) := X"00000000";
        ram_buffer(51096) := X"00621021";
        ram_buffer(51097) := X"00401821";
        ram_buffer(51098) := X"8FC20048";
        ram_buffer(51099) := X"00000000";
        ram_buffer(51100) := X"24420010";
        ram_buffer(51101) := X"0062102A";
        ram_buffer(51102) := X"1440018B";
        ram_buffer(51103) := X"00000000";
        ram_buffer(51104) := X"8FC20054";
        ram_buffer(51105) := X"00000000";
        ram_buffer(51106) := X"8C42000C";
        ram_buffer(51107) := X"00000000";
        ram_buffer(51108) := X"AFC2004C";
        ram_buffer(51109) := X"8FC20054";
        ram_buffer(51110) := X"00000000";
        ram_buffer(51111) := X"8C420008";
        ram_buffer(51112) := X"00000000";
        ram_buffer(51113) := X"AFC20050";
        ram_buffer(51114) := X"8FC20050";
        ram_buffer(51115) := X"8FC3004C";
        ram_buffer(51116) := X"00000000";
        ram_buffer(51117) := X"AC43000C";
        ram_buffer(51118) := X"8FC2004C";
        ram_buffer(51119) := X"8FC30050";
        ram_buffer(51120) := X"00000000";
        ram_buffer(51121) := X"AC430008";
        ram_buffer(51122) := X"8FC20054";
        ram_buffer(51123) := X"00000000";
        ram_buffer(51124) := X"AFC20010";
        ram_buffer(51125) := X"8FC30058";
        ram_buffer(51126) := X"8FC2001C";
        ram_buffer(51127) := X"00000000";
        ram_buffer(51128) := X"00621021";
        ram_buffer(51129) := X"8FC30014";
        ram_buffer(51130) := X"00000000";
        ram_buffer(51131) := X"00621021";
        ram_buffer(51132) := X"AFC20014";
        ram_buffer(51133) := X"8FC20010";
        ram_buffer(51134) := X"00000000";
        ram_buffer(51135) := X"24420008";
        ram_buffer(51136) := X"AFC2005C";
        ram_buffer(51137) := X"8FC20044";
        ram_buffer(51138) := X"00000000";
        ram_buffer(51139) := X"2442FFFC";
        ram_buffer(51140) := X"AFC20060";
        ram_buffer(51141) := X"8FC20060";
        ram_buffer(51142) := X"00000000";
        ram_buffer(51143) := X"2C420025";
        ram_buffer(51144) := X"10400076";
        ram_buffer(51145) := X"00000000";
        ram_buffer(51146) := X"8FC20084";
        ram_buffer(51147) := X"00000000";
        ram_buffer(51148) := X"AFC20020";
        ram_buffer(51149) := X"8FC2005C";
        ram_buffer(51150) := X"00000000";
        ram_buffer(51151) := X"AFC20024";
        ram_buffer(51152) := X"8FC20060";
        ram_buffer(51153) := X"00000000";
        ram_buffer(51154) := X"2C420014";
        ram_buffer(51155) := X"1440004D";
        ram_buffer(51156) := X"00000000";
        ram_buffer(51157) := X"8FC20024";
        ram_buffer(51158) := X"00000000";
        ram_buffer(51159) := X"24430004";
        ram_buffer(51160) := X"AFC30024";
        ram_buffer(51161) := X"8FC30020";
        ram_buffer(51162) := X"00000000";
        ram_buffer(51163) := X"24640004";
        ram_buffer(51164) := X"AFC40020";
        ram_buffer(51165) := X"8C630000";
        ram_buffer(51166) := X"00000000";
        ram_buffer(51167) := X"AC430000";
        ram_buffer(51168) := X"8FC20024";
        ram_buffer(51169) := X"00000000";
        ram_buffer(51170) := X"24430004";
        ram_buffer(51171) := X"AFC30024";
        ram_buffer(51172) := X"8FC30020";
        ram_buffer(51173) := X"00000000";
        ram_buffer(51174) := X"24640004";
        ram_buffer(51175) := X"AFC40020";
        ram_buffer(51176) := X"8C630000";
        ram_buffer(51177) := X"00000000";
        ram_buffer(51178) := X"AC430000";
        ram_buffer(51179) := X"8FC20060";
        ram_buffer(51180) := X"00000000";
        ram_buffer(51181) := X"2C42001C";
        ram_buffer(51182) := X"14400032";
        ram_buffer(51183) := X"00000000";
        ram_buffer(51184) := X"8FC20024";
        ram_buffer(51185) := X"00000000";
        ram_buffer(51186) := X"24430004";
        ram_buffer(51187) := X"AFC30024";
        ram_buffer(51188) := X"8FC30020";
        ram_buffer(51189) := X"00000000";
        ram_buffer(51190) := X"24640004";
        ram_buffer(51191) := X"AFC40020";
        ram_buffer(51192) := X"8C630000";
        ram_buffer(51193) := X"00000000";
        ram_buffer(51194) := X"AC430000";
        ram_buffer(51195) := X"8FC20024";
        ram_buffer(51196) := X"00000000";
        ram_buffer(51197) := X"24430004";
        ram_buffer(51198) := X"AFC30024";
        ram_buffer(51199) := X"8FC30020";
        ram_buffer(51200) := X"00000000";
        ram_buffer(51201) := X"24640004";
        ram_buffer(51202) := X"AFC40020";
        ram_buffer(51203) := X"8C630000";
        ram_buffer(51204) := X"00000000";
        ram_buffer(51205) := X"AC430000";
        ram_buffer(51206) := X"8FC20060";
        ram_buffer(51207) := X"00000000";
        ram_buffer(51208) := X"2C420024";
        ram_buffer(51209) := X"14400017";
        ram_buffer(51210) := X"00000000";
        ram_buffer(51211) := X"8FC20024";
        ram_buffer(51212) := X"00000000";
        ram_buffer(51213) := X"24430004";
        ram_buffer(51214) := X"AFC30024";
        ram_buffer(51215) := X"8FC30020";
        ram_buffer(51216) := X"00000000";
        ram_buffer(51217) := X"24640004";
        ram_buffer(51218) := X"AFC40020";
        ram_buffer(51219) := X"8C630000";
        ram_buffer(51220) := X"00000000";
        ram_buffer(51221) := X"AC430000";
        ram_buffer(51222) := X"8FC20024";
        ram_buffer(51223) := X"00000000";
        ram_buffer(51224) := X"24430004";
        ram_buffer(51225) := X"AFC30024";
        ram_buffer(51226) := X"8FC30020";
        ram_buffer(51227) := X"00000000";
        ram_buffer(51228) := X"24640004";
        ram_buffer(51229) := X"AFC40020";
        ram_buffer(51230) := X"8C630000";
        ram_buffer(51231) := X"00000000";
        ram_buffer(51232) := X"AC430000";
        ram_buffer(51233) := X"8FC20024";
        ram_buffer(51234) := X"00000000";
        ram_buffer(51235) := X"24430004";
        ram_buffer(51236) := X"AFC30024";
        ram_buffer(51237) := X"8FC30020";
        ram_buffer(51238) := X"00000000";
        ram_buffer(51239) := X"24640004";
        ram_buffer(51240) := X"AFC40020";
        ram_buffer(51241) := X"8C630000";
        ram_buffer(51242) := X"00000000";
        ram_buffer(51243) := X"AC430000";
        ram_buffer(51244) := X"8FC20024";
        ram_buffer(51245) := X"00000000";
        ram_buffer(51246) := X"24430004";
        ram_buffer(51247) := X"AFC30024";
        ram_buffer(51248) := X"8FC30020";
        ram_buffer(51249) := X"00000000";
        ram_buffer(51250) := X"24640004";
        ram_buffer(51251) := X"AFC40020";
        ram_buffer(51252) := X"8C630000";
        ram_buffer(51253) := X"00000000";
        ram_buffer(51254) := X"AC430000";
        ram_buffer(51255) := X"8FC20020";
        ram_buffer(51256) := X"00000000";
        ram_buffer(51257) := X"8C430000";
        ram_buffer(51258) := X"8FC20024";
        ram_buffer(51259) := X"00000000";
        ram_buffer(51260) := X"AC430000";
        ram_buffer(51261) := X"10000006";
        ram_buffer(51262) := X"00000000";
        ram_buffer(51263) := X"8FC60060";
        ram_buffer(51264) := X"8FC50084";
        ram_buffer(51265) := X"8FC4005C";
        ram_buffer(51266) := X"0C02BCED";
        ram_buffer(51267) := X"00000000";
        ram_buffer(51268) := X"3C02100D";
        ram_buffer(51269) := X"2442CBE0";
        ram_buffer(51270) := X"8FC40010";
        ram_buffer(51271) := X"8FC30048";
        ram_buffer(51272) := X"00000000";
        ram_buffer(51273) := X"00831821";
        ram_buffer(51274) := X"AC430008";
        ram_buffer(51275) := X"3C02100D";
        ram_buffer(51276) := X"2442CBE0";
        ram_buffer(51277) := X"8C420008";
        ram_buffer(51278) := X"8FC40014";
        ram_buffer(51279) := X"8FC30048";
        ram_buffer(51280) := X"00000000";
        ram_buffer(51281) := X"00831823";
        ram_buffer(51282) := X"34630001";
        ram_buffer(51283) := X"AC430004";
        ram_buffer(51284) := X"8FC20010";
        ram_buffer(51285) := X"00000000";
        ram_buffer(51286) := X"8C420004";
        ram_buffer(51287) := X"00000000";
        ram_buffer(51288) := X"30430001";
        ram_buffer(51289) := X"8FC20048";
        ram_buffer(51290) := X"00000000";
        ram_buffer(51291) := X"00621825";
        ram_buffer(51292) := X"8FC20010";
        ram_buffer(51293) := X"00000000";
        ram_buffer(51294) := X"AC430004";
        ram_buffer(51295) := X"8FC40080";
        ram_buffer(51296) := X"0C0280CD";
        ram_buffer(51297) := X"00000000";
        ram_buffer(51298) := X"8FC2005C";
        ram_buffer(51299) := X"10000283";
        ram_buffer(51300) := X"00000000";
        ram_buffer(51301) := X"8FC3001C";
        ram_buffer(51302) := X"8FC20058";
        ram_buffer(51303) := X"00000000";
        ram_buffer(51304) := X"00621821";
        ram_buffer(51305) := X"8FC20014";
        ram_buffer(51306) := X"00000000";
        ram_buffer(51307) := X"00621021";
        ram_buffer(51308) := X"00401821";
        ram_buffer(51309) := X"8FC20048";
        ram_buffer(51310) := X"00000000";
        ram_buffer(51311) := X"0062102A";
        ram_buffer(51312) := X"144000B9";
        ram_buffer(51313) := X"00000000";
        ram_buffer(51314) := X"8FC20018";
        ram_buffer(51315) := X"00000000";
        ram_buffer(51316) := X"8C42000C";
        ram_buffer(51317) := X"00000000";
        ram_buffer(51318) := X"AFC2004C";
        ram_buffer(51319) := X"8FC20018";
        ram_buffer(51320) := X"00000000";
        ram_buffer(51321) := X"8C420008";
        ram_buffer(51322) := X"00000000";
        ram_buffer(51323) := X"AFC20050";
        ram_buffer(51324) := X"8FC20050";
        ram_buffer(51325) := X"8FC3004C";
        ram_buffer(51326) := X"00000000";
        ram_buffer(51327) := X"AC43000C";
        ram_buffer(51328) := X"8FC2004C";
        ram_buffer(51329) := X"8FC30050";
        ram_buffer(51330) := X"00000000";
        ram_buffer(51331) := X"AC430008";
        ram_buffer(51332) := X"8FC20054";
        ram_buffer(51333) := X"00000000";
        ram_buffer(51334) := X"8C42000C";
        ram_buffer(51335) := X"00000000";
        ram_buffer(51336) := X"AFC2004C";
        ram_buffer(51337) := X"8FC20054";
        ram_buffer(51338) := X"00000000";
        ram_buffer(51339) := X"8C420008";
        ram_buffer(51340) := X"00000000";
        ram_buffer(51341) := X"AFC20050";
        ram_buffer(51342) := X"8FC20050";
        ram_buffer(51343) := X"8FC3004C";
        ram_buffer(51344) := X"00000000";
        ram_buffer(51345) := X"AC43000C";
        ram_buffer(51346) := X"8FC2004C";
        ram_buffer(51347) := X"8FC30050";
        ram_buffer(51348) := X"00000000";
        ram_buffer(51349) := X"AC430008";
        ram_buffer(51350) := X"8FC20054";
        ram_buffer(51351) := X"00000000";
        ram_buffer(51352) := X"AFC20010";
        ram_buffer(51353) := X"8FC3001C";
        ram_buffer(51354) := X"8FC20058";
        ram_buffer(51355) := X"00000000";
        ram_buffer(51356) := X"00621021";
        ram_buffer(51357) := X"8FC30014";
        ram_buffer(51358) := X"00000000";
        ram_buffer(51359) := X"00621021";
        ram_buffer(51360) := X"AFC20014";
        ram_buffer(51361) := X"8FC20010";
        ram_buffer(51362) := X"00000000";
        ram_buffer(51363) := X"24420008";
        ram_buffer(51364) := X"AFC2005C";
        ram_buffer(51365) := X"8FC20044";
        ram_buffer(51366) := X"00000000";
        ram_buffer(51367) := X"2442FFFC";
        ram_buffer(51368) := X"AFC20064";
        ram_buffer(51369) := X"8FC20064";
        ram_buffer(51370) := X"00000000";
        ram_buffer(51371) := X"2C420025";
        ram_buffer(51372) := X"10400076";
        ram_buffer(51373) := X"00000000";
        ram_buffer(51374) := X"8FC20084";
        ram_buffer(51375) := X"00000000";
        ram_buffer(51376) := X"AFC20028";
        ram_buffer(51377) := X"8FC2005C";
        ram_buffer(51378) := X"00000000";
        ram_buffer(51379) := X"AFC2002C";
        ram_buffer(51380) := X"8FC20064";
        ram_buffer(51381) := X"00000000";
        ram_buffer(51382) := X"2C420014";
        ram_buffer(51383) := X"1440004D";
        ram_buffer(51384) := X"00000000";
        ram_buffer(51385) := X"8FC2002C";
        ram_buffer(51386) := X"00000000";
        ram_buffer(51387) := X"24430004";
        ram_buffer(51388) := X"AFC3002C";
        ram_buffer(51389) := X"8FC30028";
        ram_buffer(51390) := X"00000000";
        ram_buffer(51391) := X"24640004";
        ram_buffer(51392) := X"AFC40028";
        ram_buffer(51393) := X"8C630000";
        ram_buffer(51394) := X"00000000";
        ram_buffer(51395) := X"AC430000";
        ram_buffer(51396) := X"8FC2002C";
        ram_buffer(51397) := X"00000000";
        ram_buffer(51398) := X"24430004";
        ram_buffer(51399) := X"AFC3002C";
        ram_buffer(51400) := X"8FC30028";
        ram_buffer(51401) := X"00000000";
        ram_buffer(51402) := X"24640004";
        ram_buffer(51403) := X"AFC40028";
        ram_buffer(51404) := X"8C630000";
        ram_buffer(51405) := X"00000000";
        ram_buffer(51406) := X"AC430000";
        ram_buffer(51407) := X"8FC20064";
        ram_buffer(51408) := X"00000000";
        ram_buffer(51409) := X"2C42001C";
        ram_buffer(51410) := X"14400032";
        ram_buffer(51411) := X"00000000";
        ram_buffer(51412) := X"8FC2002C";
        ram_buffer(51413) := X"00000000";
        ram_buffer(51414) := X"24430004";
        ram_buffer(51415) := X"AFC3002C";
        ram_buffer(51416) := X"8FC30028";
        ram_buffer(51417) := X"00000000";
        ram_buffer(51418) := X"24640004";
        ram_buffer(51419) := X"AFC40028";
        ram_buffer(51420) := X"8C630000";
        ram_buffer(51421) := X"00000000";
        ram_buffer(51422) := X"AC430000";
        ram_buffer(51423) := X"8FC2002C";
        ram_buffer(51424) := X"00000000";
        ram_buffer(51425) := X"24430004";
        ram_buffer(51426) := X"AFC3002C";
        ram_buffer(51427) := X"8FC30028";
        ram_buffer(51428) := X"00000000";
        ram_buffer(51429) := X"24640004";
        ram_buffer(51430) := X"AFC40028";
        ram_buffer(51431) := X"8C630000";
        ram_buffer(51432) := X"00000000";
        ram_buffer(51433) := X"AC430000";
        ram_buffer(51434) := X"8FC20064";
        ram_buffer(51435) := X"00000000";
        ram_buffer(51436) := X"2C420024";
        ram_buffer(51437) := X"14400017";
        ram_buffer(51438) := X"00000000";
        ram_buffer(51439) := X"8FC2002C";
        ram_buffer(51440) := X"00000000";
        ram_buffer(51441) := X"24430004";
        ram_buffer(51442) := X"AFC3002C";
        ram_buffer(51443) := X"8FC30028";
        ram_buffer(51444) := X"00000000";
        ram_buffer(51445) := X"24640004";
        ram_buffer(51446) := X"AFC40028";
        ram_buffer(51447) := X"8C630000";
        ram_buffer(51448) := X"00000000";
        ram_buffer(51449) := X"AC430000";
        ram_buffer(51450) := X"8FC2002C";
        ram_buffer(51451) := X"00000000";
        ram_buffer(51452) := X"24430004";
        ram_buffer(51453) := X"AFC3002C";
        ram_buffer(51454) := X"8FC30028";
        ram_buffer(51455) := X"00000000";
        ram_buffer(51456) := X"24640004";
        ram_buffer(51457) := X"AFC40028";
        ram_buffer(51458) := X"8C630000";
        ram_buffer(51459) := X"00000000";
        ram_buffer(51460) := X"AC430000";
        ram_buffer(51461) := X"8FC2002C";
        ram_buffer(51462) := X"00000000";
        ram_buffer(51463) := X"24430004";
        ram_buffer(51464) := X"AFC3002C";
        ram_buffer(51465) := X"8FC30028";
        ram_buffer(51466) := X"00000000";
        ram_buffer(51467) := X"24640004";
        ram_buffer(51468) := X"AFC40028";
        ram_buffer(51469) := X"8C630000";
        ram_buffer(51470) := X"00000000";
        ram_buffer(51471) := X"AC430000";
        ram_buffer(51472) := X"8FC2002C";
        ram_buffer(51473) := X"00000000";
        ram_buffer(51474) := X"24430004";
        ram_buffer(51475) := X"AFC3002C";
        ram_buffer(51476) := X"8FC30028";
        ram_buffer(51477) := X"00000000";
        ram_buffer(51478) := X"24640004";
        ram_buffer(51479) := X"AFC40028";
        ram_buffer(51480) := X"8C630000";
        ram_buffer(51481) := X"00000000";
        ram_buffer(51482) := X"AC430000";
        ram_buffer(51483) := X"8FC20028";
        ram_buffer(51484) := X"00000000";
        ram_buffer(51485) := X"8C430000";
        ram_buffer(51486) := X"8FC2002C";
        ram_buffer(51487) := X"00000000";
        ram_buffer(51488) := X"AC430000";
        ram_buffer(51489) := X"10000173";
        ram_buffer(51490) := X"00000000";
        ram_buffer(51491) := X"8FC60064";
        ram_buffer(51492) := X"8FC50084";
        ram_buffer(51493) := X"8FC4005C";
        ram_buffer(51494) := X"0C02BCED";
        ram_buffer(51495) := X"00000000";
        ram_buffer(51496) := X"1000016C";
        ram_buffer(51497) := X"00000000";
        ram_buffer(51498) := X"8FC20054";
        ram_buffer(51499) := X"00000000";
        ram_buffer(51500) := X"104000AE";
        ram_buffer(51501) := X"00000000";
        ram_buffer(51502) := X"8FC30058";
        ram_buffer(51503) := X"8FC20014";
        ram_buffer(51504) := X"00000000";
        ram_buffer(51505) := X"00621021";
        ram_buffer(51506) := X"00401821";
        ram_buffer(51507) := X"8FC20048";
        ram_buffer(51508) := X"00000000";
        ram_buffer(51509) := X"0062102A";
        ram_buffer(51510) := X"144000A4";
        ram_buffer(51511) := X"00000000";
        ram_buffer(51512) := X"8FC20054";
        ram_buffer(51513) := X"00000000";
        ram_buffer(51514) := X"8C42000C";
        ram_buffer(51515) := X"00000000";
        ram_buffer(51516) := X"AFC2004C";
        ram_buffer(51517) := X"8FC20054";
        ram_buffer(51518) := X"00000000";
        ram_buffer(51519) := X"8C420008";
        ram_buffer(51520) := X"00000000";
        ram_buffer(51521) := X"AFC20050";
        ram_buffer(51522) := X"8FC20050";
        ram_buffer(51523) := X"8FC3004C";
        ram_buffer(51524) := X"00000000";
        ram_buffer(51525) := X"AC43000C";
        ram_buffer(51526) := X"8FC2004C";
        ram_buffer(51527) := X"8FC30050";
        ram_buffer(51528) := X"00000000";
        ram_buffer(51529) := X"AC430008";
        ram_buffer(51530) := X"8FC20054";
        ram_buffer(51531) := X"00000000";
        ram_buffer(51532) := X"AFC20010";
        ram_buffer(51533) := X"8FC30014";
        ram_buffer(51534) := X"8FC20058";
        ram_buffer(51535) := X"00000000";
        ram_buffer(51536) := X"00621021";
        ram_buffer(51537) := X"AFC20014";
        ram_buffer(51538) := X"8FC20010";
        ram_buffer(51539) := X"00000000";
        ram_buffer(51540) := X"24420008";
        ram_buffer(51541) := X"AFC2005C";
        ram_buffer(51542) := X"8FC20044";
        ram_buffer(51543) := X"00000000";
        ram_buffer(51544) := X"2442FFFC";
        ram_buffer(51545) := X"AFC20068";
        ram_buffer(51546) := X"8FC20068";
        ram_buffer(51547) := X"00000000";
        ram_buffer(51548) := X"2C420025";
        ram_buffer(51549) := X"10400076";
        ram_buffer(51550) := X"00000000";
        ram_buffer(51551) := X"8FC20084";
        ram_buffer(51552) := X"00000000";
        ram_buffer(51553) := X"AFC20030";
        ram_buffer(51554) := X"8FC2005C";
        ram_buffer(51555) := X"00000000";
        ram_buffer(51556) := X"AFC20034";
        ram_buffer(51557) := X"8FC20068";
        ram_buffer(51558) := X"00000000";
        ram_buffer(51559) := X"2C420014";
        ram_buffer(51560) := X"1440004D";
        ram_buffer(51561) := X"00000000";
        ram_buffer(51562) := X"8FC20034";
        ram_buffer(51563) := X"00000000";
        ram_buffer(51564) := X"24430004";
        ram_buffer(51565) := X"AFC30034";
        ram_buffer(51566) := X"8FC30030";
        ram_buffer(51567) := X"00000000";
        ram_buffer(51568) := X"24640004";
        ram_buffer(51569) := X"AFC40030";
        ram_buffer(51570) := X"8C630000";
        ram_buffer(51571) := X"00000000";
        ram_buffer(51572) := X"AC430000";
        ram_buffer(51573) := X"8FC20034";
        ram_buffer(51574) := X"00000000";
        ram_buffer(51575) := X"24430004";
        ram_buffer(51576) := X"AFC30034";
        ram_buffer(51577) := X"8FC30030";
        ram_buffer(51578) := X"00000000";
        ram_buffer(51579) := X"24640004";
        ram_buffer(51580) := X"AFC40030";
        ram_buffer(51581) := X"8C630000";
        ram_buffer(51582) := X"00000000";
        ram_buffer(51583) := X"AC430000";
        ram_buffer(51584) := X"8FC20068";
        ram_buffer(51585) := X"00000000";
        ram_buffer(51586) := X"2C42001C";
        ram_buffer(51587) := X"14400032";
        ram_buffer(51588) := X"00000000";
        ram_buffer(51589) := X"8FC20034";
        ram_buffer(51590) := X"00000000";
        ram_buffer(51591) := X"24430004";
        ram_buffer(51592) := X"AFC30034";
        ram_buffer(51593) := X"8FC30030";
        ram_buffer(51594) := X"00000000";
        ram_buffer(51595) := X"24640004";
        ram_buffer(51596) := X"AFC40030";
        ram_buffer(51597) := X"8C630000";
        ram_buffer(51598) := X"00000000";
        ram_buffer(51599) := X"AC430000";
        ram_buffer(51600) := X"8FC20034";
        ram_buffer(51601) := X"00000000";
        ram_buffer(51602) := X"24430004";
        ram_buffer(51603) := X"AFC30034";
        ram_buffer(51604) := X"8FC30030";
        ram_buffer(51605) := X"00000000";
        ram_buffer(51606) := X"24640004";
        ram_buffer(51607) := X"AFC40030";
        ram_buffer(51608) := X"8C630000";
        ram_buffer(51609) := X"00000000";
        ram_buffer(51610) := X"AC430000";
        ram_buffer(51611) := X"8FC20068";
        ram_buffer(51612) := X"00000000";
        ram_buffer(51613) := X"2C420024";
        ram_buffer(51614) := X"14400017";
        ram_buffer(51615) := X"00000000";
        ram_buffer(51616) := X"8FC20034";
        ram_buffer(51617) := X"00000000";
        ram_buffer(51618) := X"24430004";
        ram_buffer(51619) := X"AFC30034";
        ram_buffer(51620) := X"8FC30030";
        ram_buffer(51621) := X"00000000";
        ram_buffer(51622) := X"24640004";
        ram_buffer(51623) := X"AFC40030";
        ram_buffer(51624) := X"8C630000";
        ram_buffer(51625) := X"00000000";
        ram_buffer(51626) := X"AC430000";
        ram_buffer(51627) := X"8FC20034";
        ram_buffer(51628) := X"00000000";
        ram_buffer(51629) := X"24430004";
        ram_buffer(51630) := X"AFC30034";
        ram_buffer(51631) := X"8FC30030";
        ram_buffer(51632) := X"00000000";
        ram_buffer(51633) := X"24640004";
        ram_buffer(51634) := X"AFC40030";
        ram_buffer(51635) := X"8C630000";
        ram_buffer(51636) := X"00000000";
        ram_buffer(51637) := X"AC430000";
        ram_buffer(51638) := X"8FC20034";
        ram_buffer(51639) := X"00000000";
        ram_buffer(51640) := X"24430004";
        ram_buffer(51641) := X"AFC30034";
        ram_buffer(51642) := X"8FC30030";
        ram_buffer(51643) := X"00000000";
        ram_buffer(51644) := X"24640004";
        ram_buffer(51645) := X"AFC40030";
        ram_buffer(51646) := X"8C630000";
        ram_buffer(51647) := X"00000000";
        ram_buffer(51648) := X"AC430000";
        ram_buffer(51649) := X"8FC20034";
        ram_buffer(51650) := X"00000000";
        ram_buffer(51651) := X"24430004";
        ram_buffer(51652) := X"AFC30034";
        ram_buffer(51653) := X"8FC30030";
        ram_buffer(51654) := X"00000000";
        ram_buffer(51655) := X"24640004";
        ram_buffer(51656) := X"AFC40030";
        ram_buffer(51657) := X"8C630000";
        ram_buffer(51658) := X"00000000";
        ram_buffer(51659) := X"AC430000";
        ram_buffer(51660) := X"8FC20030";
        ram_buffer(51661) := X"00000000";
        ram_buffer(51662) := X"8C430000";
        ram_buffer(51663) := X"8FC20034";
        ram_buffer(51664) := X"00000000";
        ram_buffer(51665) := X"AC430000";
        ram_buffer(51666) := X"100000C2";
        ram_buffer(51667) := X"00000000";
        ram_buffer(51668) := X"8FC60068";
        ram_buffer(51669) := X"8FC50084";
        ram_buffer(51670) := X"8FC4005C";
        ram_buffer(51671) := X"0C02BCED";
        ram_buffer(51672) := X"00000000";
        ram_buffer(51673) := X"100000BB";
        ram_buffer(51674) := X"00000000";
        ram_buffer(51675) := X"8FC50088";
        ram_buffer(51676) := X"8FC40080";
        ram_buffer(51677) := X"0C027B8F";
        ram_buffer(51678) := X"00000000";
        ram_buffer(51679) := X"AFC2005C";
        ram_buffer(51680) := X"8FC2005C";
        ram_buffer(51681) := X"00000000";
        ram_buffer(51682) := X"14400007";
        ram_buffer(51683) := X"00000000";
        ram_buffer(51684) := X"8FC40080";
        ram_buffer(51685) := X"0C0280CD";
        ram_buffer(51686) := X"00000000";
        ram_buffer(51687) := X"00001021";
        ram_buffer(51688) := X"100000FE";
        ram_buffer(51689) := X"00000000";
        ram_buffer(51690) := X"8FC2005C";
        ram_buffer(51691) := X"00000000";
        ram_buffer(51692) := X"2442FFF8";
        ram_buffer(51693) := X"AFC20010";
        ram_buffer(51694) := X"8FC20040";
        ram_buffer(51695) := X"00000000";
        ram_buffer(51696) := X"8C430004";
        ram_buffer(51697) := X"2402FFFE";
        ram_buffer(51698) := X"00621024";
        ram_buffer(51699) := X"8FC30040";
        ram_buffer(51700) := X"00000000";
        ram_buffer(51701) := X"00621021";
        ram_buffer(51702) := X"8FC30010";
        ram_buffer(51703) := X"00000000";
        ram_buffer(51704) := X"1462000F";
        ram_buffer(51705) := X"00000000";
        ram_buffer(51706) := X"8FC20010";
        ram_buffer(51707) := X"00000000";
        ram_buffer(51708) := X"8C430004";
        ram_buffer(51709) := X"2402FFFC";
        ram_buffer(51710) := X"00621024";
        ram_buffer(51711) := X"8FC30014";
        ram_buffer(51712) := X"00000000";
        ram_buffer(51713) := X"00621021";
        ram_buffer(51714) := X"AFC20014";
        ram_buffer(51715) := X"8FC20040";
        ram_buffer(51716) := X"00000000";
        ram_buffer(51717) := X"AFC20010";
        ram_buffer(51718) := X"1000008E";
        ram_buffer(51719) := X"00000000";
        ram_buffer(51720) := X"8FC20044";
        ram_buffer(51721) := X"00000000";
        ram_buffer(51722) := X"2442FFFC";
        ram_buffer(51723) := X"AFC2006C";
        ram_buffer(51724) := X"8FC2006C";
        ram_buffer(51725) := X"00000000";
        ram_buffer(51726) := X"2C420025";
        ram_buffer(51727) := X"10400076";
        ram_buffer(51728) := X"00000000";
        ram_buffer(51729) := X"8FC20084";
        ram_buffer(51730) := X"00000000";
        ram_buffer(51731) := X"AFC20038";
        ram_buffer(51732) := X"8FC2005C";
        ram_buffer(51733) := X"00000000";
        ram_buffer(51734) := X"AFC2003C";
        ram_buffer(51735) := X"8FC2006C";
        ram_buffer(51736) := X"00000000";
        ram_buffer(51737) := X"2C420014";
        ram_buffer(51738) := X"1440004D";
        ram_buffer(51739) := X"00000000";
        ram_buffer(51740) := X"8FC2003C";
        ram_buffer(51741) := X"00000000";
        ram_buffer(51742) := X"24430004";
        ram_buffer(51743) := X"AFC3003C";
        ram_buffer(51744) := X"8FC30038";
        ram_buffer(51745) := X"00000000";
        ram_buffer(51746) := X"24640004";
        ram_buffer(51747) := X"AFC40038";
        ram_buffer(51748) := X"8C630000";
        ram_buffer(51749) := X"00000000";
        ram_buffer(51750) := X"AC430000";
        ram_buffer(51751) := X"8FC2003C";
        ram_buffer(51752) := X"00000000";
        ram_buffer(51753) := X"24430004";
        ram_buffer(51754) := X"AFC3003C";
        ram_buffer(51755) := X"8FC30038";
        ram_buffer(51756) := X"00000000";
        ram_buffer(51757) := X"24640004";
        ram_buffer(51758) := X"AFC40038";
        ram_buffer(51759) := X"8C630000";
        ram_buffer(51760) := X"00000000";
        ram_buffer(51761) := X"AC430000";
        ram_buffer(51762) := X"8FC2006C";
        ram_buffer(51763) := X"00000000";
        ram_buffer(51764) := X"2C42001C";
        ram_buffer(51765) := X"14400032";
        ram_buffer(51766) := X"00000000";
        ram_buffer(51767) := X"8FC2003C";
        ram_buffer(51768) := X"00000000";
        ram_buffer(51769) := X"24430004";
        ram_buffer(51770) := X"AFC3003C";
        ram_buffer(51771) := X"8FC30038";
        ram_buffer(51772) := X"00000000";
        ram_buffer(51773) := X"24640004";
        ram_buffer(51774) := X"AFC40038";
        ram_buffer(51775) := X"8C630000";
        ram_buffer(51776) := X"00000000";
        ram_buffer(51777) := X"AC430000";
        ram_buffer(51778) := X"8FC2003C";
        ram_buffer(51779) := X"00000000";
        ram_buffer(51780) := X"24430004";
        ram_buffer(51781) := X"AFC3003C";
        ram_buffer(51782) := X"8FC30038";
        ram_buffer(51783) := X"00000000";
        ram_buffer(51784) := X"24640004";
        ram_buffer(51785) := X"AFC40038";
        ram_buffer(51786) := X"8C630000";
        ram_buffer(51787) := X"00000000";
        ram_buffer(51788) := X"AC430000";
        ram_buffer(51789) := X"8FC2006C";
        ram_buffer(51790) := X"00000000";
        ram_buffer(51791) := X"2C420024";
        ram_buffer(51792) := X"14400017";
        ram_buffer(51793) := X"00000000";
        ram_buffer(51794) := X"8FC2003C";
        ram_buffer(51795) := X"00000000";
        ram_buffer(51796) := X"24430004";
        ram_buffer(51797) := X"AFC3003C";
        ram_buffer(51798) := X"8FC30038";
        ram_buffer(51799) := X"00000000";
        ram_buffer(51800) := X"24640004";
        ram_buffer(51801) := X"AFC40038";
        ram_buffer(51802) := X"8C630000";
        ram_buffer(51803) := X"00000000";
        ram_buffer(51804) := X"AC430000";
        ram_buffer(51805) := X"8FC2003C";
        ram_buffer(51806) := X"00000000";
        ram_buffer(51807) := X"24430004";
        ram_buffer(51808) := X"AFC3003C";
        ram_buffer(51809) := X"8FC30038";
        ram_buffer(51810) := X"00000000";
        ram_buffer(51811) := X"24640004";
        ram_buffer(51812) := X"AFC40038";
        ram_buffer(51813) := X"8C630000";
        ram_buffer(51814) := X"00000000";
        ram_buffer(51815) := X"AC430000";
        ram_buffer(51816) := X"8FC2003C";
        ram_buffer(51817) := X"00000000";
        ram_buffer(51818) := X"24430004";
        ram_buffer(51819) := X"AFC3003C";
        ram_buffer(51820) := X"8FC30038";
        ram_buffer(51821) := X"00000000";
        ram_buffer(51822) := X"24640004";
        ram_buffer(51823) := X"AFC40038";
        ram_buffer(51824) := X"8C630000";
        ram_buffer(51825) := X"00000000";
        ram_buffer(51826) := X"AC430000";
        ram_buffer(51827) := X"8FC2003C";
        ram_buffer(51828) := X"00000000";
        ram_buffer(51829) := X"24430004";
        ram_buffer(51830) := X"AFC3003C";
        ram_buffer(51831) := X"8FC30038";
        ram_buffer(51832) := X"00000000";
        ram_buffer(51833) := X"24640004";
        ram_buffer(51834) := X"AFC40038";
        ram_buffer(51835) := X"8C630000";
        ram_buffer(51836) := X"00000000";
        ram_buffer(51837) := X"AC430000";
        ram_buffer(51838) := X"8FC20038";
        ram_buffer(51839) := X"00000000";
        ram_buffer(51840) := X"8C430000";
        ram_buffer(51841) := X"8FC2003C";
        ram_buffer(51842) := X"00000000";
        ram_buffer(51843) := X"AC430000";
        ram_buffer(51844) := X"10000006";
        ram_buffer(51845) := X"00000000";
        ram_buffer(51846) := X"8FC6006C";
        ram_buffer(51847) := X"8FC50084";
        ram_buffer(51848) := X"8FC4005C";
        ram_buffer(51849) := X"0C02BCED";
        ram_buffer(51850) := X"00000000";
        ram_buffer(51851) := X"8FC50084";
        ram_buffer(51852) := X"8FC40080";
        ram_buffer(51853) := X"0C027301";
        ram_buffer(51854) := X"00000000";
        ram_buffer(51855) := X"8FC40080";
        ram_buffer(51856) := X"0C0280CD";
        ram_buffer(51857) := X"00000000";
        ram_buffer(51858) := X"8FC2005C";
        ram_buffer(51859) := X"10000053";
        ram_buffer(51860) := X"00000000";
        ram_buffer(51861) := X"8FC30014";
        ram_buffer(51862) := X"8FC20048";
        ram_buffer(51863) := X"00000000";
        ram_buffer(51864) := X"00621023";
        ram_buffer(51865) := X"AFC20070";
        ram_buffer(51866) := X"8FC20070";
        ram_buffer(51867) := X"00000000";
        ram_buffer(51868) := X"2C420010";
        ram_buffer(51869) := X"1440002C";
        ram_buffer(51870) := X"00000000";
        ram_buffer(51871) := X"8FC30010";
        ram_buffer(51872) := X"8FC20048";
        ram_buffer(51873) := X"00000000";
        ram_buffer(51874) := X"00621021";
        ram_buffer(51875) := X"AFC20074";
        ram_buffer(51876) := X"8FC20010";
        ram_buffer(51877) := X"00000000";
        ram_buffer(51878) := X"8C420004";
        ram_buffer(51879) := X"00000000";
        ram_buffer(51880) := X"30430001";
        ram_buffer(51881) := X"8FC20048";
        ram_buffer(51882) := X"00000000";
        ram_buffer(51883) := X"00621825";
        ram_buffer(51884) := X"8FC20010";
        ram_buffer(51885) := X"00000000";
        ram_buffer(51886) := X"AC430004";
        ram_buffer(51887) := X"8FC20070";
        ram_buffer(51888) := X"00000000";
        ram_buffer(51889) := X"34430001";
        ram_buffer(51890) := X"8FC20074";
        ram_buffer(51891) := X"00000000";
        ram_buffer(51892) := X"AC430004";
        ram_buffer(51893) := X"8FC30074";
        ram_buffer(51894) := X"8FC20070";
        ram_buffer(51895) := X"00000000";
        ram_buffer(51896) := X"00621021";
        ram_buffer(51897) := X"8FC40074";
        ram_buffer(51898) := X"8FC30070";
        ram_buffer(51899) := X"00000000";
        ram_buffer(51900) := X"00831821";
        ram_buffer(51901) := X"8C630004";
        ram_buffer(51902) := X"00000000";
        ram_buffer(51903) := X"34630001";
        ram_buffer(51904) := X"AC430004";
        ram_buffer(51905) := X"8FC20074";
        ram_buffer(51906) := X"00000000";
        ram_buffer(51907) := X"24420008";
        ram_buffer(51908) := X"00402821";
        ram_buffer(51909) := X"8FC40080";
        ram_buffer(51910) := X"0C027301";
        ram_buffer(51911) := X"00000000";
        ram_buffer(51912) := X"10000018";
        ram_buffer(51913) := X"00000000";
        ram_buffer(51914) := X"8FC20010";
        ram_buffer(51915) := X"00000000";
        ram_buffer(51916) := X"8C420004";
        ram_buffer(51917) := X"00000000";
        ram_buffer(51918) := X"30430001";
        ram_buffer(51919) := X"8FC20014";
        ram_buffer(51920) := X"00000000";
        ram_buffer(51921) := X"00621825";
        ram_buffer(51922) := X"8FC20010";
        ram_buffer(51923) := X"00000000";
        ram_buffer(51924) := X"AC430004";
        ram_buffer(51925) := X"8FC30010";
        ram_buffer(51926) := X"8FC20014";
        ram_buffer(51927) := X"00000000";
        ram_buffer(51928) := X"00621021";
        ram_buffer(51929) := X"8FC40010";
        ram_buffer(51930) := X"8FC30014";
        ram_buffer(51931) := X"00000000";
        ram_buffer(51932) := X"00831821";
        ram_buffer(51933) := X"8C630004";
        ram_buffer(51934) := X"00000000";
        ram_buffer(51935) := X"34630001";
        ram_buffer(51936) := X"AC430004";
        ram_buffer(51937) := X"8FC40080";
        ram_buffer(51938) := X"0C0280CD";
        ram_buffer(51939) := X"00000000";
        ram_buffer(51940) := X"8FC20010";
        ram_buffer(51941) := X"00000000";
        ram_buffer(51942) := X"24420008";
        ram_buffer(51943) := X"03C0E821";
        ram_buffer(51944) := X"8FBF007C";
        ram_buffer(51945) := X"8FBE0078";
        ram_buffer(51946) := X"27BD0080";
        ram_buffer(51947) := X"03E00008";
        ram_buffer(51948) := X"00000000";
        ram_buffer(51949) := X"27BDFFE8";
        ram_buffer(51950) := X"AFBE0014";
        ram_buffer(51951) := X"03A0F021";
        ram_buffer(51952) := X"AFC5001C";
        ram_buffer(51953) := X"AFC40018";
        ram_buffer(51954) := X"8FC3001C";
        ram_buffer(51955) := X"8FC20018";
        ram_buffer(51956) := X"AFC3000C";
        ram_buffer(51957) := X"AFC20008";
        ram_buffer(51958) := X"8FC20008";
        ram_buffer(51959) := X"00000000";
        ram_buffer(51960) := X"AFC20000";
        ram_buffer(51961) := X"8FC2000C";
        ram_buffer(51962) := X"00000000";
        ram_buffer(51963) := X"AFC20004";
        ram_buffer(51964) := X"8FC20000";
        ram_buffer(51965) := X"00000000";
        ram_buffer(51966) := X"14400005";
        ram_buffer(51967) := X"00000000";
        ram_buffer(51968) := X"8FC20004";
        ram_buffer(51969) := X"00000000";
        ram_buffer(51970) := X"10400009";
        ram_buffer(51971) := X"00000000";
        ram_buffer(51972) := X"8FC30000";
        ram_buffer(51973) := X"3C028000";
        ram_buffer(51974) := X"14620008";
        ram_buffer(51975) := X"00000000";
        ram_buffer(51976) := X"8FC20004";
        ram_buffer(51977) := X"00000000";
        ram_buffer(51978) := X"14400004";
        ram_buffer(51979) := X"00000000";
        ram_buffer(51980) := X"24020002";
        ram_buffer(51981) := X"1000003D";
        ram_buffer(51982) := X"00000000";
        ram_buffer(51983) := X"8FC30000";
        ram_buffer(51984) := X"3C020010";
        ram_buffer(51985) := X"0062102B";
        ram_buffer(51986) := X"14400006";
        ram_buffer(51987) := X"00000000";
        ram_buffer(51988) := X"8FC30000";
        ram_buffer(51989) := X"3C027FF0";
        ram_buffer(51990) := X"0062102B";
        ram_buffer(51991) := X"1440000B";
        ram_buffer(51992) := X"00000000";
        ram_buffer(51993) := X"8FC30000";
        ram_buffer(51994) := X"3C028010";
        ram_buffer(51995) := X"0062102B";
        ram_buffer(51996) := X"14400009";
        ram_buffer(51997) := X"00000000";
        ram_buffer(51998) := X"8FC30000";
        ram_buffer(51999) := X"3C02FFF0";
        ram_buffer(52000) := X"0062102B";
        ram_buffer(52001) := X"10400004";
        ram_buffer(52002) := X"00000000";
        ram_buffer(52003) := X"24020004";
        ram_buffer(52004) := X"10000026";
        ram_buffer(52005) := X"00000000";
        ram_buffer(52006) := X"8FC30000";
        ram_buffer(52007) := X"3C020010";
        ram_buffer(52008) := X"0062102B";
        ram_buffer(52009) := X"1440000A";
        ram_buffer(52010) := X"00000000";
        ram_buffer(52011) := X"8FC20000";
        ram_buffer(52012) := X"00000000";
        ram_buffer(52013) := X"04410009";
        ram_buffer(52014) := X"00000000";
        ram_buffer(52015) := X"8FC30000";
        ram_buffer(52016) := X"3C028010";
        ram_buffer(52017) := X"0062102B";
        ram_buffer(52018) := X"10400004";
        ram_buffer(52019) := X"00000000";
        ram_buffer(52020) := X"24020003";
        ram_buffer(52021) := X"10000015";
        ram_buffer(52022) := X"00000000";
        ram_buffer(52023) := X"8FC30000";
        ram_buffer(52024) := X"3C027FF0";
        ram_buffer(52025) := X"14620005";
        ram_buffer(52026) := X"00000000";
        ram_buffer(52027) := X"8FC20004";
        ram_buffer(52028) := X"00000000";
        ram_buffer(52029) := X"10400009";
        ram_buffer(52030) := X"00000000";
        ram_buffer(52031) := X"8FC30000";
        ram_buffer(52032) := X"3C02FFF0";
        ram_buffer(52033) := X"14620008";
        ram_buffer(52034) := X"00000000";
        ram_buffer(52035) := X"8FC20004";
        ram_buffer(52036) := X"00000000";
        ram_buffer(52037) := X"14400004";
        ram_buffer(52038) := X"00000000";
        ram_buffer(52039) := X"24020001";
        ram_buffer(52040) := X"10000002";
        ram_buffer(52041) := X"00000000";
        ram_buffer(52042) := X"00001021";
        ram_buffer(52043) := X"03C0E821";
        ram_buffer(52044) := X"8FBE0014";
        ram_buffer(52045) := X"27BD0018";
        ram_buffer(52046) := X"03E00008";
        ram_buffer(52047) := X"00000000";
        ram_buffer(52048) := X"27BDFFC0";
        ram_buffer(52049) := X"AFBF003C";
        ram_buffer(52050) := X"AFBE0038";
        ram_buffer(52051) := X"03A0F021";
        ram_buffer(52052) := X"AFC50044";
        ram_buffer(52053) := X"AFC40040";
        ram_buffer(52054) := X"AFC60048";
        ram_buffer(52055) := X"8FC30044";
        ram_buffer(52056) := X"8FC20040";
        ram_buffer(52057) := X"AFC30024";
        ram_buffer(52058) := X"AFC20020";
        ram_buffer(52059) := X"8FC20020";
        ram_buffer(52060) := X"00000000";
        ram_buffer(52061) := X"AFC20010";
        ram_buffer(52062) := X"8FC20024";
        ram_buffer(52063) := X"00000000";
        ram_buffer(52064) := X"AFC20018";
        ram_buffer(52065) := X"8FC30010";
        ram_buffer(52066) := X"3C027FFF";
        ram_buffer(52067) := X"3442FFFF";
        ram_buffer(52068) := X"00621024";
        ram_buffer(52069) := X"AFC20014";
        ram_buffer(52070) := X"8FC20048";
        ram_buffer(52071) := X"00000000";
        ram_buffer(52072) := X"AC400000";
        ram_buffer(52073) := X"8FC30014";
        ram_buffer(52074) := X"3C027FF0";
        ram_buffer(52075) := X"0062102A";
        ram_buffer(52076) := X"10400007";
        ram_buffer(52077) := X"00000000";
        ram_buffer(52078) := X"8FC30014";
        ram_buffer(52079) := X"8FC20018";
        ram_buffer(52080) := X"00000000";
        ram_buffer(52081) := X"00621025";
        ram_buffer(52082) := X"14400005";
        ram_buffer(52083) := X"00000000";
        ram_buffer(52084) := X"8FC30044";
        ram_buffer(52085) := X"8FC20040";
        ram_buffer(52086) := X"1000003E";
        ram_buffer(52087) := X"00000000";
        ram_buffer(52088) := X"8FC30014";
        ram_buffer(52089) := X"3C020010";
        ram_buffer(52090) := X"0062102A";
        ram_buffer(52091) := X"1040001A";
        ram_buffer(52092) := X"00000000";
        ram_buffer(52093) := X"8F83814C";
        ram_buffer(52094) := X"8F828148";
        ram_buffer(52095) := X"00603821";
        ram_buffer(52096) := X"00403021";
        ram_buffer(52097) := X"8FC50044";
        ram_buffer(52098) := X"8FC40040";
        ram_buffer(52099) := X"0C03174A";
        ram_buffer(52100) := X"00000000";
        ram_buffer(52101) := X"AFC30044";
        ram_buffer(52102) := X"AFC20040";
        ram_buffer(52103) := X"8FC30044";
        ram_buffer(52104) := X"8FC20040";
        ram_buffer(52105) := X"AFC3002C";
        ram_buffer(52106) := X"AFC20028";
        ram_buffer(52107) := X"8FC20028";
        ram_buffer(52108) := X"00000000";
        ram_buffer(52109) := X"AFC20010";
        ram_buffer(52110) := X"8FC30010";
        ram_buffer(52111) := X"3C027FFF";
        ram_buffer(52112) := X"3442FFFF";
        ram_buffer(52113) := X"00621024";
        ram_buffer(52114) := X"AFC20014";
        ram_buffer(52115) := X"8FC20048";
        ram_buffer(52116) := X"2403FFCA";
        ram_buffer(52117) := X"AC430000";
        ram_buffer(52118) := X"8FC20048";
        ram_buffer(52119) := X"00000000";
        ram_buffer(52120) := X"8C430000";
        ram_buffer(52121) := X"8FC20014";
        ram_buffer(52122) := X"00000000";
        ram_buffer(52123) := X"00021503";
        ram_buffer(52124) := X"2442FC02";
        ram_buffer(52125) := X"00621821";
        ram_buffer(52126) := X"8FC20048";
        ram_buffer(52127) := X"00000000";
        ram_buffer(52128) := X"AC430000";
        ram_buffer(52129) := X"8FC30010";
        ram_buffer(52130) := X"3C02800F";
        ram_buffer(52131) := X"3442FFFF";
        ram_buffer(52132) := X"00621824";
        ram_buffer(52133) := X"3C023FE0";
        ram_buffer(52134) := X"00621025";
        ram_buffer(52135) := X"AFC20010";
        ram_buffer(52136) := X"8FC30044";
        ram_buffer(52137) := X"8FC20040";
        ram_buffer(52138) := X"AFC30034";
        ram_buffer(52139) := X"AFC20030";
        ram_buffer(52140) := X"8FC20010";
        ram_buffer(52141) := X"00000000";
        ram_buffer(52142) := X"AFC20030";
        ram_buffer(52143) := X"8FC30034";
        ram_buffer(52144) := X"8FC20030";
        ram_buffer(52145) := X"AFC30044";
        ram_buffer(52146) := X"AFC20040";
        ram_buffer(52147) := X"8FC30044";
        ram_buffer(52148) := X"8FC20040";
        ram_buffer(52149) := X"03C0E821";
        ram_buffer(52150) := X"8FBF003C";
        ram_buffer(52151) := X"8FBE0038";
        ram_buffer(52152) := X"27BD0040";
        ram_buffer(52153) := X"03E00008";
        ram_buffer(52154) := X"00000000";
        ram_buffer(52155) := X"27BDFFF0";
        ram_buffer(52156) := X"AFBE000C";
        ram_buffer(52157) := X"AFB20008";
        ram_buffer(52158) := X"AFB10004";
        ram_buffer(52159) := X"AFB00000";
        ram_buffer(52160) := X"03A0F021";
        ram_buffer(52161) := X"00801821";
        ram_buffer(52162) := X"00A01021";
        ram_buffer(52163) := X"00402021";
        ram_buffer(52164) := X"24820001";
        ram_buffer(52165) := X"90840000";
        ram_buffer(52166) := X"00000000";
        ram_buffer(52167) := X"00808821";
        ram_buffer(52168) := X"2404005E";
        ram_buffer(52169) := X"16240009";
        ram_buffer(52170) := X"00000000";
        ram_buffer(52171) := X"24120001";
        ram_buffer(52172) := X"00402021";
        ram_buffer(52173) := X"24820001";
        ram_buffer(52174) := X"90840000";
        ram_buffer(52175) := X"00000000";
        ram_buffer(52176) := X"00808821";
        ram_buffer(52177) := X"10000002";
        ram_buffer(52178) := X"00000000";
        ram_buffer(52179) := X"00009021";
        ram_buffer(52180) := X"00008021";
        ram_buffer(52181) := X"10000007";
        ram_buffer(52182) := X"00000000";
        ram_buffer(52183) := X"02002021";
        ram_buffer(52184) := X"00642021";
        ram_buffer(52185) := X"00122E00";
        ram_buffer(52186) := X"00052E03";
        ram_buffer(52187) := X"A0850000";
        ram_buffer(52188) := X"26100001";
        ram_buffer(52189) := X"2A040100";
        ram_buffer(52190) := X"1480FFF8";
        ram_buffer(52191) := X"00000000";
        ram_buffer(52192) := X"16200004";
        ram_buffer(52193) := X"00000000";
        ram_buffer(52194) := X"2442FFFF";
        ram_buffer(52195) := X"10000036";
        ram_buffer(52196) := X"00000000";
        ram_buffer(52197) := X"24040001";
        ram_buffer(52198) := X"00929023";
        ram_buffer(52199) := X"02202021";
        ram_buffer(52200) := X"00642021";
        ram_buffer(52201) := X"00122E00";
        ram_buffer(52202) := X"00052E03";
        ram_buffer(52203) := X"A0850000";
        ram_buffer(52204) := X"00402021";
        ram_buffer(52205) := X"24820001";
        ram_buffer(52206) := X"90840000";
        ram_buffer(52207) := X"00000000";
        ram_buffer(52208) := X"00808021";
        ram_buffer(52209) := X"2404002D";
        ram_buffer(52210) := X"12040009";
        ram_buffer(52211) := X"00000000";
        ram_buffer(52212) := X"2404005D";
        ram_buffer(52213) := X"1204001E";
        ram_buffer(52214) := X"00000000";
        ram_buffer(52215) := X"1600001E";
        ram_buffer(52216) := X"00000000";
        ram_buffer(52217) := X"2442FFFF";
        ram_buffer(52218) := X"1000001F";
        ram_buffer(52219) := X"00000000";
        ram_buffer(52220) := X"90440000";
        ram_buffer(52221) := X"00000000";
        ram_buffer(52222) := X"00808021";
        ram_buffer(52223) := X"2404005D";
        ram_buffer(52224) := X"12040004";
        ram_buffer(52225) := X"00000000";
        ram_buffer(52226) := X"0211202A";
        ram_buffer(52227) := X"10800004";
        ram_buffer(52228) := X"00000000";
        ram_buffer(52229) := X"2411002D";
        ram_buffer(52230) := X"10000011";
        ram_buffer(52231) := X"00000000";
        ram_buffer(52232) := X"24420001";
        ram_buffer(52233) := X"26310001";
        ram_buffer(52234) := X"02202021";
        ram_buffer(52235) := X"00642021";
        ram_buffer(52236) := X"00122E00";
        ram_buffer(52237) := X"00052E03";
        ram_buffer(52238) := X"A0850000";
        ram_buffer(52239) := X"0230202A";
        ram_buffer(52240) := X"1480FFF8";
        ram_buffer(52241) := X"00000000";
        ram_buffer(52242) := X"1000FFD9";
        ram_buffer(52243) := X"00000000";
        ram_buffer(52244) := X"10000005";
        ram_buffer(52245) := X"00000000";
        ram_buffer(52246) := X"02008821";
        ram_buffer(52247) := X"00000000";
        ram_buffer(52248) := X"1000FFCE";
        ram_buffer(52249) := X"00000000";
        ram_buffer(52250) := X"03C0E821";
        ram_buffer(52251) := X"8FBE000C";
        ram_buffer(52252) := X"8FB20008";
        ram_buffer(52253) := X"8FB10004";
        ram_buffer(52254) := X"8FB00000";
        ram_buffer(52255) := X"27BD0010";
        ram_buffer(52256) := X"03E00008";
        ram_buffer(52257) := X"00000000";
        ram_buffer(52258) := X"27BDFFF0";
        ram_buffer(52259) := X"AFBE000C";
        ram_buffer(52260) := X"03A0F021";
        ram_buffer(52261) := X"AFC40010";
        ram_buffer(52262) := X"8F828150";
        ram_buffer(52263) := X"00000000";
        ram_buffer(52264) := X"AFC20000";
        ram_buffer(52265) := X"8FC20000";
        ram_buffer(52266) := X"03C0E821";
        ram_buffer(52267) := X"8FBE000C";
        ram_buffer(52268) := X"27BD0010";
        ram_buffer(52269) := X"03E00008";
        ram_buffer(52270) := X"00000000";
        ram_buffer(52271) := X"00854025";
        ram_buffer(52272) := X"31080003";
        ram_buffer(52273) := X"1500005E";
        ram_buffer(52274) := X"3C180101";
        ram_buffer(52275) := X"37180101";
        ram_buffer(52276) := X"3C197F7F";
        ram_buffer(52277) := X"37397F7F";
        ram_buffer(52278) := X"8C820000";
        ram_buffer(52279) := X"8CA30000";
        ram_buffer(52280) := X"00584023";
        ram_buffer(52281) := X"14430040";
        ram_buffer(52282) := X"00594827";
        ram_buffer(52283) := X"01094024";
        ram_buffer(52284) := X"1500003B";
        ram_buffer(52285) := X"00000000";
        ram_buffer(52286) := X"8C820004";
        ram_buffer(52287) := X"8CA30004";
        ram_buffer(52288) := X"00584023";
        ram_buffer(52289) := X"14430038";
        ram_buffer(52290) := X"00594827";
        ram_buffer(52291) := X"01094024";
        ram_buffer(52292) := X"15000033";
        ram_buffer(52293) := X"00000000";
        ram_buffer(52294) := X"8C820008";
        ram_buffer(52295) := X"8CA30008";
        ram_buffer(52296) := X"00584023";
        ram_buffer(52297) := X"14430030";
        ram_buffer(52298) := X"00594827";
        ram_buffer(52299) := X"01094024";
        ram_buffer(52300) := X"1500002B";
        ram_buffer(52301) := X"00000000";
        ram_buffer(52302) := X"8C82000C";
        ram_buffer(52303) := X"8CA3000C";
        ram_buffer(52304) := X"00584023";
        ram_buffer(52305) := X"14430028";
        ram_buffer(52306) := X"00594827";
        ram_buffer(52307) := X"01094024";
        ram_buffer(52308) := X"15000023";
        ram_buffer(52309) := X"00000000";
        ram_buffer(52310) := X"8C820010";
        ram_buffer(52311) := X"8CA30010";
        ram_buffer(52312) := X"00584023";
        ram_buffer(52313) := X"14430020";
        ram_buffer(52314) := X"00594827";
        ram_buffer(52315) := X"01094024";
        ram_buffer(52316) := X"1500001B";
        ram_buffer(52317) := X"00000000";
        ram_buffer(52318) := X"8C820014";
        ram_buffer(52319) := X"8CA30014";
        ram_buffer(52320) := X"00584023";
        ram_buffer(52321) := X"14430018";
        ram_buffer(52322) := X"00594827";
        ram_buffer(52323) := X"01094024";
        ram_buffer(52324) := X"15000013";
        ram_buffer(52325) := X"00000000";
        ram_buffer(52326) := X"8C820018";
        ram_buffer(52327) := X"8CA30018";
        ram_buffer(52328) := X"00584023";
        ram_buffer(52329) := X"14430010";
        ram_buffer(52330) := X"00594827";
        ram_buffer(52331) := X"01094024";
        ram_buffer(52332) := X"1500000B";
        ram_buffer(52333) := X"00000000";
        ram_buffer(52334) := X"8C82001C";
        ram_buffer(52335) := X"8CA3001C";
        ram_buffer(52336) := X"00584023";
        ram_buffer(52337) := X"14430008";
        ram_buffer(52338) := X"00594827";
        ram_buffer(52339) := X"01094024";
        ram_buffer(52340) := X"15000003";
        ram_buffer(52341) := X"24840020";
        ram_buffer(52342) := X"1000FFBF";
        ram_buffer(52343) := X"24A50020";
        ram_buffer(52344) := X"03E00008";
        ram_buffer(52345) := X"00001021";
        ram_buffer(52346) := X"00024602";
        ram_buffer(52347) := X"11000012";
        ram_buffer(52348) := X"00034E02";
        ram_buffer(52349) := X"15090010";
        ram_buffer(52350) := X"0002C402";
        ram_buffer(52351) := X"0003CC02";
        ram_buffer(52352) := X"331800FF";
        ram_buffer(52353) := X"1300000A";
        ram_buffer(52354) := X"333900FF";
        ram_buffer(52355) := X"17190008";
        ram_buffer(52356) := X"00024202";
        ram_buffer(52357) := X"00034A02";
        ram_buffer(52358) := X"310800FF";
        ram_buffer(52359) := X"11000006";
        ram_buffer(52360) := X"312900FF";
        ram_buffer(52361) := X"15090004";
        ram_buffer(52362) := X"305800FF";
        ram_buffer(52363) := X"307900FF";
        ram_buffer(52364) := X"03E00008";
        ram_buffer(52365) := X"03191023";
        ram_buffer(52366) := X"03E00008";
        ram_buffer(52367) := X"01091023";
        ram_buffer(52368) := X"90820000";
        ram_buffer(52369) := X"90A30000";
        ram_buffer(52370) := X"10400028";
        ram_buffer(52371) := X"00000000";
        ram_buffer(52372) := X"14430026";
        ram_buffer(52373) := X"90980001";
        ram_buffer(52374) := X"90B90001";
        ram_buffer(52375) := X"13000025";
        ram_buffer(52376) := X"00000000";
        ram_buffer(52377) := X"17190023";
        ram_buffer(52378) := X"90820002";
        ram_buffer(52379) := X"90A30002";
        ram_buffer(52380) := X"1040001E";
        ram_buffer(52381) := X"00000000";
        ram_buffer(52382) := X"1443001C";
        ram_buffer(52383) := X"90980003";
        ram_buffer(52384) := X"90B90003";
        ram_buffer(52385) := X"1300001B";
        ram_buffer(52386) := X"00000000";
        ram_buffer(52387) := X"17190019";
        ram_buffer(52388) := X"90820004";
        ram_buffer(52389) := X"90A30004";
        ram_buffer(52390) := X"10400014";
        ram_buffer(52391) := X"00000000";
        ram_buffer(52392) := X"14430012";
        ram_buffer(52393) := X"90980005";
        ram_buffer(52394) := X"90B90005";
        ram_buffer(52395) := X"13000011";
        ram_buffer(52396) := X"00000000";
        ram_buffer(52397) := X"1719000F";
        ram_buffer(52398) := X"90820006";
        ram_buffer(52399) := X"90A30006";
        ram_buffer(52400) := X"1040000A";
        ram_buffer(52401) := X"00000000";
        ram_buffer(52402) := X"14430008";
        ram_buffer(52403) := X"90980007";
        ram_buffer(52404) := X"90B90007";
        ram_buffer(52405) := X"13000007";
        ram_buffer(52406) := X"00000000";
        ram_buffer(52407) := X"17190005";
        ram_buffer(52408) := X"24840008";
        ram_buffer(52409) := X"1000FFD6";
        ram_buffer(52410) := X"24A50008";
        ram_buffer(52411) := X"03E00008";
        ram_buffer(52412) := X"00431023";
        ram_buffer(52413) := X"03E00008";
        ram_buffer(52414) := X"03191023";
        ram_buffer(52415) := X"27BDFFD0";
        ram_buffer(52416) := X"AFBE002C";
        ram_buffer(52417) := X"03A0F021";
        ram_buffer(52418) := X"AFC40030";
        ram_buffer(52419) := X"AFC50034";
        ram_buffer(52420) := X"AFC60038";
        ram_buffer(52421) := X"8FC20030";
        ram_buffer(52422) := X"00000000";
        ram_buffer(52423) := X"AFC20000";
        ram_buffer(52424) := X"8FC20034";
        ram_buffer(52425) := X"00000000";
        ram_buffer(52426) := X"AFC20004";
        ram_buffer(52427) := X"1000002C";
        ram_buffer(52428) := X"00000000";
        ram_buffer(52429) := X"8FC20000";
        ram_buffer(52430) := X"00000000";
        ram_buffer(52431) := X"24430001";
        ram_buffer(52432) := X"AFC30000";
        ram_buffer(52433) := X"8FC30004";
        ram_buffer(52434) := X"00000000";
        ram_buffer(52435) := X"24640001";
        ram_buffer(52436) := X"AFC40004";
        ram_buffer(52437) := X"90630000";
        ram_buffer(52438) := X"00000000";
        ram_buffer(52439) := X"AFC30008";
        ram_buffer(52440) := X"8FC30008";
        ram_buffer(52441) := X"00000000";
        ram_buffer(52442) := X"306300FF";
        ram_buffer(52443) := X"A0430000";
        ram_buffer(52444) := X"8FC20038";
        ram_buffer(52445) := X"00000000";
        ram_buffer(52446) := X"2442FFFF";
        ram_buffer(52447) := X"AFC20038";
        ram_buffer(52448) := X"8FC20008";
        ram_buffer(52449) := X"00000000";
        ram_buffer(52450) := X"14400015";
        ram_buffer(52451) := X"00000000";
        ram_buffer(52452) := X"8FC30000";
        ram_buffer(52453) := X"8FC20038";
        ram_buffer(52454) := X"00000000";
        ram_buffer(52455) := X"00621021";
        ram_buffer(52456) := X"AFC2000C";
        ram_buffer(52457) := X"10000006";
        ram_buffer(52458) := X"00000000";
        ram_buffer(52459) := X"8FC20000";
        ram_buffer(52460) := X"00000000";
        ram_buffer(52461) := X"24430001";
        ram_buffer(52462) := X"AFC30000";
        ram_buffer(52463) := X"A0400000";
        ram_buffer(52464) := X"8FC30000";
        ram_buffer(52465) := X"8FC2000C";
        ram_buffer(52466) := X"00000000";
        ram_buffer(52467) := X"1462FFF7";
        ram_buffer(52468) := X"00000000";
        ram_buffer(52469) := X"8FC20030";
        ram_buffer(52470) := X"10000139";
        ram_buffer(52471) := X"00000000";
        ram_buffer(52472) := X"8FC20004";
        ram_buffer(52473) := X"00000000";
        ram_buffer(52474) := X"30420003";
        ram_buffer(52475) := X"10400005";
        ram_buffer(52476) := X"00000000";
        ram_buffer(52477) := X"8FC20038";
        ram_buffer(52478) := X"00000000";
        ram_buffer(52479) := X"1440FFCD";
        ram_buffer(52480) := X"00000000";
        ram_buffer(52481) := X"8FC20038";
        ram_buffer(52482) := X"00000000";
        ram_buffer(52483) := X"2C420004";
        ram_buffer(52484) := X"38420001";
        ram_buffer(52485) := X"304200FF";
        ram_buffer(52486) := X"1040005F";
        ram_buffer(52487) := X"00000000";
        ram_buffer(52488) := X"8FC20038";
        ram_buffer(52489) := X"00000000";
        ram_buffer(52490) := X"30420003";
        ram_buffer(52491) := X"AFC20010";
        ram_buffer(52492) := X"8FC20010";
        ram_buffer(52493) := X"8FC30038";
        ram_buffer(52494) := X"00000000";
        ram_buffer(52495) := X"00621023";
        ram_buffer(52496) := X"AFC20038";
        ram_buffer(52497) := X"8FC20004";
        ram_buffer(52498) := X"00000000";
        ram_buffer(52499) := X"90420000";
        ram_buffer(52500) := X"00000000";
        ram_buffer(52501) := X"AFC20014";
        ram_buffer(52502) := X"8FC20004";
        ram_buffer(52503) := X"00000000";
        ram_buffer(52504) := X"24420001";
        ram_buffer(52505) := X"90420000";
        ram_buffer(52506) := X"00000000";
        ram_buffer(52507) := X"AFC20018";
        ram_buffer(52508) := X"8FC20004";
        ram_buffer(52509) := X"00000000";
        ram_buffer(52510) := X"24420002";
        ram_buffer(52511) := X"90420000";
        ram_buffer(52512) := X"00000000";
        ram_buffer(52513) := X"AFC2001C";
        ram_buffer(52514) := X"8FC20004";
        ram_buffer(52515) := X"00000000";
        ram_buffer(52516) := X"24420003";
        ram_buffer(52517) := X"90420000";
        ram_buffer(52518) := X"00000000";
        ram_buffer(52519) := X"AFC20020";
        ram_buffer(52520) := X"8FC20004";
        ram_buffer(52521) := X"00000000";
        ram_buffer(52522) := X"24420004";
        ram_buffer(52523) := X"AFC20004";
        ram_buffer(52524) := X"8FC20038";
        ram_buffer(52525) := X"00000000";
        ram_buffer(52526) := X"2442FFFC";
        ram_buffer(52527) := X"AFC20038";
        ram_buffer(52528) := X"8FC20014";
        ram_buffer(52529) := X"00000000";
        ram_buffer(52530) := X"304300FF";
        ram_buffer(52531) := X"8FC20000";
        ram_buffer(52532) := X"00000000";
        ram_buffer(52533) := X"A0430000";
        ram_buffer(52534) := X"8FC20014";
        ram_buffer(52535) := X"00000000";
        ram_buffer(52536) := X"1040005D";
        ram_buffer(52537) := X"00000000";
        ram_buffer(52538) := X"8FC20000";
        ram_buffer(52539) := X"00000000";
        ram_buffer(52540) := X"24420001";
        ram_buffer(52541) := X"8FC30018";
        ram_buffer(52542) := X"00000000";
        ram_buffer(52543) := X"306300FF";
        ram_buffer(52544) := X"A0430000";
        ram_buffer(52545) := X"8FC20018";
        ram_buffer(52546) := X"00000000";
        ram_buffer(52547) := X"1040005D";
        ram_buffer(52548) := X"00000000";
        ram_buffer(52549) := X"8FC20000";
        ram_buffer(52550) := X"00000000";
        ram_buffer(52551) := X"24420002";
        ram_buffer(52552) := X"8FC3001C";
        ram_buffer(52553) := X"00000000";
        ram_buffer(52554) := X"306300FF";
        ram_buffer(52555) := X"A0430000";
        ram_buffer(52556) := X"8FC2001C";
        ram_buffer(52557) := X"00000000";
        ram_buffer(52558) := X"1040005D";
        ram_buffer(52559) := X"00000000";
        ram_buffer(52560) := X"8FC20000";
        ram_buffer(52561) := X"00000000";
        ram_buffer(52562) := X"24420003";
        ram_buffer(52563) := X"8FC30020";
        ram_buffer(52564) := X"00000000";
        ram_buffer(52565) := X"306300FF";
        ram_buffer(52566) := X"A0430000";
        ram_buffer(52567) := X"8FC20020";
        ram_buffer(52568) := X"00000000";
        ram_buffer(52569) := X"1040005D";
        ram_buffer(52570) := X"00000000";
        ram_buffer(52571) := X"8FC20000";
        ram_buffer(52572) := X"00000000";
        ram_buffer(52573) := X"24420004";
        ram_buffer(52574) := X"AFC20000";
        ram_buffer(52575) := X"8FC20038";
        ram_buffer(52576) := X"00000000";
        ram_buffer(52577) := X"1440FFAF";
        ram_buffer(52578) := X"00000000";
        ram_buffer(52579) := X"8FC20010";
        ram_buffer(52580) := X"00000000";
        ram_buffer(52581) := X"AFC20038";
        ram_buffer(52582) := X"8FC30000";
        ram_buffer(52583) := X"8FC20038";
        ram_buffer(52584) := X"00000000";
        ram_buffer(52585) := X"00621021";
        ram_buffer(52586) := X"AFC2000C";
        ram_buffer(52587) := X"10000022";
        ram_buffer(52588) := X"00000000";
        ram_buffer(52589) := X"8FC20000";
        ram_buffer(52590) := X"00000000";
        ram_buffer(52591) := X"24430001";
        ram_buffer(52592) := X"AFC30000";
        ram_buffer(52593) := X"8FC30004";
        ram_buffer(52594) := X"00000000";
        ram_buffer(52595) := X"24640001";
        ram_buffer(52596) := X"AFC40004";
        ram_buffer(52597) := X"90630000";
        ram_buffer(52598) := X"00000000";
        ram_buffer(52599) := X"AFC30008";
        ram_buffer(52600) := X"8FC30008";
        ram_buffer(52601) := X"00000000";
        ram_buffer(52602) := X"306300FF";
        ram_buffer(52603) := X"A0430000";
        ram_buffer(52604) := X"8FC20008";
        ram_buffer(52605) := X"00000000";
        ram_buffer(52606) := X"1440000F";
        ram_buffer(52607) := X"00000000";
        ram_buffer(52608) := X"10000006";
        ram_buffer(52609) := X"00000000";
        ram_buffer(52610) := X"8FC20000";
        ram_buffer(52611) := X"00000000";
        ram_buffer(52612) := X"24430001";
        ram_buffer(52613) := X"AFC30000";
        ram_buffer(52614) := X"A0400000";
        ram_buffer(52615) := X"8FC30000";
        ram_buffer(52616) := X"8FC2000C";
        ram_buffer(52617) := X"00000000";
        ram_buffer(52618) := X"1462FFF7";
        ram_buffer(52619) := X"00000000";
        ram_buffer(52620) := X"10000006";
        ram_buffer(52621) := X"00000000";
        ram_buffer(52622) := X"8FC30000";
        ram_buffer(52623) := X"8FC2000C";
        ram_buffer(52624) := X"00000000";
        ram_buffer(52625) := X"1462FFDB";
        ram_buffer(52626) := X"00000000";
        ram_buffer(52627) := X"8FC20030";
        ram_buffer(52628) := X"1000009B";
        ram_buffer(52629) := X"00000000";
        ram_buffer(52630) := X"00000000";
        ram_buffer(52631) := X"8FC20038";
        ram_buffer(52632) := X"00000000";
        ram_buffer(52633) := X"24420001";
        ram_buffer(52634) := X"AFC20038";
        ram_buffer(52635) := X"8FC20000";
        ram_buffer(52636) := X"00000000";
        ram_buffer(52637) := X"2442FFFF";
        ram_buffer(52638) := X"AFC20000";
        ram_buffer(52639) := X"10000002";
        ram_buffer(52640) := X"00000000";
        ram_buffer(52641) := X"00000000";
        ram_buffer(52642) := X"8FC20038";
        ram_buffer(52643) := X"00000000";
        ram_buffer(52644) := X"24420001";
        ram_buffer(52645) := X"AFC20038";
        ram_buffer(52646) := X"8FC20000";
        ram_buffer(52647) := X"00000000";
        ram_buffer(52648) := X"2442FFFF";
        ram_buffer(52649) := X"AFC20000";
        ram_buffer(52650) := X"10000002";
        ram_buffer(52651) := X"00000000";
        ram_buffer(52652) := X"00000000";
        ram_buffer(52653) := X"8FC20038";
        ram_buffer(52654) := X"00000000";
        ram_buffer(52655) := X"24420001";
        ram_buffer(52656) := X"AFC20038";
        ram_buffer(52657) := X"8FC20000";
        ram_buffer(52658) := X"00000000";
        ram_buffer(52659) := X"2442FFFF";
        ram_buffer(52660) := X"AFC20000";
        ram_buffer(52661) := X"10000002";
        ram_buffer(52662) := X"00000000";
        ram_buffer(52663) := X"00000000";
        ram_buffer(52664) := X"8FC20010";
        ram_buffer(52665) := X"8FC30038";
        ram_buffer(52666) := X"00000000";
        ram_buffer(52667) := X"00621021";
        ram_buffer(52668) := X"AFC20038";
        ram_buffer(52669) := X"8FC20000";
        ram_buffer(52670) := X"00000000";
        ram_buffer(52671) := X"24420004";
        ram_buffer(52672) := X"AFC20000";
        ram_buffer(52673) := X"1000000A";
        ram_buffer(52674) := X"00000000";
        ram_buffer(52675) := X"8FC20038";
        ram_buffer(52676) := X"00000000";
        ram_buffer(52677) := X"2442FFFF";
        ram_buffer(52678) := X"AFC20038";
        ram_buffer(52679) := X"8FC20000";
        ram_buffer(52680) := X"00000000";
        ram_buffer(52681) := X"24430001";
        ram_buffer(52682) := X"AFC30000";
        ram_buffer(52683) := X"A0400000";
        ram_buffer(52684) := X"8FC20038";
        ram_buffer(52685) := X"00000000";
        ram_buffer(52686) := X"10400020";
        ram_buffer(52687) := X"00000000";
        ram_buffer(52688) := X"8FC20000";
        ram_buffer(52689) := X"00000000";
        ram_buffer(52690) := X"30420003";
        ram_buffer(52691) := X"1440FFEF";
        ram_buffer(52692) := X"00000000";
        ram_buffer(52693) := X"10000019";
        ram_buffer(52694) := X"00000000";
        ram_buffer(52695) := X"8FC20038";
        ram_buffer(52696) := X"00000000";
        ram_buffer(52697) := X"2442FFF0";
        ram_buffer(52698) := X"AFC20038";
        ram_buffer(52699) := X"8FC20000";
        ram_buffer(52700) := X"00000000";
        ram_buffer(52701) := X"24420010";
        ram_buffer(52702) := X"AFC20000";
        ram_buffer(52703) := X"8FC20000";
        ram_buffer(52704) := X"00000000";
        ram_buffer(52705) := X"2442FFF0";
        ram_buffer(52706) := X"AC400000";
        ram_buffer(52707) := X"8FC20000";
        ram_buffer(52708) := X"00000000";
        ram_buffer(52709) := X"2442FFF4";
        ram_buffer(52710) := X"AC400000";
        ram_buffer(52711) := X"8FC20000";
        ram_buffer(52712) := X"00000000";
        ram_buffer(52713) := X"2442FFF8";
        ram_buffer(52714) := X"AC400000";
        ram_buffer(52715) := X"8FC20000";
        ram_buffer(52716) := X"00000000";
        ram_buffer(52717) := X"2442FFFC";
        ram_buffer(52718) := X"AC400000";
        ram_buffer(52719) := X"8FC20038";
        ram_buffer(52720) := X"00000000";
        ram_buffer(52721) := X"2C420010";
        ram_buffer(52722) := X"1040FFE4";
        ram_buffer(52723) := X"00000000";
        ram_buffer(52724) := X"8FC20038";
        ram_buffer(52725) := X"00000000";
        ram_buffer(52726) := X"2C420008";
        ram_buffer(52727) := X"14400010";
        ram_buffer(52728) := X"00000000";
        ram_buffer(52729) := X"8FC20038";
        ram_buffer(52730) := X"00000000";
        ram_buffer(52731) := X"2442FFF8";
        ram_buffer(52732) := X"AFC20038";
        ram_buffer(52733) := X"8FC20000";
        ram_buffer(52734) := X"00000000";
        ram_buffer(52735) := X"AC400000";
        ram_buffer(52736) := X"8FC20000";
        ram_buffer(52737) := X"00000000";
        ram_buffer(52738) := X"24420004";
        ram_buffer(52739) := X"AC400000";
        ram_buffer(52740) := X"8FC20000";
        ram_buffer(52741) := X"00000000";
        ram_buffer(52742) := X"24420008";
        ram_buffer(52743) := X"AFC20000";
        ram_buffer(52744) := X"8FC20038";
        ram_buffer(52745) := X"00000000";
        ram_buffer(52746) := X"2C420004";
        ram_buffer(52747) := X"1440000C";
        ram_buffer(52748) := X"00000000";
        ram_buffer(52749) := X"8FC20038";
        ram_buffer(52750) := X"00000000";
        ram_buffer(52751) := X"2442FFFC";
        ram_buffer(52752) := X"AFC20038";
        ram_buffer(52753) := X"8FC20000";
        ram_buffer(52754) := X"00000000";
        ram_buffer(52755) := X"AC400000";
        ram_buffer(52756) := X"8FC20000";
        ram_buffer(52757) := X"00000000";
        ram_buffer(52758) := X"24420004";
        ram_buffer(52759) := X"AFC20000";
        ram_buffer(52760) := X"8FC20038";
        ram_buffer(52761) := X"00000000";
        ram_buffer(52762) := X"2C420002";
        ram_buffer(52763) := X"1440000C";
        ram_buffer(52764) := X"00000000";
        ram_buffer(52765) := X"8FC20038";
        ram_buffer(52766) := X"00000000";
        ram_buffer(52767) := X"2442FFFE";
        ram_buffer(52768) := X"AFC20038";
        ram_buffer(52769) := X"8FC20000";
        ram_buffer(52770) := X"00000000";
        ram_buffer(52771) := X"A4400000";
        ram_buffer(52772) := X"8FC20000";
        ram_buffer(52773) := X"00000000";
        ram_buffer(52774) := X"24420002";
        ram_buffer(52775) := X"AFC20000";
        ram_buffer(52776) := X"8FC20038";
        ram_buffer(52777) := X"00000000";
        ram_buffer(52778) := X"10400004";
        ram_buffer(52779) := X"00000000";
        ram_buffer(52780) := X"8FC20000";
        ram_buffer(52781) := X"00000000";
        ram_buffer(52782) := X"A0400000";
        ram_buffer(52783) := X"8FC20030";
        ram_buffer(52784) := X"03C0E821";
        ram_buffer(52785) := X"8FBE002C";
        ram_buffer(52786) := X"27BD0030";
        ram_buffer(52787) := X"03E00008";
        ram_buffer(52788) := X"00000000";
        ram_buffer(52789) := X"27BDFFD0";
        ram_buffer(52790) := X"AFBF002C";
        ram_buffer(52791) := X"AFBE0028";
        ram_buffer(52792) := X"03A0F021";
        ram_buffer(52793) := X"AFC50034";
        ram_buffer(52794) := X"AFC40030";
        ram_buffer(52795) := X"AFC60038";
        ram_buffer(52796) := X"8FC30034";
        ram_buffer(52797) := X"8FC20030";
        ram_buffer(52798) := X"00602821";
        ram_buffer(52799) := X"00402021";
        ram_buffer(52800) := X"0C02C3B7";
        ram_buffer(52801) := X"00000000";
        ram_buffer(52802) := X"AFC30014";
        ram_buffer(52803) := X"AFC20010";
        ram_buffer(52804) := X"8FC20038";
        ram_buffer(52805) := X"00000000";
        ram_buffer(52806) := X"1040000C";
        ram_buffer(52807) := X"00000000";
        ram_buffer(52808) := X"8FC30030";
        ram_buffer(52809) := X"3C027FF0";
        ram_buffer(52810) := X"00621024";
        ram_buffer(52811) := X"00021502";
        ram_buffer(52812) := X"2403006B";
        ram_buffer(52813) := X"00621023";
        ram_buffer(52814) := X"AFC20018";
        ram_buffer(52815) := X"8FC20018";
        ram_buffer(52816) := X"00000000";
        ram_buffer(52817) := X"1C400005";
        ram_buffer(52818) := X"00000000";
        ram_buffer(52819) := X"8FC30014";
        ram_buffer(52820) := X"8FC20010";
        ram_buffer(52821) := X"10000011";
        ram_buffer(52822) := X"00000000";
        ram_buffer(52823) := X"8FC20018";
        ram_buffer(52824) := X"00000000";
        ram_buffer(52825) := X"00021500";
        ram_buffer(52826) := X"00401821";
        ram_buffer(52827) := X"3C023FF0";
        ram_buffer(52828) := X"00621021";
        ram_buffer(52829) := X"AFC20020";
        ram_buffer(52830) := X"AFC00024";
        ram_buffer(52831) := X"8FC30024";
        ram_buffer(52832) := X"8FC20020";
        ram_buffer(52833) := X"8FC70014";
        ram_buffer(52834) := X"8FC60010";
        ram_buffer(52835) := X"00602821";
        ram_buffer(52836) := X"00402021";
        ram_buffer(52837) := X"0C03174A";
        ram_buffer(52838) := X"00000000";
        ram_buffer(52839) := X"03C0E821";
        ram_buffer(52840) := X"8FBF002C";
        ram_buffer(52841) := X"8FBE0028";
        ram_buffer(52842) := X"27BD0030";
        ram_buffer(52843) := X"03E00008";
        ram_buffer(52844) := X"00000000";
        ram_buffer(52845) := X"27BDFFF8";
        ram_buffer(52846) := X"AFBE0004";
        ram_buffer(52847) := X"03A0F021";
        ram_buffer(52848) := X"AFC40008";
        ram_buffer(52849) := X"AFC5000C";
        ram_buffer(52850) := X"AFC60010";
        ram_buffer(52851) := X"AFC70014";
        ram_buffer(52852) := X"8FC20014";
        ram_buffer(52853) := X"00000000";
        ram_buffer(52854) := X"30420007";
        ram_buffer(52855) := X"2C430007";
        ram_buffer(52856) := X"1060004E";
        ram_buffer(52857) := X"00000000";
        ram_buffer(52858) := X"00021880";
        ram_buffer(52859) := X"3C02100D";
        ram_buffer(52860) := X"2442AA88";
        ram_buffer(52861) := X"00621021";
        ram_buffer(52862) := X"8C420000";
        ram_buffer(52863) := X"00000000";
        ram_buffer(52864) := X"00400008";
        ram_buffer(52865) := X"00000000";
        ram_buffer(52866) := X"8FC20008";
        ram_buffer(52867) := X"00000000";
        ram_buffer(52868) := X"24420004";
        ram_buffer(52869) := X"AC400000";
        ram_buffer(52870) := X"8C430000";
        ram_buffer(52871) := X"8FC20008";
        ram_buffer(52872) := X"00000000";
        ram_buffer(52873) := X"AC430000";
        ram_buffer(52874) := X"1000003C";
        ram_buffer(52875) := X"00000000";
        ram_buffer(52876) := X"8FC20008";
        ram_buffer(52877) := X"00000000";
        ram_buffer(52878) := X"24420004";
        ram_buffer(52879) := X"8FC3000C";
        ram_buffer(52880) := X"00000000";
        ram_buffer(52881) := X"8C630000";
        ram_buffer(52882) := X"00000000";
        ram_buffer(52883) := X"AC430000";
        ram_buffer(52884) := X"8FC2000C";
        ram_buffer(52885) := X"00000000";
        ram_buffer(52886) := X"8C430004";
        ram_buffer(52887) := X"8FC20008";
        ram_buffer(52888) := X"00000000";
        ram_buffer(52889) := X"AC430000";
        ram_buffer(52890) := X"1000002C";
        ram_buffer(52891) := X"00000000";
        ram_buffer(52892) := X"8FC20008";
        ram_buffer(52893) := X"00000000";
        ram_buffer(52894) := X"24420004";
        ram_buffer(52895) := X"8FC3000C";
        ram_buffer(52896) := X"00000000";
        ram_buffer(52897) := X"8C630000";
        ram_buffer(52898) := X"00000000";
        ram_buffer(52899) := X"AC430000";
        ram_buffer(52900) := X"8FC2000C";
        ram_buffer(52901) := X"00000000";
        ram_buffer(52902) := X"24420004";
        ram_buffer(52903) := X"8C430000";
        ram_buffer(52904) := X"3C02FFEF";
        ram_buffer(52905) := X"3442FFFF";
        ram_buffer(52906) := X"00621024";
        ram_buffer(52907) := X"8FC30010";
        ram_buffer(52908) := X"00000000";
        ram_buffer(52909) := X"24630433";
        ram_buffer(52910) := X"00031D00";
        ram_buffer(52911) := X"00431825";
        ram_buffer(52912) := X"8FC20008";
        ram_buffer(52913) := X"00000000";
        ram_buffer(52914) := X"AC430000";
        ram_buffer(52915) := X"10000013";
        ram_buffer(52916) := X"00000000";
        ram_buffer(52917) := X"8FC20008";
        ram_buffer(52918) := X"3C037FF0";
        ram_buffer(52919) := X"AC430000";
        ram_buffer(52920) := X"8FC20008";
        ram_buffer(52921) := X"00000000";
        ram_buffer(52922) := X"24420004";
        ram_buffer(52923) := X"AC400000";
        ram_buffer(52924) := X"1000000A";
        ram_buffer(52925) := X"00000000";
        ram_buffer(52926) := X"8FC20008";
        ram_buffer(52927) := X"3C037FFF";
        ram_buffer(52928) := X"3463FFFF";
        ram_buffer(52929) := X"AC430000";
        ram_buffer(52930) := X"8FC20008";
        ram_buffer(52931) := X"00000000";
        ram_buffer(52932) := X"24420004";
        ram_buffer(52933) := X"2403FFFF";
        ram_buffer(52934) := X"AC430000";
        ram_buffer(52935) := X"8FC20014";
        ram_buffer(52936) := X"00000000";
        ram_buffer(52937) := X"30420008";
        ram_buffer(52938) := X"10400009";
        ram_buffer(52939) := X"00000000";
        ram_buffer(52940) := X"8FC20008";
        ram_buffer(52941) := X"00000000";
        ram_buffer(52942) := X"8C430000";
        ram_buffer(52943) := X"3C028000";
        ram_buffer(52944) := X"00621825";
        ram_buffer(52945) := X"8FC20008";
        ram_buffer(52946) := X"00000000";
        ram_buffer(52947) := X"AC430000";
        ram_buffer(52948) := X"00000000";
        ram_buffer(52949) := X"03C0E821";
        ram_buffer(52950) := X"8FBE0004";
        ram_buffer(52951) := X"27BD0008";
        ram_buffer(52952) := X"03E00008";
        ram_buffer(52953) := X"00000000";
        ram_buffer(52954) := X"27BDFFE8";
        ram_buffer(52955) := X"AFBE0014";
        ram_buffer(52956) := X"03A0F021";
        ram_buffer(52957) := X"AFC40018";
        ram_buffer(52958) := X"AFC5001C";
        ram_buffer(52959) := X"8FC20018";
        ram_buffer(52960) := X"00000000";
        ram_buffer(52961) := X"8C420000";
        ram_buffer(52962) := X"00000000";
        ram_buffer(52963) := X"AFC20004";
        ram_buffer(52964) := X"10000020";
        ram_buffer(52965) := X"00000000";
        ram_buffer(52966) := X"8FC20004";
        ram_buffer(52967) := X"00000000";
        ram_buffer(52968) := X"24420001";
        ram_buffer(52969) := X"AFC20004";
        ram_buffer(52970) := X"8FC20004";
        ram_buffer(52971) := X"00000000";
        ram_buffer(52972) := X"80420000";
        ram_buffer(52973) := X"00000000";
        ram_buffer(52974) := X"AFC20000";
        ram_buffer(52975) := X"8FC20000";
        ram_buffer(52976) := X"00000000";
        ram_buffer(52977) := X"28420041";
        ram_buffer(52978) := X"1440000A";
        ram_buffer(52979) := X"00000000";
        ram_buffer(52980) := X"8FC20000";
        ram_buffer(52981) := X"00000000";
        ram_buffer(52982) := X"2842005B";
        ram_buffer(52983) := X"10400005";
        ram_buffer(52984) := X"00000000";
        ram_buffer(52985) := X"8FC20000";
        ram_buffer(52986) := X"00000000";
        ram_buffer(52987) := X"24420020";
        ram_buffer(52988) := X"AFC20000";
        ram_buffer(52989) := X"8FC30000";
        ram_buffer(52990) := X"8FC20008";
        ram_buffer(52991) := X"00000000";
        ram_buffer(52992) := X"10620004";
        ram_buffer(52993) := X"00000000";
        ram_buffer(52994) := X"00001021";
        ram_buffer(52995) := X"10000013";
        ram_buffer(52996) := X"00000000";
        ram_buffer(52997) := X"8FC2001C";
        ram_buffer(52998) := X"00000000";
        ram_buffer(52999) := X"24430001";
        ram_buffer(53000) := X"AFC3001C";
        ram_buffer(53001) := X"80420000";
        ram_buffer(53002) := X"00000000";
        ram_buffer(53003) := X"AFC20008";
        ram_buffer(53004) := X"8FC20008";
        ram_buffer(53005) := X"00000000";
        ram_buffer(53006) := X"1440FFD7";
        ram_buffer(53007) := X"00000000";
        ram_buffer(53008) := X"8FC20004";
        ram_buffer(53009) := X"00000000";
        ram_buffer(53010) := X"24430001";
        ram_buffer(53011) := X"8FC20018";
        ram_buffer(53012) := X"00000000";
        ram_buffer(53013) := X"AC430000";
        ram_buffer(53014) := X"24020001";
        ram_buffer(53015) := X"03C0E821";
        ram_buffer(53016) := X"8FBE0014";
        ram_buffer(53017) := X"27BD0018";
        ram_buffer(53018) := X"03E00008";
        ram_buffer(53019) := X"00000000";
        ram_buffer(53020) := X"27BDFED8";
        ram_buffer(53021) := X"AFBF0124";
        ram_buffer(53022) := X"AFBE0120";
        ram_buffer(53023) := X"AFB7011C";
        ram_buffer(53024) := X"AFB60118";
        ram_buffer(53025) := X"AFB50114";
        ram_buffer(53026) := X"AFB40110";
        ram_buffer(53027) := X"AFB3010C";
        ram_buffer(53028) := X"AFB20108";
        ram_buffer(53029) := X"AFB10104";
        ram_buffer(53030) := X"AFB00100";
        ram_buffer(53031) := X"03A0F021";
        ram_buffer(53032) := X"AFC40128";
        ram_buffer(53033) := X"AFC5012C";
        ram_buffer(53034) := X"AFC60130";
        ram_buffer(53035) := X"AFC000D8";
        ram_buffer(53036) := X"AFC0007C";
        ram_buffer(53037) := X"AFC00084";
        ram_buffer(53038) := X"AFC00088";
        ram_buffer(53039) := X"AFC0007C";
        ram_buffer(53040) := X"8FC2007C";
        ram_buffer(53041) := X"00000000";
        ram_buffer(53042) := X"AFC20084";
        ram_buffer(53043) := X"8FC20084";
        ram_buffer(53044) := X"00000000";
        ram_buffer(53045) := X"AFC20088";
        ram_buffer(53046) := X"AFC00034";
        ram_buffer(53047) := X"8FC20034";
        ram_buffer(53048) := X"00000000";
        ram_buffer(53049) := X"AFC20058";
        ram_buffer(53050) := X"8FC20058";
        ram_buffer(53051) := X"00000000";
        ram_buffer(53052) := X"AFC2005C";
        ram_buffer(53053) := X"8FC2005C";
        ram_buffer(53054) := X"00000000";
        ram_buffer(53055) := X"AFC20060";
        ram_buffer(53056) := X"AFC000CC";
        ram_buffer(53057) := X"AFC000C8";
        ram_buffer(53058) := X"8FC2012C";
        ram_buffer(53059) := X"00000000";
        ram_buffer(53060) := X"AFC200B8";
        ram_buffer(53061) := X"8FC200B8";
        ram_buffer(53062) := X"00000000";
        ram_buffer(53063) := X"80420000";
        ram_buffer(53064) := X"00000000";
        ram_buffer(53065) := X"2C43002E";
        ram_buffer(53066) := X"1060001D";
        ram_buffer(53067) := X"00000000";
        ram_buffer(53068) := X"00021880";
        ram_buffer(53069) := X"3C02100D";
        ram_buffer(53070) := X"2442AAB4";
        ram_buffer(53071) := X"00621021";
        ram_buffer(53072) := X"8C420000";
        ram_buffer(53073) := X"00000000";
        ram_buffer(53074) := X"00400008";
        ram_buffer(53075) := X"00000000";
        ram_buffer(53076) := X"24020001";
        ram_buffer(53077) := X"AFC20060";
        ram_buffer(53078) := X"8FC200B8";
        ram_buffer(53079) := X"00000000";
        ram_buffer(53080) := X"24420001";
        ram_buffer(53081) := X"AFC200B8";
        ram_buffer(53082) := X"8FC200B8";
        ram_buffer(53083) := X"00000000";
        ram_buffer(53084) := X"80420000";
        ram_buffer(53085) := X"00000000";
        ram_buffer(53086) := X"10400286";
        ram_buffer(53087) := X"00000000";
        ram_buffer(53088) := X"10000008";
        ram_buffer(53089) := X"00000000";
        ram_buffer(53090) := X"8FC200B8";
        ram_buffer(53091) := X"00000000";
        ram_buffer(53092) := X"24420001";
        ram_buffer(53093) := X"AFC200B8";
        ram_buffer(53094) := X"1000FFDE";
        ram_buffer(53095) := X"00000000";
        ram_buffer(53096) := X"00000000";
        ram_buffer(53097) := X"8FC200B8";
        ram_buffer(53098) := X"00000000";
        ram_buffer(53099) := X"80430000";
        ram_buffer(53100) := X"24020030";
        ram_buffer(53101) := X"1462005E";
        ram_buffer(53102) := X"00000000";
        ram_buffer(53103) := X"8FC200B8";
        ram_buffer(53104) := X"00000000";
        ram_buffer(53105) := X"24420001";
        ram_buffer(53106) := X"80420000";
        ram_buffer(53107) := X"24030058";
        ram_buffer(53108) := X"10430004";
        ram_buffer(53109) := X"00000000";
        ram_buffer(53110) := X"24030078";
        ram_buffer(53111) := X"14430041";
        ram_buffer(53112) := X"00000000";
        ram_buffer(53113) := X"8FC200B8";
        ram_buffer(53114) := X"00000000";
        ram_buffer(53115) := X"24420001";
        ram_buffer(53116) := X"AFC2012C";
        ram_buffer(53117) := X"27C400DC";
        ram_buffer(53118) := X"27C300B8";
        ram_buffer(53119) := X"8FC20060";
        ram_buffer(53120) := X"00000000";
        ram_buffer(53121) := X"AFA20014";
        ram_buffer(53122) := X"27C200D8";
        ram_buffer(53123) := X"AFA20010";
        ram_buffer(53124) := X"00803821";
        ram_buffer(53125) := X"3C02100D";
        ram_buffer(53126) := X"2446AB6C";
        ram_buffer(53127) := X"00602821";
        ram_buffer(53128) := X"8FC40128";
        ram_buffer(53129) := X"0C02F4DF";
        ram_buffer(53130) := X"00000000";
        ram_buffer(53131) := X"AFC20044";
        ram_buffer(53132) := X"8FC20044";
        ram_buffer(53133) := X"00000000";
        ram_buffer(53134) := X"30420007";
        ram_buffer(53135) := X"1040086C";
        ram_buffer(53136) := X"00000000";
        ram_buffer(53137) := X"24030006";
        ram_buffer(53138) := X"14430008";
        ram_buffer(53139) := X"00000000";
        ram_buffer(53140) := X"8FC2012C";
        ram_buffer(53141) := X"00000000";
        ram_buffer(53142) := X"AFC200B8";
        ram_buffer(53143) := X"AFC00060";
        ram_buffer(53144) := X"00000000";
        ram_buffer(53145) := X"10000862";
        ram_buffer(53146) := X"00000000";
        ram_buffer(53147) := X"8FC200D8";
        ram_buffer(53148) := X"00000000";
        ram_buffer(53149) := X"10400010";
        ram_buffer(53150) := X"00000000";
        ram_buffer(53151) := X"3C02100D";
        ram_buffer(53152) := X"8C43AB6C";
        ram_buffer(53153) := X"8FC400D8";
        ram_buffer(53154) := X"27C200E0";
        ram_buffer(53155) := X"00803021";
        ram_buffer(53156) := X"00602821";
        ram_buffer(53157) := X"00402021";
        ram_buffer(53158) := X"0C02C5D4";
        ram_buffer(53159) := X"00000000";
        ram_buffer(53160) := X"8FC200D8";
        ram_buffer(53161) := X"00000000";
        ram_buffer(53162) := X"00402821";
        ram_buffer(53163) := X"8FC40128";
        ram_buffer(53164) := X"0C02BE10";
        ram_buffer(53165) := X"00000000";
        ram_buffer(53166) := X"8FC400DC";
        ram_buffer(53167) := X"27C300E0";
        ram_buffer(53168) := X"27C200C8";
        ram_buffer(53169) := X"8FC70044";
        ram_buffer(53170) := X"00803021";
        ram_buffer(53171) := X"00602821";
        ram_buffer(53172) := X"00402021";
        ram_buffer(53173) := X"0C02CE6D";
        ram_buffer(53174) := X"00000000";
        ram_buffer(53175) := X"10000854";
        ram_buffer(53176) := X"00000000";
        ram_buffer(53177) := X"24020001";
        ram_buffer(53178) := X"AFC2005C";
        ram_buffer(53179) := X"00000000";
        ram_buffer(53180) := X"8FC200B8";
        ram_buffer(53181) := X"00000000";
        ram_buffer(53182) := X"24420001";
        ram_buffer(53183) := X"AFC200B8";
        ram_buffer(53184) := X"8FC200B8";
        ram_buffer(53185) := X"00000000";
        ram_buffer(53186) := X"80430000";
        ram_buffer(53187) := X"24020030";
        ram_buffer(53188) := X"1062FFF7";
        ram_buffer(53189) := X"00000000";
        ram_buffer(53190) := X"8FC200B8";
        ram_buffer(53191) := X"00000000";
        ram_buffer(53192) := X"80420000";
        ram_buffer(53193) := X"00000000";
        ram_buffer(53194) := X"10400834";
        ram_buffer(53195) := X"00000000";
        ram_buffer(53196) := X"8FC200B8";
        ram_buffer(53197) := X"00000000";
        ram_buffer(53198) := X"AFC20064";
        ram_buffer(53199) := X"AFC00078";
        ram_buffer(53200) := X"8FC20078";
        ram_buffer(53201) := X"00000000";
        ram_buffer(53202) := X"AFC20074";
        ram_buffer(53203) := X"AFC00054";
        ram_buffer(53204) := X"8FC20054";
        ram_buffer(53205) := X"00000000";
        ram_buffer(53206) := X"AFC2004C";
        ram_buffer(53207) := X"10000024";
        ram_buffer(53208) := X"00000000";
        ram_buffer(53209) := X"8FC2004C";
        ram_buffer(53210) := X"00000000";
        ram_buffer(53211) := X"28420009";
        ram_buffer(53212) := X"1040000D";
        ram_buffer(53213) := X"00000000";
        ram_buffer(53214) := X"8FC20074";
        ram_buffer(53215) := X"00000000";
        ram_buffer(53216) := X"00021040";
        ram_buffer(53217) := X"00021880";
        ram_buffer(53218) := X"00431821";
        ram_buffer(53219) := X"8FC20030";
        ram_buffer(53220) := X"00000000";
        ram_buffer(53221) := X"00621021";
        ram_buffer(53222) := X"2442FFD0";
        ram_buffer(53223) := X"AFC20074";
        ram_buffer(53224) := X"1000000B";
        ram_buffer(53225) := X"00000000";
        ram_buffer(53226) := X"8FC20078";
        ram_buffer(53227) := X"00000000";
        ram_buffer(53228) := X"00021040";
        ram_buffer(53229) := X"00021880";
        ram_buffer(53230) := X"00431821";
        ram_buffer(53231) := X"8FC20030";
        ram_buffer(53232) := X"00000000";
        ram_buffer(53233) := X"00621021";
        ram_buffer(53234) := X"2442FFD0";
        ram_buffer(53235) := X"AFC20078";
        ram_buffer(53236) := X"8FC2004C";
        ram_buffer(53237) := X"00000000";
        ram_buffer(53238) := X"24420001";
        ram_buffer(53239) := X"AFC2004C";
        ram_buffer(53240) := X"8FC200B8";
        ram_buffer(53241) := X"00000000";
        ram_buffer(53242) := X"24420001";
        ram_buffer(53243) := X"AFC200B8";
        ram_buffer(53244) := X"8FC200B8";
        ram_buffer(53245) := X"00000000";
        ram_buffer(53246) := X"80420000";
        ram_buffer(53247) := X"00000000";
        ram_buffer(53248) := X"AFC20030";
        ram_buffer(53249) := X"8FC20030";
        ram_buffer(53250) := X"00000000";
        ram_buffer(53251) := X"28420030";
        ram_buffer(53252) := X"14400006";
        ram_buffer(53253) := X"00000000";
        ram_buffer(53254) := X"8FC20030";
        ram_buffer(53255) := X"00000000";
        ram_buffer(53256) := X"2842003A";
        ram_buffer(53257) := X"1440FFCF";
        ram_buffer(53258) := X"00000000";
        ram_buffer(53259) := X"8FC2004C";
        ram_buffer(53260) := X"00000000";
        ram_buffer(53261) := X"AFC20050";
        ram_buffer(53262) := X"8FC200B8";
        ram_buffer(53263) := X"00000000";
        ram_buffer(53264) := X"AFC200F0";
        ram_buffer(53265) := X"8FC40128";
        ram_buffer(53266) := X"0C02BB25";
        ram_buffer(53267) := X"00000000";
        ram_buffer(53268) := X"8C430000";
        ram_buffer(53269) := X"00000000";
        ram_buffer(53270) := X"AFC300F8";
        ram_buffer(53271) := X"8FC40128";
        ram_buffer(53272) := X"0C02BB25";
        ram_buffer(53273) := X"00000000";
        ram_buffer(53274) := X"8C420000";
        ram_buffer(53275) := X"00000000";
        ram_buffer(53276) := X"00402021";
        ram_buffer(53277) := X"0C02851E";
        ram_buffer(53278) := X"00000000";
        ram_buffer(53279) := X"00403021";
        ram_buffer(53280) := X"8FC500F8";
        ram_buffer(53281) := X"8FC400F0";
        ram_buffer(53282) := X"0C028525";
        ram_buffer(53283) := X"00000000";
        ram_buffer(53284) := X"144000B0";
        ram_buffer(53285) := X"00000000";
        ram_buffer(53286) := X"24020001";
        ram_buffer(53287) := X"AFC20034";
        ram_buffer(53288) := X"8FC40128";
        ram_buffer(53289) := X"0C02BB25";
        ram_buffer(53290) := X"00000000";
        ram_buffer(53291) := X"8C420000";
        ram_buffer(53292) := X"00000000";
        ram_buffer(53293) := X"00402021";
        ram_buffer(53294) := X"0C02851E";
        ram_buffer(53295) := X"00000000";
        ram_buffer(53296) := X"00401821";
        ram_buffer(53297) := X"8FC200B8";
        ram_buffer(53298) := X"00000000";
        ram_buffer(53299) := X"00431021";
        ram_buffer(53300) := X"AFC200B8";
        ram_buffer(53301) := X"8FC200B8";
        ram_buffer(53302) := X"00000000";
        ram_buffer(53303) := X"80420000";
        ram_buffer(53304) := X"00000000";
        ram_buffer(53305) := X"AFC20030";
        ram_buffer(53306) := X"8FC2004C";
        ram_buffer(53307) := X"00000000";
        ram_buffer(53308) := X"1440008B";
        ram_buffer(53309) := X"00000000";
        ram_buffer(53310) := X"1000000E";
        ram_buffer(53311) := X"00000000";
        ram_buffer(53312) := X"8FC20058";
        ram_buffer(53313) := X"00000000";
        ram_buffer(53314) := X"24420001";
        ram_buffer(53315) := X"AFC20058";
        ram_buffer(53316) := X"8FC200B8";
        ram_buffer(53317) := X"00000000";
        ram_buffer(53318) := X"24420001";
        ram_buffer(53319) := X"AFC200B8";
        ram_buffer(53320) := X"8FC200B8";
        ram_buffer(53321) := X"00000000";
        ram_buffer(53322) := X"80420000";
        ram_buffer(53323) := X"00000000";
        ram_buffer(53324) := X"AFC20030";
        ram_buffer(53325) := X"8FC30030";
        ram_buffer(53326) := X"24020030";
        ram_buffer(53327) := X"1062FFF0";
        ram_buffer(53328) := X"00000000";
        ram_buffer(53329) := X"8FC20030";
        ram_buffer(53330) := X"00000000";
        ram_buffer(53331) := X"28420031";
        ram_buffer(53332) := X"1440007F";
        ram_buffer(53333) := X"00000000";
        ram_buffer(53334) := X"8FC20030";
        ram_buffer(53335) := X"00000000";
        ram_buffer(53336) := X"2842003A";
        ram_buffer(53337) := X"1040007A";
        ram_buffer(53338) := X"00000000";
        ram_buffer(53339) := X"8FC200B8";
        ram_buffer(53340) := X"00000000";
        ram_buffer(53341) := X"AFC20064";
        ram_buffer(53342) := X"8FC30054";
        ram_buffer(53343) := X"8FC20058";
        ram_buffer(53344) := X"00000000";
        ram_buffer(53345) := X"00621021";
        ram_buffer(53346) := X"AFC20054";
        ram_buffer(53347) := X"AFC00058";
        ram_buffer(53348) := X"00000000";
        ram_buffer(53349) := X"8FC20058";
        ram_buffer(53350) := X"00000000";
        ram_buffer(53351) := X"24420001";
        ram_buffer(53352) := X"AFC20058";
        ram_buffer(53353) := X"8FC20030";
        ram_buffer(53354) := X"00000000";
        ram_buffer(53355) := X"2442FFD0";
        ram_buffer(53356) := X"AFC20030";
        ram_buffer(53357) := X"8FC20030";
        ram_buffer(53358) := X"00000000";
        ram_buffer(53359) := X"1040004F";
        ram_buffer(53360) := X"00000000";
        ram_buffer(53361) := X"8FC30054";
        ram_buffer(53362) := X"8FC20058";
        ram_buffer(53363) := X"00000000";
        ram_buffer(53364) := X"00621021";
        ram_buffer(53365) := X"AFC20054";
        ram_buffer(53366) := X"24020001";
        ram_buffer(53367) := X"AFC20044";
        ram_buffer(53368) := X"1000001F";
        ram_buffer(53369) := X"00000000";
        ram_buffer(53370) := X"8FC2004C";
        ram_buffer(53371) := X"00000000";
        ram_buffer(53372) := X"24430001";
        ram_buffer(53373) := X"AFC3004C";
        ram_buffer(53374) := X"28420009";
        ram_buffer(53375) := X"10400009";
        ram_buffer(53376) := X"00000000";
        ram_buffer(53377) := X"8FC20074";
        ram_buffer(53378) := X"00000000";
        ram_buffer(53379) := X"00021040";
        ram_buffer(53380) := X"00021880";
        ram_buffer(53381) := X"00431021";
        ram_buffer(53382) := X"AFC20074";
        ram_buffer(53383) := X"1000000C";
        ram_buffer(53384) := X"00000000";
        ram_buffer(53385) := X"8FC2004C";
        ram_buffer(53386) := X"00000000";
        ram_buffer(53387) := X"28420011";
        ram_buffer(53388) := X"10400007";
        ram_buffer(53389) := X"00000000";
        ram_buffer(53390) := X"8FC20078";
        ram_buffer(53391) := X"00000000";
        ram_buffer(53392) := X"00021040";
        ram_buffer(53393) := X"00021880";
        ram_buffer(53394) := X"00431021";
        ram_buffer(53395) := X"AFC20078";
        ram_buffer(53396) := X"8FC20044";
        ram_buffer(53397) := X"00000000";
        ram_buffer(53398) := X"24420001";
        ram_buffer(53399) := X"AFC20044";
        ram_buffer(53400) := X"8FC30044";
        ram_buffer(53401) := X"8FC20058";
        ram_buffer(53402) := X"00000000";
        ram_buffer(53403) := X"0062102A";
        ram_buffer(53404) := X"1440FFDD";
        ram_buffer(53405) := X"00000000";
        ram_buffer(53406) := X"8FC2004C";
        ram_buffer(53407) := X"00000000";
        ram_buffer(53408) := X"24430001";
        ram_buffer(53409) := X"AFC3004C";
        ram_buffer(53410) := X"28420009";
        ram_buffer(53411) := X"1040000C";
        ram_buffer(53412) := X"00000000";
        ram_buffer(53413) := X"8FC20074";
        ram_buffer(53414) := X"00000000";
        ram_buffer(53415) := X"00021040";
        ram_buffer(53416) := X"00021880";
        ram_buffer(53417) := X"00431821";
        ram_buffer(53418) := X"8FC20030";
        ram_buffer(53419) := X"00000000";
        ram_buffer(53420) := X"00621021";
        ram_buffer(53421) := X"AFC20074";
        ram_buffer(53422) := X"1000000F";
        ram_buffer(53423) := X"00000000";
        ram_buffer(53424) := X"8FC2004C";
        ram_buffer(53425) := X"00000000";
        ram_buffer(53426) := X"28420011";
        ram_buffer(53427) := X"1040000A";
        ram_buffer(53428) := X"00000000";
        ram_buffer(53429) := X"8FC20078";
        ram_buffer(53430) := X"00000000";
        ram_buffer(53431) := X"00021040";
        ram_buffer(53432) := X"00021880";
        ram_buffer(53433) := X"00431821";
        ram_buffer(53434) := X"8FC20030";
        ram_buffer(53435) := X"00000000";
        ram_buffer(53436) := X"00621021";
        ram_buffer(53437) := X"AFC20078";
        ram_buffer(53438) := X"AFC00058";
        ram_buffer(53439) := X"8FC200B8";
        ram_buffer(53440) := X"00000000";
        ram_buffer(53441) := X"24420001";
        ram_buffer(53442) := X"AFC200B8";
        ram_buffer(53443) := X"8FC200B8";
        ram_buffer(53444) := X"00000000";
        ram_buffer(53445) := X"80420000";
        ram_buffer(53446) := X"00000000";
        ram_buffer(53447) := X"AFC20030";
        ram_buffer(53448) := X"8FC20030";
        ram_buffer(53449) := X"00000000";
        ram_buffer(53450) := X"28420030";
        ram_buffer(53451) := X"14400009";
        ram_buffer(53452) := X"00000000";
        ram_buffer(53453) := X"8FC20030";
        ram_buffer(53454) := X"00000000";
        ram_buffer(53455) := X"2842003A";
        ram_buffer(53456) := X"1440FF94";
        ram_buffer(53457) := X"00000000";
        ram_buffer(53458) := X"10000002";
        ram_buffer(53459) := X"00000000";
        ram_buffer(53460) := X"00000000";
        ram_buffer(53461) := X"AFC00038";
        ram_buffer(53462) := X"8FC30030";
        ram_buffer(53463) := X"24020065";
        ram_buffer(53464) := X"10620005";
        ram_buffer(53465) := X"00000000";
        ram_buffer(53466) := X"8FC30030";
        ram_buffer(53467) := X"24020045";
        ram_buffer(53468) := X"1462009C";
        ram_buffer(53469) := X"00000000";
        ram_buffer(53470) := X"8FC2004C";
        ram_buffer(53471) := X"00000000";
        ram_buffer(53472) := X"14400009";
        ram_buffer(53473) := X"00000000";
        ram_buffer(53474) := X"8FC20058";
        ram_buffer(53475) := X"00000000";
        ram_buffer(53476) := X"14400005";
        ram_buffer(53477) := X"00000000";
        ram_buffer(53478) := X"8FC2005C";
        ram_buffer(53479) := X"00000000";
        ram_buffer(53480) := X"104000FF";
        ram_buffer(53481) := X"00000000";
        ram_buffer(53482) := X"8FC200B8";
        ram_buffer(53483) := X"00000000";
        ram_buffer(53484) := X"AFC2012C";
        ram_buffer(53485) := X"AFC00040";
        ram_buffer(53486) := X"8FC200B8";
        ram_buffer(53487) := X"00000000";
        ram_buffer(53488) := X"24420001";
        ram_buffer(53489) := X"AFC200B8";
        ram_buffer(53490) := X"8FC200B8";
        ram_buffer(53491) := X"00000000";
        ram_buffer(53492) := X"80420000";
        ram_buffer(53493) := X"00000000";
        ram_buffer(53494) := X"AFC20030";
        ram_buffer(53495) := X"8FC20030";
        ram_buffer(53496) := X"2403002B";
        ram_buffer(53497) := X"10430006";
        ram_buffer(53498) := X"00000000";
        ram_buffer(53499) := X"2403002D";
        ram_buffer(53500) := X"1443000C";
        ram_buffer(53501) := X"00000000";
        ram_buffer(53502) := X"24020001";
        ram_buffer(53503) := X"AFC20040";
        ram_buffer(53504) := X"8FC200B8";
        ram_buffer(53505) := X"00000000";
        ram_buffer(53506) := X"24420001";
        ram_buffer(53507) := X"AFC200B8";
        ram_buffer(53508) := X"8FC200B8";
        ram_buffer(53509) := X"00000000";
        ram_buffer(53510) := X"80420000";
        ram_buffer(53511) := X"00000000";
        ram_buffer(53512) := X"AFC20030";
        ram_buffer(53513) := X"8FC20030";
        ram_buffer(53514) := X"00000000";
        ram_buffer(53515) := X"28420030";
        ram_buffer(53516) := X"14400069";
        ram_buffer(53517) := X"00000000";
        ram_buffer(53518) := X"8FC20030";
        ram_buffer(53519) := X"00000000";
        ram_buffer(53520) := X"2842003A";
        ram_buffer(53521) := X"10400064";
        ram_buffer(53522) := X"00000000";
        ram_buffer(53523) := X"1000000A";
        ram_buffer(53524) := X"00000000";
        ram_buffer(53525) := X"8FC200B8";
        ram_buffer(53526) := X"00000000";
        ram_buffer(53527) := X"24420001";
        ram_buffer(53528) := X"AFC200B8";
        ram_buffer(53529) := X"8FC200B8";
        ram_buffer(53530) := X"00000000";
        ram_buffer(53531) := X"80420000";
        ram_buffer(53532) := X"00000000";
        ram_buffer(53533) := X"AFC20030";
        ram_buffer(53534) := X"8FC30030";
        ram_buffer(53535) := X"24020030";
        ram_buffer(53536) := X"1062FFF4";
        ram_buffer(53537) := X"00000000";
        ram_buffer(53538) := X"8FC20030";
        ram_buffer(53539) := X"00000000";
        ram_buffer(53540) := X"28420031";
        ram_buffer(53541) := X"1440004B";
        ram_buffer(53542) := X"00000000";
        ram_buffer(53543) := X"8FC20030";
        ram_buffer(53544) := X"00000000";
        ram_buffer(53545) := X"2842003A";
        ram_buffer(53546) := X"10400046";
        ram_buffer(53547) := X"00000000";
        ram_buffer(53548) := X"8FC20030";
        ram_buffer(53549) := X"00000000";
        ram_buffer(53550) := X"2442FFD0";
        ram_buffer(53551) := X"AFC20070";
        ram_buffer(53552) := X"8FC200B8";
        ram_buffer(53553) := X"00000000";
        ram_buffer(53554) := X"AFC20094";
        ram_buffer(53555) := X"1000000B";
        ram_buffer(53556) := X"00000000";
        ram_buffer(53557) := X"8FC20070";
        ram_buffer(53558) := X"00000000";
        ram_buffer(53559) := X"00021040";
        ram_buffer(53560) := X"00021880";
        ram_buffer(53561) := X"00431821";
        ram_buffer(53562) := X"8FC20030";
        ram_buffer(53563) := X"00000000";
        ram_buffer(53564) := X"00621021";
        ram_buffer(53565) := X"2442FFD0";
        ram_buffer(53566) := X"AFC20070";
        ram_buffer(53567) := X"8FC200B8";
        ram_buffer(53568) := X"00000000";
        ram_buffer(53569) := X"24420001";
        ram_buffer(53570) := X"AFC200B8";
        ram_buffer(53571) := X"8FC200B8";
        ram_buffer(53572) := X"00000000";
        ram_buffer(53573) := X"80420000";
        ram_buffer(53574) := X"00000000";
        ram_buffer(53575) := X"AFC20030";
        ram_buffer(53576) := X"8FC20030";
        ram_buffer(53577) := X"00000000";
        ram_buffer(53578) := X"28420030";
        ram_buffer(53579) := X"14400006";
        ram_buffer(53580) := X"00000000";
        ram_buffer(53581) := X"8FC20030";
        ram_buffer(53582) := X"00000000";
        ram_buffer(53583) := X"2842003A";
        ram_buffer(53584) := X"1440FFE4";
        ram_buffer(53585) := X"00000000";
        ram_buffer(53586) := X"8FC200B8";
        ram_buffer(53587) := X"00000000";
        ram_buffer(53588) := X"00401821";
        ram_buffer(53589) := X"8FC20094";
        ram_buffer(53590) := X"00000000";
        ram_buffer(53591) := X"00621023";
        ram_buffer(53592) := X"28420009";
        ram_buffer(53593) := X"10400006";
        ram_buffer(53594) := X"00000000";
        ram_buffer(53595) := X"8FC20070";
        ram_buffer(53596) := X"00000000";
        ram_buffer(53597) := X"28424E20";
        ram_buffer(53598) := X"14400005";
        ram_buffer(53599) := X"00000000";
        ram_buffer(53600) := X"24024E1F";
        ram_buffer(53601) := X"AFC20038";
        ram_buffer(53602) := X"10000004";
        ram_buffer(53603) := X"00000000";
        ram_buffer(53604) := X"8FC20070";
        ram_buffer(53605) := X"00000000";
        ram_buffer(53606) := X"AFC20038";
        ram_buffer(53607) := X"8FC20040";
        ram_buffer(53608) := X"00000000";
        ram_buffer(53609) := X"1040000A";
        ram_buffer(53610) := X"00000000";
        ram_buffer(53611) := X"8FC20038";
        ram_buffer(53612) := X"00000000";
        ram_buffer(53613) := X"00021023";
        ram_buffer(53614) := X"AFC20038";
        ram_buffer(53615) := X"10000004";
        ram_buffer(53616) := X"00000000";
        ram_buffer(53617) := X"AFC00038";
        ram_buffer(53618) := X"10000006";
        ram_buffer(53619) := X"00000000";
        ram_buffer(53620) := X"10000004";
        ram_buffer(53621) := X"00000000";
        ram_buffer(53622) := X"8FC2012C";
        ram_buffer(53623) := X"00000000";
        ram_buffer(53624) := X"AFC200B8";
        ram_buffer(53625) := X"8FC2004C";
        ram_buffer(53626) := X"00000000";
        ram_buffer(53627) := X"14400076";
        ram_buffer(53628) := X"00000000";
        ram_buffer(53629) := X"8FC20058";
        ram_buffer(53630) := X"00000000";
        ram_buffer(53631) := X"14400682";
        ram_buffer(53632) := X"00000000";
        ram_buffer(53633) := X"8FC2005C";
        ram_buffer(53634) := X"00000000";
        ram_buffer(53635) := X"1440067E";
        ram_buffer(53636) := X"00000000";
        ram_buffer(53637) := X"8FC20034";
        ram_buffer(53638) := X"00000000";
        ram_buffer(53639) := X"14400064";
        ram_buffer(53640) := X"00000000";
        ram_buffer(53641) := X"8FC20030";
        ram_buffer(53642) := X"2403004E";
        ram_buffer(53643) := X"1043002E";
        ram_buffer(53644) := X"00000000";
        ram_buffer(53645) := X"2843004F";
        ram_buffer(53646) := X"10600006";
        ram_buffer(53647) := X"00000000";
        ram_buffer(53648) := X"24030049";
        ram_buffer(53649) := X"1043000B";
        ram_buffer(53650) := X"00000000";
        ram_buffer(53651) := X"10000058";
        ram_buffer(53652) := X"00000000";
        ram_buffer(53653) := X"24030069";
        ram_buffer(53654) := X"10430006";
        ram_buffer(53655) := X"00000000";
        ram_buffer(53656) := X"2403006E";
        ram_buffer(53657) := X"10430020";
        ram_buffer(53658) := X"00000000";
        ram_buffer(53659) := X"10000050";
        ram_buffer(53660) := X"00000000";
        ram_buffer(53661) := X"27C300B8";
        ram_buffer(53662) := X"3C02100D";
        ram_buffer(53663) := X"2445AAA4";
        ram_buffer(53664) := X"00602021";
        ram_buffer(53665) := X"0C02CEDA";
        ram_buffer(53666) := X"00000000";
        ram_buffer(53667) := X"10400047";
        ram_buffer(53668) := X"00000000";
        ram_buffer(53669) := X"8FC200B8";
        ram_buffer(53670) := X"00000000";
        ram_buffer(53671) := X"2442FFFF";
        ram_buffer(53672) := X"AFC200B8";
        ram_buffer(53673) := X"27C300B8";
        ram_buffer(53674) := X"3C02100D";
        ram_buffer(53675) := X"2445AAA8";
        ram_buffer(53676) := X"00602021";
        ram_buffer(53677) := X"0C02CEDA";
        ram_buffer(53678) := X"00000000";
        ram_buffer(53679) := X"14400005";
        ram_buffer(53680) := X"00000000";
        ram_buffer(53681) := X"8FC200B8";
        ram_buffer(53682) := X"00000000";
        ram_buffer(53683) := X"24420001";
        ram_buffer(53684) := X"AFC200B8";
        ram_buffer(53685) := X"3C027FF0";
        ram_buffer(53686) := X"AFC200C8";
        ram_buffer(53687) := X"AFC000CC";
        ram_buffer(53688) := X"10000653";
        ram_buffer(53689) := X"00000000";
        ram_buffer(53690) := X"27C300B8";
        ram_buffer(53691) := X"3C02100D";
        ram_buffer(53692) := X"2445AAB0";
        ram_buffer(53693) := X"00602021";
        ram_buffer(53694) := X"0C02CEDA";
        ram_buffer(53695) := X"00000000";
        ram_buffer(53696) := X"1040002B";
        ram_buffer(53697) := X"00000000";
        ram_buffer(53698) := X"8FC200B8";
        ram_buffer(53699) := X"00000000";
        ram_buffer(53700) := X"80430000";
        ram_buffer(53701) := X"24020028";
        ram_buffer(53702) := X"14620016";
        ram_buffer(53703) := X"00000000";
        ram_buffer(53704) := X"27C200E8";
        ram_buffer(53705) := X"27C300B8";
        ram_buffer(53706) := X"00403021";
        ram_buffer(53707) := X"3C02100D";
        ram_buffer(53708) := X"2445AB80";
        ram_buffer(53709) := X"00602021";
        ram_buffer(53710) := X"0C02F8D0";
        ram_buffer(53711) := X"00000000";
        ram_buffer(53712) := X"00401821";
        ram_buffer(53713) := X"24020005";
        ram_buffer(53714) := X"1462000A";
        ram_buffer(53715) := X"00000000";
        ram_buffer(53716) := X"8FC300EC";
        ram_buffer(53717) := X"3C027FF0";
        ram_buffer(53718) := X"00621025";
        ram_buffer(53719) := X"AFC200C8";
        ram_buffer(53720) := X"8FC200E8";
        ram_buffer(53721) := X"00000000";
        ram_buffer(53722) := X"AFC200CC";
        ram_buffer(53723) := X"10000630";
        ram_buffer(53724) := X"00000000";
        ram_buffer(53725) := X"3C027FF7";
        ram_buffer(53726) := X"3442FFFF";
        ram_buffer(53727) := X"AFC200C8";
        ram_buffer(53728) := X"2402FFFF";
        ram_buffer(53729) := X"AFC200CC";
        ram_buffer(53730) := X"00000000";
        ram_buffer(53731) := X"10000628";
        ram_buffer(53732) := X"00000000";
        ram_buffer(53733) := X"00000000";
        ram_buffer(53734) := X"10000005";
        ram_buffer(53735) := X"00000000";
        ram_buffer(53736) := X"00000000";
        ram_buffer(53737) := X"10000002";
        ram_buffer(53738) := X"00000000";
        ram_buffer(53739) := X"00000000";
        ram_buffer(53740) := X"8FC2012C";
        ram_buffer(53741) := X"00000000";
        ram_buffer(53742) := X"AFC200B8";
        ram_buffer(53743) := X"AFC00060";
        ram_buffer(53744) := X"10000611";
        ram_buffer(53745) := X"00000000";
        ram_buffer(53746) := X"8FC30038";
        ram_buffer(53747) := X"8FC20054";
        ram_buffer(53748) := X"00000000";
        ram_buffer(53749) := X"00621023";
        ram_buffer(53750) := X"AFC20038";
        ram_buffer(53751) := X"8FC20038";
        ram_buffer(53752) := X"00000000";
        ram_buffer(53753) := X"AFC2003C";
        ram_buffer(53754) := X"8FC20050";
        ram_buffer(53755) := X"00000000";
        ram_buffer(53756) := X"14400004";
        ram_buffer(53757) := X"00000000";
        ram_buffer(53758) := X"8FC2004C";
        ram_buffer(53759) := X"00000000";
        ram_buffer(53760) := X"AFC20050";
        ram_buffer(53761) := X"8FC2004C";
        ram_buffer(53762) := X"00000000";
        ram_buffer(53763) := X"28430011";
        ram_buffer(53764) := X"14600002";
        ram_buffer(53765) := X"00000000";
        ram_buffer(53766) := X"24020010";
        ram_buffer(53767) := X"AFC20098";
        ram_buffer(53768) := X"8FC40074";
        ram_buffer(53769) := X"0C031BBD";
        ram_buffer(53770) := X"00000000";
        ram_buffer(53771) := X"AFC300CC";
        ram_buffer(53772) := X"AFC200C8";
        ram_buffer(53773) := X"8FC20098";
        ram_buffer(53774) := X"00000000";
        ram_buffer(53775) := X"2842000A";
        ram_buffer(53776) := X"1440001F";
        ram_buffer(53777) := X"00000000";
        ram_buffer(53778) := X"8FC20098";
        ram_buffer(53779) := X"00000000";
        ram_buffer(53780) := X"2443FFF7";
        ram_buffer(53781) := X"3C02100D";
        ram_buffer(53782) := X"000318C0";
        ram_buffer(53783) := X"2442A938";
        ram_buffer(53784) := X"00621021";
        ram_buffer(53785) := X"8C430004";
        ram_buffer(53786) := X"8C420000";
        ram_buffer(53787) := X"8FC500CC";
        ram_buffer(53788) := X"8FC400C8";
        ram_buffer(53789) := X"00A03821";
        ram_buffer(53790) := X"00803021";
        ram_buffer(53791) := X"00602821";
        ram_buffer(53792) := X"00402021";
        ram_buffer(53793) := X"0C03174A";
        ram_buffer(53794) := X"00000000";
        ram_buffer(53795) := X"AFC300F4";
        ram_buffer(53796) := X"AFC200F0";
        ram_buffer(53797) := X"8FC40078";
        ram_buffer(53798) := X"0C031BBD";
        ram_buffer(53799) := X"00000000";
        ram_buffer(53800) := X"00603821";
        ram_buffer(53801) := X"00403021";
        ram_buffer(53802) := X"8FC500F4";
        ram_buffer(53803) := X"8FC400F0";
        ram_buffer(53804) := X"0C0311FC";
        ram_buffer(53805) := X"00000000";
        ram_buffer(53806) := X"AFC300CC";
        ram_buffer(53807) := X"AFC200C8";
        ram_buffer(53808) := X"AFC00080";
        ram_buffer(53809) := X"8FC2004C";
        ram_buffer(53810) := X"00000000";
        ram_buffer(53811) := X"28420010";
        ram_buffer(53812) := X"10400074";
        ram_buffer(53813) := X"00000000";
        ram_buffer(53814) := X"8FC20038";
        ram_buffer(53815) := X"00000000";
        ram_buffer(53816) := X"104005CC";
        ram_buffer(53817) := X"00000000";
        ram_buffer(53818) := X"8FC20038";
        ram_buffer(53819) := X"00000000";
        ram_buffer(53820) := X"18400052";
        ram_buffer(53821) := X"00000000";
        ram_buffer(53822) := X"8FC20038";
        ram_buffer(53823) := X"00000000";
        ram_buffer(53824) := X"28420017";
        ram_buffer(53825) := X"10400015";
        ram_buffer(53826) := X"00000000";
        ram_buffer(53827) := X"8FC300CC";
        ram_buffer(53828) := X"8FC200C8";
        ram_buffer(53829) := X"3C04100D";
        ram_buffer(53830) := X"8FC50038";
        ram_buffer(53831) := X"00000000";
        ram_buffer(53832) := X"000528C0";
        ram_buffer(53833) := X"2484A938";
        ram_buffer(53834) := X"00A42021";
        ram_buffer(53835) := X"8C850004";
        ram_buffer(53836) := X"8C840000";
        ram_buffer(53837) := X"00A03821";
        ram_buffer(53838) := X"00803021";
        ram_buffer(53839) := X"00602821";
        ram_buffer(53840) := X"00402021";
        ram_buffer(53841) := X"0C03174A";
        ram_buffer(53842) := X"00000000";
        ram_buffer(53843) := X"AFC300CC";
        ram_buffer(53844) := X"AFC200C8";
        ram_buffer(53845) := X"100005B6";
        ram_buffer(53846) := X"00000000";
        ram_buffer(53847) := X"2403000F";
        ram_buffer(53848) := X"8FC2004C";
        ram_buffer(53849) := X"00000000";
        ram_buffer(53850) := X"00621023";
        ram_buffer(53851) := X"AFC20044";
        ram_buffer(53852) := X"8FC20044";
        ram_buffer(53853) := X"00000000";
        ram_buffer(53854) := X"24430016";
        ram_buffer(53855) := X"8FC20038";
        ram_buffer(53856) := X"00000000";
        ram_buffer(53857) := X"0062102A";
        ram_buffer(53858) := X"14400046";
        ram_buffer(53859) := X"00000000";
        ram_buffer(53860) := X"8FC30038";
        ram_buffer(53861) := X"8FC20044";
        ram_buffer(53862) := X"00000000";
        ram_buffer(53863) := X"00621023";
        ram_buffer(53864) := X"AFC20038";
        ram_buffer(53865) := X"8FC300CC";
        ram_buffer(53866) := X"8FC200C8";
        ram_buffer(53867) := X"3C04100D";
        ram_buffer(53868) := X"8FC50044";
        ram_buffer(53869) := X"00000000";
        ram_buffer(53870) := X"000528C0";
        ram_buffer(53871) := X"2484A938";
        ram_buffer(53872) := X"00A42021";
        ram_buffer(53873) := X"8C850004";
        ram_buffer(53874) := X"8C840000";
        ram_buffer(53875) := X"00A03821";
        ram_buffer(53876) := X"00803021";
        ram_buffer(53877) := X"00602821";
        ram_buffer(53878) := X"00402021";
        ram_buffer(53879) := X"0C03174A";
        ram_buffer(53880) := X"00000000";
        ram_buffer(53881) := X"AFC300CC";
        ram_buffer(53882) := X"AFC200C8";
        ram_buffer(53883) := X"8FC300CC";
        ram_buffer(53884) := X"8FC200C8";
        ram_buffer(53885) := X"3C04100D";
        ram_buffer(53886) := X"8FC50038";
        ram_buffer(53887) := X"00000000";
        ram_buffer(53888) := X"000528C0";
        ram_buffer(53889) := X"2484A938";
        ram_buffer(53890) := X"00A42021";
        ram_buffer(53891) := X"8C850004";
        ram_buffer(53892) := X"8C840000";
        ram_buffer(53893) := X"00A03821";
        ram_buffer(53894) := X"00803021";
        ram_buffer(53895) := X"00602821";
        ram_buffer(53896) := X"00402021";
        ram_buffer(53897) := X"0C03174A";
        ram_buffer(53898) := X"00000000";
        ram_buffer(53899) := X"AFC300CC";
        ram_buffer(53900) := X"AFC200C8";
        ram_buffer(53901) := X"1000057E";
        ram_buffer(53902) := X"00000000";
        ram_buffer(53903) := X"8FC20038";
        ram_buffer(53904) := X"00000000";
        ram_buffer(53905) := X"2842FFEA";
        ram_buffer(53906) := X"14400016";
        ram_buffer(53907) := X"00000000";
        ram_buffer(53908) := X"8FC300CC";
        ram_buffer(53909) := X"8FC200C8";
        ram_buffer(53910) := X"8FC40038";
        ram_buffer(53911) := X"00000000";
        ram_buffer(53912) := X"00042823";
        ram_buffer(53913) := X"3C04100D";
        ram_buffer(53914) := X"000528C0";
        ram_buffer(53915) := X"2484A938";
        ram_buffer(53916) := X"00A42021";
        ram_buffer(53917) := X"8C850004";
        ram_buffer(53918) := X"8C840000";
        ram_buffer(53919) := X"00A03821";
        ram_buffer(53920) := X"00803021";
        ram_buffer(53921) := X"00602821";
        ram_buffer(53922) := X"00402021";
        ram_buffer(53923) := X"0C03144F";
        ram_buffer(53924) := X"00000000";
        ram_buffer(53925) := X"AFC300CC";
        ram_buffer(53926) := X"AFC200C8";
        ram_buffer(53927) := X"10000564";
        ram_buffer(53928) := X"00000000";
        ram_buffer(53929) := X"8FC3004C";
        ram_buffer(53930) := X"8FC20098";
        ram_buffer(53931) := X"00000000";
        ram_buffer(53932) := X"00621023";
        ram_buffer(53933) := X"8FC3003C";
        ram_buffer(53934) := X"00000000";
        ram_buffer(53935) := X"00621021";
        ram_buffer(53936) := X"AFC2003C";
        ram_buffer(53937) := X"AFC00018";
        ram_buffer(53938) := X"8FC2003C";
        ram_buffer(53939) := X"00000000";
        ram_buffer(53940) := X"184000BC";
        ram_buffer(53941) := X"00000000";
        ram_buffer(53942) := X"8FC2003C";
        ram_buffer(53943) := X"00000000";
        ram_buffer(53944) := X"3042000F";
        ram_buffer(53945) := X"AFC20044";
        ram_buffer(53946) := X"8FC20044";
        ram_buffer(53947) := X"00000000";
        ram_buffer(53948) := X"10400013";
        ram_buffer(53949) := X"00000000";
        ram_buffer(53950) := X"8FC300CC";
        ram_buffer(53951) := X"8FC200C8";
        ram_buffer(53952) := X"3C04100D";
        ram_buffer(53953) := X"8FC50044";
        ram_buffer(53954) := X"00000000";
        ram_buffer(53955) := X"000528C0";
        ram_buffer(53956) := X"2484A938";
        ram_buffer(53957) := X"00A42021";
        ram_buffer(53958) := X"8C850004";
        ram_buffer(53959) := X"8C840000";
        ram_buffer(53960) := X"00A03821";
        ram_buffer(53961) := X"00803021";
        ram_buffer(53962) := X"00602821";
        ram_buffer(53963) := X"00402021";
        ram_buffer(53964) := X"0C03174A";
        ram_buffer(53965) := X"00000000";
        ram_buffer(53966) := X"AFC300CC";
        ram_buffer(53967) := X"AFC200C8";
        ram_buffer(53968) := X"8FC3003C";
        ram_buffer(53969) := X"2402FFF0";
        ram_buffer(53970) := X"00621024";
        ram_buffer(53971) := X"AFC2003C";
        ram_buffer(53972) := X"8FC2003C";
        ram_buffer(53973) := X"00000000";
        ram_buffer(53974) := X"10400146";
        ram_buffer(53975) := X"00000000";
        ram_buffer(53976) := X"8FC2003C";
        ram_buffer(53977) := X"00000000";
        ram_buffer(53978) := X"28420135";
        ram_buffer(53979) := X"14400037";
        ram_buffer(53980) := X"00000000";
        ram_buffer(53981) := X"10000029";
        ram_buffer(53982) := X"00000000";
        ram_buffer(53983) := X"00000000";
        ram_buffer(53984) := X"10000026";
        ram_buffer(53985) := X"00000000";
        ram_buffer(53986) := X"00000000";
        ram_buffer(53987) := X"10000023";
        ram_buffer(53988) := X"00000000";
        ram_buffer(53989) := X"00000000";
        ram_buffer(53990) := X"10000020";
        ram_buffer(53991) := X"00000000";
        ram_buffer(53992) := X"00000000";
        ram_buffer(53993) := X"1000001D";
        ram_buffer(53994) := X"00000000";
        ram_buffer(53995) := X"00000000";
        ram_buffer(53996) := X"1000001A";
        ram_buffer(53997) := X"00000000";
        ram_buffer(53998) := X"00000000";
        ram_buffer(53999) := X"10000017";
        ram_buffer(54000) := X"00000000";
        ram_buffer(54001) := X"00000000";
        ram_buffer(54002) := X"10000014";
        ram_buffer(54003) := X"00000000";
        ram_buffer(54004) := X"00000000";
        ram_buffer(54005) := X"10000011";
        ram_buffer(54006) := X"00000000";
        ram_buffer(54007) := X"00000000";
        ram_buffer(54008) := X"1000000E";
        ram_buffer(54009) := X"00000000";
        ram_buffer(54010) := X"00000000";
        ram_buffer(54011) := X"1000000B";
        ram_buffer(54012) := X"00000000";
        ram_buffer(54013) := X"00000000";
        ram_buffer(54014) := X"10000008";
        ram_buffer(54015) := X"00000000";
        ram_buffer(54016) := X"00000000";
        ram_buffer(54017) := X"10000005";
        ram_buffer(54018) := X"00000000";
        ram_buffer(54019) := X"00000000";
        ram_buffer(54020) := X"10000002";
        ram_buffer(54021) := X"00000000";
        ram_buffer(54022) := X"00000000";
        ram_buffer(54023) := X"8FC20128";
        ram_buffer(54024) := X"24030022";
        ram_buffer(54025) := X"AC430000";
        ram_buffer(54026) := X"3C027FF0";
        ram_buffer(54027) := X"AFC200C8";
        ram_buffer(54028) := X"AFC000CC";
        ram_buffer(54029) := X"8FC20080";
        ram_buffer(54030) := X"00000000";
        ram_buffer(54031) := X"104004F8";
        ram_buffer(54032) := X"00000000";
        ram_buffer(54033) := X"100004D2";
        ram_buffer(54034) := X"00000000";
        ram_buffer(54035) := X"8FC2003C";
        ram_buffer(54036) := X"00000000";
        ram_buffer(54037) := X"00021103";
        ram_buffer(54038) := X"AFC2003C";
        ram_buffer(54039) := X"AFC00048";
        ram_buffer(54040) := X"10000020";
        ram_buffer(54041) := X"00000000";
        ram_buffer(54042) := X"8FC2003C";
        ram_buffer(54043) := X"00000000";
        ram_buffer(54044) := X"30420001";
        ram_buffer(54045) := X"10400013";
        ram_buffer(54046) := X"00000000";
        ram_buffer(54047) := X"8FC300CC";
        ram_buffer(54048) := X"8FC200C8";
        ram_buffer(54049) := X"3C04100D";
        ram_buffer(54050) := X"8FC50048";
        ram_buffer(54051) := X"00000000";
        ram_buffer(54052) := X"000528C0";
        ram_buffer(54053) := X"2484AA00";
        ram_buffer(54054) := X"00A42021";
        ram_buffer(54055) := X"8C850004";
        ram_buffer(54056) := X"8C840000";
        ram_buffer(54057) := X"00A03821";
        ram_buffer(54058) := X"00803021";
        ram_buffer(54059) := X"00602821";
        ram_buffer(54060) := X"00402021";
        ram_buffer(54061) := X"0C03174A";
        ram_buffer(54062) := X"00000000";
        ram_buffer(54063) := X"AFC300CC";
        ram_buffer(54064) := X"AFC200C8";
        ram_buffer(54065) := X"8FC20048";
        ram_buffer(54066) := X"00000000";
        ram_buffer(54067) := X"24420001";
        ram_buffer(54068) := X"AFC20048";
        ram_buffer(54069) := X"8FC2003C";
        ram_buffer(54070) := X"00000000";
        ram_buffer(54071) := X"00021043";
        ram_buffer(54072) := X"AFC2003C";
        ram_buffer(54073) := X"8FC2003C";
        ram_buffer(54074) := X"00000000";
        ram_buffer(54075) := X"28420002";
        ram_buffer(54076) := X"1040FFDD";
        ram_buffer(54077) := X"00000000";
        ram_buffer(54078) := X"8FC300C8";
        ram_buffer(54079) := X"3C02FCB0";
        ram_buffer(54080) := X"00621021";
        ram_buffer(54081) := X"AFC200C8";
        ram_buffer(54082) := X"8FC300CC";
        ram_buffer(54083) := X"8FC200C8";
        ram_buffer(54084) := X"3C04100D";
        ram_buffer(54085) := X"8FC50048";
        ram_buffer(54086) := X"00000000";
        ram_buffer(54087) := X"000528C0";
        ram_buffer(54088) := X"2484AA00";
        ram_buffer(54089) := X"00A42021";
        ram_buffer(54090) := X"8C850004";
        ram_buffer(54091) := X"8C840000";
        ram_buffer(54092) := X"00A03821";
        ram_buffer(54093) := X"00803021";
        ram_buffer(54094) := X"00602821";
        ram_buffer(54095) := X"00402021";
        ram_buffer(54096) := X"0C03174A";
        ram_buffer(54097) := X"00000000";
        ram_buffer(54098) := X"AFC300CC";
        ram_buffer(54099) := X"AFC200C8";
        ram_buffer(54100) := X"8FC300C8";
        ram_buffer(54101) := X"3C027FF0";
        ram_buffer(54102) := X"00621024";
        ram_buffer(54103) := X"AFC20078";
        ram_buffer(54104) := X"8FC30078";
        ram_buffer(54105) := X"3C027CA0";
        ram_buffer(54106) := X"34420001";
        ram_buffer(54107) := X"0062102B";
        ram_buffer(54108) := X"1040FF82";
        ram_buffer(54109) := X"00000000";
        ram_buffer(54110) := X"8FC30078";
        ram_buffer(54111) := X"3C027C90";
        ram_buffer(54112) := X"34420001";
        ram_buffer(54113) := X"0062102B";
        ram_buffer(54114) := X"14400008";
        ram_buffer(54115) := X"00000000";
        ram_buffer(54116) := X"3C027FEF";
        ram_buffer(54117) := X"3442FFFF";
        ram_buffer(54118) := X"AFC200C8";
        ram_buffer(54119) := X"2402FFFF";
        ram_buffer(54120) := X"AFC200CC";
        ram_buffer(54121) := X"100000B3";
        ram_buffer(54122) := X"00000000";
        ram_buffer(54123) := X"8FC300C8";
        ram_buffer(54124) := X"3C020350";
        ram_buffer(54125) := X"00621021";
        ram_buffer(54126) := X"AFC200C8";
        ram_buffer(54127) := X"100000AD";
        ram_buffer(54128) := X"00000000";
        ram_buffer(54129) := X"8FC2003C";
        ram_buffer(54130) := X"00000000";
        ram_buffer(54131) := X"044100A9";
        ram_buffer(54132) := X"00000000";
        ram_buffer(54133) := X"8FC2003C";
        ram_buffer(54134) := X"00000000";
        ram_buffer(54135) := X"00021023";
        ram_buffer(54136) := X"AFC2003C";
        ram_buffer(54137) := X"8FC2003C";
        ram_buffer(54138) := X"00000000";
        ram_buffer(54139) := X"3042000F";
        ram_buffer(54140) := X"AFC20044";
        ram_buffer(54141) := X"8FC20044";
        ram_buffer(54142) := X"00000000";
        ram_buffer(54143) := X"10400013";
        ram_buffer(54144) := X"00000000";
        ram_buffer(54145) := X"8FC300CC";
        ram_buffer(54146) := X"8FC200C8";
        ram_buffer(54147) := X"3C04100D";
        ram_buffer(54148) := X"8FC50044";
        ram_buffer(54149) := X"00000000";
        ram_buffer(54150) := X"000528C0";
        ram_buffer(54151) := X"2484A938";
        ram_buffer(54152) := X"00A42021";
        ram_buffer(54153) := X"8C850004";
        ram_buffer(54154) := X"8C840000";
        ram_buffer(54155) := X"00A03821";
        ram_buffer(54156) := X"00803021";
        ram_buffer(54157) := X"00602821";
        ram_buffer(54158) := X"00402021";
        ram_buffer(54159) := X"0C03144F";
        ram_buffer(54160) := X"00000000";
        ram_buffer(54161) := X"AFC300CC";
        ram_buffer(54162) := X"AFC200C8";
        ram_buffer(54163) := X"8FC2003C";
        ram_buffer(54164) := X"00000000";
        ram_buffer(54165) := X"00021103";
        ram_buffer(54166) := X"AFC2003C";
        ram_buffer(54167) := X"8FC2003C";
        ram_buffer(54168) := X"00000000";
        ram_buffer(54169) := X"10400083";
        ram_buffer(54170) := X"00000000";
        ram_buffer(54171) := X"8FC2003C";
        ram_buffer(54172) := X"00000000";
        ram_buffer(54173) := X"28420020";
        ram_buffer(54174) := X"10400069";
        ram_buffer(54175) := X"00000000";
        ram_buffer(54176) := X"8FC2003C";
        ram_buffer(54177) := X"00000000";
        ram_buffer(54178) := X"30420010";
        ram_buffer(54179) := X"10400003";
        ram_buffer(54180) := X"00000000";
        ram_buffer(54181) := X"2402006A";
        ram_buffer(54182) := X"AFC20018";
        ram_buffer(54183) := X"AFC00048";
        ram_buffer(54184) := X"10000020";
        ram_buffer(54185) := X"00000000";
        ram_buffer(54186) := X"8FC2003C";
        ram_buffer(54187) := X"00000000";
        ram_buffer(54188) := X"30420001";
        ram_buffer(54189) := X"10400013";
        ram_buffer(54190) := X"00000000";
        ram_buffer(54191) := X"8FC300CC";
        ram_buffer(54192) := X"8FC200C8";
        ram_buffer(54193) := X"3C04100D";
        ram_buffer(54194) := X"8FC50048";
        ram_buffer(54195) := X"00000000";
        ram_buffer(54196) := X"000528C0";
        ram_buffer(54197) := X"2484AA60";
        ram_buffer(54198) := X"00A42021";
        ram_buffer(54199) := X"8C850004";
        ram_buffer(54200) := X"8C840000";
        ram_buffer(54201) := X"00A03821";
        ram_buffer(54202) := X"00803021";
        ram_buffer(54203) := X"00602821";
        ram_buffer(54204) := X"00402021";
        ram_buffer(54205) := X"0C03174A";
        ram_buffer(54206) := X"00000000";
        ram_buffer(54207) := X"AFC300CC";
        ram_buffer(54208) := X"AFC200C8";
        ram_buffer(54209) := X"8FC20048";
        ram_buffer(54210) := X"00000000";
        ram_buffer(54211) := X"24420001";
        ram_buffer(54212) := X"AFC20048";
        ram_buffer(54213) := X"8FC2003C";
        ram_buffer(54214) := X"00000000";
        ram_buffer(54215) := X"00021043";
        ram_buffer(54216) := X"AFC2003C";
        ram_buffer(54217) := X"8FC2003C";
        ram_buffer(54218) := X"00000000";
        ram_buffer(54219) := X"1C40FFDE";
        ram_buffer(54220) := X"00000000";
        ram_buffer(54221) := X"8FC20018";
        ram_buffer(54222) := X"00000000";
        ram_buffer(54223) := X"1040002C";
        ram_buffer(54224) := X"00000000";
        ram_buffer(54225) := X"8FC300C8";
        ram_buffer(54226) := X"3C027FF0";
        ram_buffer(54227) := X"00621024";
        ram_buffer(54228) := X"00021502";
        ram_buffer(54229) := X"2403006B";
        ram_buffer(54230) := X"00621023";
        ram_buffer(54231) := X"AFC20048";
        ram_buffer(54232) := X"8FC20048";
        ram_buffer(54233) := X"00000000";
        ram_buffer(54234) := X"18400021";
        ram_buffer(54235) := X"00000000";
        ram_buffer(54236) := X"8FC20048";
        ram_buffer(54237) := X"00000000";
        ram_buffer(54238) := X"28420020";
        ram_buffer(54239) := X"14400015";
        ram_buffer(54240) := X"00000000";
        ram_buffer(54241) := X"AFC000CC";
        ram_buffer(54242) := X"8FC20048";
        ram_buffer(54243) := X"00000000";
        ram_buffer(54244) := X"28420035";
        ram_buffer(54245) := X"14400005";
        ram_buffer(54246) := X"00000000";
        ram_buffer(54247) := X"3C020370";
        ram_buffer(54248) := X"AFC200C8";
        ram_buffer(54249) := X"10000012";
        ram_buffer(54250) := X"00000000";
        ram_buffer(54251) := X"8FC300C8";
        ram_buffer(54252) := X"8FC20048";
        ram_buffer(54253) := X"00000000";
        ram_buffer(54254) := X"2442FFE0";
        ram_buffer(54255) := X"2404FFFF";
        ram_buffer(54256) := X"00441004";
        ram_buffer(54257) := X"00621024";
        ram_buffer(54258) := X"AFC200C8";
        ram_buffer(54259) := X"10000008";
        ram_buffer(54260) := X"00000000";
        ram_buffer(54261) := X"8FC300CC";
        ram_buffer(54262) := X"2404FFFF";
        ram_buffer(54263) := X"8FC20048";
        ram_buffer(54264) := X"00000000";
        ram_buffer(54265) := X"00441004";
        ram_buffer(54266) := X"00621024";
        ram_buffer(54267) := X"AFC200CC";
        ram_buffer(54268) := X"8FC300CC";
        ram_buffer(54269) := X"8FC200C8";
        ram_buffer(54270) := X"00003821";
        ram_buffer(54271) := X"00003021";
        ram_buffer(54272) := X"00602821";
        ram_buffer(54273) := X"00402021";
        ram_buffer(54274) := X"0C03167F";
        ram_buffer(54275) := X"00000000";
        ram_buffer(54276) := X"14400018";
        ram_buffer(54277) := X"00000000";
        ram_buffer(54278) := X"1000000B";
        ram_buffer(54279) := X"00000000";
        ram_buffer(54280) := X"00000000";
        ram_buffer(54281) := X"10000008";
        ram_buffer(54282) := X"00000000";
        ram_buffer(54283) := X"00000000";
        ram_buffer(54284) := X"10000005";
        ram_buffer(54285) := X"00000000";
        ram_buffer(54286) := X"00000000";
        ram_buffer(54287) := X"10000002";
        ram_buffer(54288) := X"00000000";
        ram_buffer(54289) := X"00000000";
        ram_buffer(54290) := X"AFC000CC";
        ram_buffer(54291) := X"AFC000C8";
        ram_buffer(54292) := X"8FC20128";
        ram_buffer(54293) := X"24030022";
        ram_buffer(54294) := X"AC430000";
        ram_buffer(54295) := X"8FC20080";
        ram_buffer(54296) := X"00000000";
        ram_buffer(54297) := X"104003F1";
        ram_buffer(54298) := X"00000000";
        ram_buffer(54299) := X"100003C8";
        ram_buffer(54300) := X"00000000";
        ram_buffer(54301) := X"8FC20074";
        ram_buffer(54302) := X"00000000";
        ram_buffer(54303) := X"AFA20010";
        ram_buffer(54304) := X"8FC7004C";
        ram_buffer(54305) := X"8FC60050";
        ram_buffer(54306) := X"8FC50064";
        ram_buffer(54307) := X"8FC40128";
        ram_buffer(54308) := X"0C02BEC2";
        ram_buffer(54309) := X"00000000";
        ram_buffer(54310) := X"AFC20080";
        ram_buffer(54311) := X"8FC20080";
        ram_buffer(54312) := X"00000000";
        ram_buffer(54313) := X"1040FEB8";
        ram_buffer(54314) := X"00000000";
        ram_buffer(54315) := X"8FC20080";
        ram_buffer(54316) := X"00000000";
        ram_buffer(54317) := X"8C420004";
        ram_buffer(54318) := X"00000000";
        ram_buffer(54319) := X"00402821";
        ram_buffer(54320) := X"8FC40128";
        ram_buffer(54321) := X"0C02BDA8";
        ram_buffer(54322) := X"00000000";
        ram_buffer(54323) := X"AFC2007C";
        ram_buffer(54324) := X"8FC2007C";
        ram_buffer(54325) := X"00000000";
        ram_buffer(54326) := X"1040FEAE";
        ram_buffer(54327) := X"00000000";
        ram_buffer(54328) := X"8FC2007C";
        ram_buffer(54329) := X"00000000";
        ram_buffer(54330) := X"2443000C";
        ram_buffer(54331) := X"8FC20080";
        ram_buffer(54332) := X"00000000";
        ram_buffer(54333) := X"2444000C";
        ram_buffer(54334) := X"8FC20080";
        ram_buffer(54335) := X"00000000";
        ram_buffer(54336) := X"8C420010";
        ram_buffer(54337) := X"00000000";
        ram_buffer(54338) := X"24420002";
        ram_buffer(54339) := X"00021080";
        ram_buffer(54340) := X"00403021";
        ram_buffer(54341) := X"00802821";
        ram_buffer(54342) := X"00602021";
        ram_buffer(54343) := X"0C027F93";
        ram_buffer(54344) := X"00000000";
        ram_buffer(54345) := X"8FC300CC";
        ram_buffer(54346) := X"8FC200C8";
        ram_buffer(54347) := X"27C400B4";
        ram_buffer(54348) := X"AFA40014";
        ram_buffer(54349) := X"27C400B0";
        ram_buffer(54350) := X"AFA40010";
        ram_buffer(54351) := X"00603821";
        ram_buffer(54352) := X"00403021";
        ram_buffer(54353) := X"8FC40128";
        ram_buffer(54354) := X"0C02C49D";
        ram_buffer(54355) := X"00000000";
        ram_buffer(54356) := X"AFC200D8";
        ram_buffer(54357) := X"8FC200D8";
        ram_buffer(54358) := X"00000000";
        ram_buffer(54359) := X"1040FE90";
        ram_buffer(54360) := X"00000000";
        ram_buffer(54361) := X"24050001";
        ram_buffer(54362) := X"8FC40128";
        ram_buffer(54363) := X"0C02BFBF";
        ram_buffer(54364) := X"00000000";
        ram_buffer(54365) := X"AFC20084";
        ram_buffer(54366) := X"8FC20084";
        ram_buffer(54367) := X"00000000";
        ram_buffer(54368) := X"1040FE8A";
        ram_buffer(54369) := X"00000000";
        ram_buffer(54370) := X"8FC20038";
        ram_buffer(54371) := X"00000000";
        ram_buffer(54372) := X"0440000D";
        ram_buffer(54373) := X"00000000";
        ram_buffer(54374) := X"AFC00020";
        ram_buffer(54375) := X"8FC20020";
        ram_buffer(54376) := X"00000000";
        ram_buffer(54377) := X"AFC2001C";
        ram_buffer(54378) := X"8FC20038";
        ram_buffer(54379) := X"00000000";
        ram_buffer(54380) := X"AFC20028";
        ram_buffer(54381) := X"8FC20028";
        ram_buffer(54382) := X"00000000";
        ram_buffer(54383) := X"AFC20024";
        ram_buffer(54384) := X"1000000C";
        ram_buffer(54385) := X"00000000";
        ram_buffer(54386) := X"8FC20038";
        ram_buffer(54387) := X"00000000";
        ram_buffer(54388) := X"00021023";
        ram_buffer(54389) := X"AFC20020";
        ram_buffer(54390) := X"8FC20020";
        ram_buffer(54391) := X"00000000";
        ram_buffer(54392) := X"AFC2001C";
        ram_buffer(54393) := X"AFC00028";
        ram_buffer(54394) := X"8FC20028";
        ram_buffer(54395) := X"00000000";
        ram_buffer(54396) := X"AFC20024";
        ram_buffer(54397) := X"8FC200B0";
        ram_buffer(54398) := X"00000000";
        ram_buffer(54399) := X"04400008";
        ram_buffer(54400) := X"00000000";
        ram_buffer(54401) := X"8FC200B0";
        ram_buffer(54402) := X"8FC3001C";
        ram_buffer(54403) := X"00000000";
        ram_buffer(54404) := X"00621021";
        ram_buffer(54405) := X"AFC2001C";
        ram_buffer(54406) := X"10000006";
        ram_buffer(54407) := X"00000000";
        ram_buffer(54408) := X"8FC200B0";
        ram_buffer(54409) := X"8FC30024";
        ram_buffer(54410) := X"00000000";
        ram_buffer(54411) := X"00621023";
        ram_buffer(54412) := X"AFC20024";
        ram_buffer(54413) := X"8FC2001C";
        ram_buffer(54414) := X"00000000";
        ram_buffer(54415) := X"AFC2002C";
        ram_buffer(54416) := X"24020001";
        ram_buffer(54417) := X"AFC2008C";
        ram_buffer(54418) := X"AFC00090";
        ram_buffer(54419) := X"8FC300B0";
        ram_buffer(54420) := X"8FC20018";
        ram_buffer(54421) := X"00000000";
        ram_buffer(54422) := X"00621023";
        ram_buffer(54423) := X"AFC20048";
        ram_buffer(54424) := X"8FC300B4";
        ram_buffer(54425) := X"8FC20048";
        ram_buffer(54426) := X"00000000";
        ram_buffer(54427) := X"00621021";
        ram_buffer(54428) := X"2442FFFF";
        ram_buffer(54429) := X"AFC20044";
        ram_buffer(54430) := X"8FC200B4";
        ram_buffer(54431) := X"24030036";
        ram_buffer(54432) := X"00621023";
        ram_buffer(54433) := X"AFC20048";
        ram_buffer(54434) := X"8FC20044";
        ram_buffer(54435) := X"00000000";
        ram_buffer(54436) := X"2842FC02";
        ram_buffer(54437) := X"1040001E";
        ram_buffer(54438) := X"00000000";
        ram_buffer(54439) := X"2403FC02";
        ram_buffer(54440) := X"8FC20044";
        ram_buffer(54441) := X"00000000";
        ram_buffer(54442) := X"00621023";
        ram_buffer(54443) := X"AFC20044";
        ram_buffer(54444) := X"8FC30048";
        ram_buffer(54445) := X"8FC20044";
        ram_buffer(54446) := X"00000000";
        ram_buffer(54447) := X"00621023";
        ram_buffer(54448) := X"AFC20048";
        ram_buffer(54449) := X"8FC20044";
        ram_buffer(54450) := X"00000000";
        ram_buffer(54451) := X"28420020";
        ram_buffer(54452) := X"10400008";
        ram_buffer(54453) := X"00000000";
        ram_buffer(54454) := X"8FC3008C";
        ram_buffer(54455) := X"8FC20044";
        ram_buffer(54456) := X"00000000";
        ram_buffer(54457) := X"00431004";
        ram_buffer(54458) := X"AFC2008C";
        ram_buffer(54459) := X"10000008";
        ram_buffer(54460) := X"00000000";
        ram_buffer(54461) := X"8FC20044";
        ram_buffer(54462) := X"00000000";
        ram_buffer(54463) := X"2442FFE0";
        ram_buffer(54464) := X"8FC3008C";
        ram_buffer(54465) := X"00000000";
        ram_buffer(54466) := X"00431004";
        ram_buffer(54467) := X"AFC20090";
        ram_buffer(54468) := X"8FC3001C";
        ram_buffer(54469) := X"8FC20048";
        ram_buffer(54470) := X"00000000";
        ram_buffer(54471) := X"00621021";
        ram_buffer(54472) := X"AFC2001C";
        ram_buffer(54473) := X"8FC30024";
        ram_buffer(54474) := X"8FC20048";
        ram_buffer(54475) := X"00000000";
        ram_buffer(54476) := X"00621021";
        ram_buffer(54477) := X"AFC20024";
        ram_buffer(54478) := X"8FC30024";
        ram_buffer(54479) := X"8FC20018";
        ram_buffer(54480) := X"00000000";
        ram_buffer(54481) := X"00621021";
        ram_buffer(54482) := X"AFC20024";
        ram_buffer(54483) := X"8FC3001C";
        ram_buffer(54484) := X"8FC20024";
        ram_buffer(54485) := X"00000000";
        ram_buffer(54486) := X"0062202A";
        ram_buffer(54487) := X"10800002";
        ram_buffer(54488) := X"00000000";
        ram_buffer(54489) := X"00601021";
        ram_buffer(54490) := X"AFC20044";
        ram_buffer(54491) := X"8FC30044";
        ram_buffer(54492) := X"8FC2002C";
        ram_buffer(54493) := X"00000000";
        ram_buffer(54494) := X"0043102A";
        ram_buffer(54495) := X"10400004";
        ram_buffer(54496) := X"00000000";
        ram_buffer(54497) := X"8FC2002C";
        ram_buffer(54498) := X"00000000";
        ram_buffer(54499) := X"AFC20044";
        ram_buffer(54500) := X"8FC20044";
        ram_buffer(54501) := X"00000000";
        ram_buffer(54502) := X"18400010";
        ram_buffer(54503) := X"00000000";
        ram_buffer(54504) := X"8FC3001C";
        ram_buffer(54505) := X"8FC20044";
        ram_buffer(54506) := X"00000000";
        ram_buffer(54507) := X"00621023";
        ram_buffer(54508) := X"AFC2001C";
        ram_buffer(54509) := X"8FC30024";
        ram_buffer(54510) := X"8FC20044";
        ram_buffer(54511) := X"00000000";
        ram_buffer(54512) := X"00621023";
        ram_buffer(54513) := X"AFC20024";
        ram_buffer(54514) := X"8FC3002C";
        ram_buffer(54515) := X"8FC20044";
        ram_buffer(54516) := X"00000000";
        ram_buffer(54517) := X"00621023";
        ram_buffer(54518) := X"AFC2002C";
        ram_buffer(54519) := X"8FC20020";
        ram_buffer(54520) := X"00000000";
        ram_buffer(54521) := X"18400020";
        ram_buffer(54522) := X"00000000";
        ram_buffer(54523) := X"8FC60020";
        ram_buffer(54524) := X"8FC50084";
        ram_buffer(54525) := X"8FC40128";
        ram_buffer(54526) := X"0C02C138";
        ram_buffer(54527) := X"00000000";
        ram_buffer(54528) := X"AFC20084";
        ram_buffer(54529) := X"8FC20084";
        ram_buffer(54530) := X"00000000";
        ram_buffer(54531) := X"1040FDEA";
        ram_buffer(54532) := X"00000000";
        ram_buffer(54533) := X"8FC200D8";
        ram_buffer(54534) := X"00000000";
        ram_buffer(54535) := X"00403021";
        ram_buffer(54536) := X"8FC50084";
        ram_buffer(54537) := X"8FC40128";
        ram_buffer(54538) := X"0C02BFD8";
        ram_buffer(54539) := X"00000000";
        ram_buffer(54540) := X"AFC2009C";
        ram_buffer(54541) := X"8FC2009C";
        ram_buffer(54542) := X"00000000";
        ram_buffer(54543) := X"1040FDE1";
        ram_buffer(54544) := X"00000000";
        ram_buffer(54545) := X"8FC200D8";
        ram_buffer(54546) := X"00000000";
        ram_buffer(54547) := X"00402821";
        ram_buffer(54548) := X"8FC40128";
        ram_buffer(54549) := X"0C02BE10";
        ram_buffer(54550) := X"00000000";
        ram_buffer(54551) := X"8FC2009C";
        ram_buffer(54552) := X"00000000";
        ram_buffer(54553) := X"AFC200D8";
        ram_buffer(54554) := X"8FC2001C";
        ram_buffer(54555) := X"00000000";
        ram_buffer(54556) := X"1840000C";
        ram_buffer(54557) := X"00000000";
        ram_buffer(54558) := X"8FC200D8";
        ram_buffer(54559) := X"8FC6001C";
        ram_buffer(54560) := X"00402821";
        ram_buffer(54561) := X"8FC40128";
        ram_buffer(54562) := X"0C02C1BB";
        ram_buffer(54563) := X"00000000";
        ram_buffer(54564) := X"AFC200D8";
        ram_buffer(54565) := X"8FC200D8";
        ram_buffer(54566) := X"00000000";
        ram_buffer(54567) := X"1040FDCC";
        ram_buffer(54568) := X"00000000";
        ram_buffer(54569) := X"8FC20028";
        ram_buffer(54570) := X"00000000";
        ram_buffer(54571) := X"1840000B";
        ram_buffer(54572) := X"00000000";
        ram_buffer(54573) := X"8FC60028";
        ram_buffer(54574) := X"8FC5007C";
        ram_buffer(54575) := X"8FC40128";
        ram_buffer(54576) := X"0C02C138";
        ram_buffer(54577) := X"00000000";
        ram_buffer(54578) := X"AFC2007C";
        ram_buffer(54579) := X"8FC2007C";
        ram_buffer(54580) := X"00000000";
        ram_buffer(54581) := X"1040FDC1";
        ram_buffer(54582) := X"00000000";
        ram_buffer(54583) := X"8FC20024";
        ram_buffer(54584) := X"00000000";
        ram_buffer(54585) := X"1840000B";
        ram_buffer(54586) := X"00000000";
        ram_buffer(54587) := X"8FC60024";
        ram_buffer(54588) := X"8FC5007C";
        ram_buffer(54589) := X"8FC40128";
        ram_buffer(54590) := X"0C02C1BB";
        ram_buffer(54591) := X"00000000";
        ram_buffer(54592) := X"AFC2007C";
        ram_buffer(54593) := X"8FC2007C";
        ram_buffer(54594) := X"00000000";
        ram_buffer(54595) := X"1040FDB6";
        ram_buffer(54596) := X"00000000";
        ram_buffer(54597) := X"8FC2002C";
        ram_buffer(54598) := X"00000000";
        ram_buffer(54599) := X"1840000B";
        ram_buffer(54600) := X"00000000";
        ram_buffer(54601) := X"8FC6002C";
        ram_buffer(54602) := X"8FC50084";
        ram_buffer(54603) := X"8FC40128";
        ram_buffer(54604) := X"0C02C1BB";
        ram_buffer(54605) := X"00000000";
        ram_buffer(54606) := X"AFC20084";
        ram_buffer(54607) := X"8FC20084";
        ram_buffer(54608) := X"00000000";
        ram_buffer(54609) := X"1040FDAB";
        ram_buffer(54610) := X"00000000";
        ram_buffer(54611) := X"8FC200D8";
        ram_buffer(54612) := X"8FC6007C";
        ram_buffer(54613) := X"00402821";
        ram_buffer(54614) := X"8FC40128";
        ram_buffer(54615) := X"0C02C2CE";
        ram_buffer(54616) := X"00000000";
        ram_buffer(54617) := X"AFC20088";
        ram_buffer(54618) := X"8FC20088";
        ram_buffer(54619) := X"00000000";
        ram_buffer(54620) := X"1040FDA3";
        ram_buffer(54621) := X"00000000";
        ram_buffer(54622) := X"8FC20088";
        ram_buffer(54623) := X"00000000";
        ram_buffer(54624) := X"8C42000C";
        ram_buffer(54625) := X"00000000";
        ram_buffer(54626) := X"AFC200A0";
        ram_buffer(54627) := X"8FC20088";
        ram_buffer(54628) := X"00000000";
        ram_buffer(54629) := X"AC40000C";
        ram_buffer(54630) := X"8FC50084";
        ram_buffer(54631) := X"8FC40088";
        ram_buffer(54632) := X"0C02C26D";
        ram_buffer(54633) := X"00000000";
        ram_buffer(54634) := X"AFC20044";
        ram_buffer(54635) := X"8FC20044";
        ram_buffer(54636) := X"00000000";
        ram_buffer(54637) := X"04410032";
        ram_buffer(54638) := X"00000000";
        ram_buffer(54639) := X"8FC200A0";
        ram_buffer(54640) := X"00000000";
        ram_buffer(54641) := X"14400254";
        ram_buffer(54642) := X"00000000";
        ram_buffer(54643) := X"8FC200CC";
        ram_buffer(54644) := X"00000000";
        ram_buffer(54645) := X"14400250";
        ram_buffer(54646) := X"00000000";
        ram_buffer(54647) := X"8FC300C8";
        ram_buffer(54648) := X"3C02000F";
        ram_buffer(54649) := X"3442FFFF";
        ram_buffer(54650) := X"00621024";
        ram_buffer(54651) := X"1440024A";
        ram_buffer(54652) := X"00000000";
        ram_buffer(54653) := X"8FC300C8";
        ram_buffer(54654) := X"3C027FF0";
        ram_buffer(54655) := X"00621824";
        ram_buffer(54656) := X"3C0206B0";
        ram_buffer(54657) := X"34420001";
        ram_buffer(54658) := X"0062102B";
        ram_buffer(54659) := X"14400242";
        ram_buffer(54660) := X"00000000";
        ram_buffer(54661) := X"8FC20088";
        ram_buffer(54662) := X"00000000";
        ram_buffer(54663) := X"8C420014";
        ram_buffer(54664) := X"00000000";
        ram_buffer(54665) := X"14400008";
        ram_buffer(54666) := X"00000000";
        ram_buffer(54667) := X"8FC20088";
        ram_buffer(54668) := X"00000000";
        ram_buffer(54669) := X"8C420010";
        ram_buffer(54670) := X"00000000";
        ram_buffer(54671) := X"28420002";
        ram_buffer(54672) := X"1440022B";
        ram_buffer(54673) := X"00000000";
        ram_buffer(54674) := X"24060001";
        ram_buffer(54675) := X"8FC50088";
        ram_buffer(54676) := X"8FC40128";
        ram_buffer(54677) := X"0C02C1BB";
        ram_buffer(54678) := X"00000000";
        ram_buffer(54679) := X"AFC20088";
        ram_buffer(54680) := X"8FC50084";
        ram_buffer(54681) := X"8FC40088";
        ram_buffer(54682) := X"0C02C26D";
        ram_buffer(54683) := X"00000000";
        ram_buffer(54684) := X"18400222";
        ram_buffer(54685) := X"00000000";
        ram_buffer(54686) := X"10000049";
        ram_buffer(54687) := X"00000000";
        ram_buffer(54688) := X"8FC20044";
        ram_buffer(54689) := X"00000000";
        ram_buffer(54690) := X"144000B7";
        ram_buffer(54691) := X"00000000";
        ram_buffer(54692) := X"8FC200A0";
        ram_buffer(54693) := X"00000000";
        ram_buffer(54694) := X"10400037";
        ram_buffer(54695) := X"00000000";
        ram_buffer(54696) := X"8FC300C8";
        ram_buffer(54697) := X"3C02000F";
        ram_buffer(54698) := X"3442FFFF";
        ram_buffer(54699) := X"00621824";
        ram_buffer(54700) := X"3C02000F";
        ram_buffer(54701) := X"3442FFFF";
        ram_buffer(54702) := X"14620060";
        ram_buffer(54703) := X"00000000";
        ram_buffer(54704) := X"8FC300CC";
        ram_buffer(54705) := X"8FC20018";
        ram_buffer(54706) := X"00000000";
        ram_buffer(54707) := X"10400014";
        ram_buffer(54708) := X"00000000";
        ram_buffer(54709) := X"8FC400C8";
        ram_buffer(54710) := X"3C027FF0";
        ram_buffer(54711) := X"00821024";
        ram_buffer(54712) := X"AFC20074";
        ram_buffer(54713) := X"8FC40074";
        ram_buffer(54714) := X"3C0206A0";
        ram_buffer(54715) := X"34420001";
        ram_buffer(54716) := X"0082102B";
        ram_buffer(54717) := X"1040000A";
        ram_buffer(54718) := X"00000000";
        ram_buffer(54719) := X"8FC20074";
        ram_buffer(54720) := X"00000000";
        ram_buffer(54721) := X"00021502";
        ram_buffer(54722) := X"2404006B";
        ram_buffer(54723) := X"00821023";
        ram_buffer(54724) := X"2404FFFF";
        ram_buffer(54725) := X"00441004";
        ram_buffer(54726) := X"10000002";
        ram_buffer(54727) := X"00000000";
        ram_buffer(54728) := X"2402FFFF";
        ram_buffer(54729) := X"14620045";
        ram_buffer(54730) := X"00000000";
        ram_buffer(54731) := X"8FC300C8";
        ram_buffer(54732) := X"3C027FEF";
        ram_buffer(54733) := X"3442FFFF";
        ram_buffer(54734) := X"14620005";
        ram_buffer(54735) := X"00000000";
        ram_buffer(54736) := X"8FC300CC";
        ram_buffer(54737) := X"2402FFFF";
        ram_buffer(54738) := X"1062FD30";
        ram_buffer(54739) := X"00000000";
        ram_buffer(54740) := X"8FC300C8";
        ram_buffer(54741) := X"3C027FF0";
        ram_buffer(54742) := X"00621824";
        ram_buffer(54743) := X"3C020010";
        ram_buffer(54744) := X"00621021";
        ram_buffer(54745) := X"AFC200C8";
        ram_buffer(54746) := X"AFC000CC";
        ram_buffer(54747) := X"AFC000A0";
        ram_buffer(54748) := X"100001E9";
        ram_buffer(54749) := X"00000000";
        ram_buffer(54750) := X"8FC300C8";
        ram_buffer(54751) := X"3C02000F";
        ram_buffer(54752) := X"3442FFFF";
        ram_buffer(54753) := X"00621024";
        ram_buffer(54754) := X"1440002C";
        ram_buffer(54755) := X"00000000";
        ram_buffer(54756) := X"8FC200CC";
        ram_buffer(54757) := X"00000000";
        ram_buffer(54758) := X"14400028";
        ram_buffer(54759) := X"00000000";
        ram_buffer(54760) := X"8FC20018";
        ram_buffer(54761) := X"00000000";
        ram_buffer(54762) := X"10400015";
        ram_buffer(54763) := X"00000000";
        ram_buffer(54764) := X"8FC200C8";
        ram_buffer(54765) := X"00000000";
        ram_buffer(54766) := X"00401821";
        ram_buffer(54767) := X"3C027FF0";
        ram_buffer(54768) := X"00621024";
        ram_buffer(54769) := X"AFC20070";
        ram_buffer(54770) := X"8FC30070";
        ram_buffer(54771) := X"3C0206B0";
        ram_buffer(54772) := X"34420001";
        ram_buffer(54773) := X"0062102B";
        ram_buffer(54774) := X"10400009";
        ram_buffer(54775) := X"00000000";
        ram_buffer(54776) := X"8FC30070";
        ram_buffer(54777) := X"3C020370";
        ram_buffer(54778) := X"34420001";
        ram_buffer(54779) := X"0062102B";
        ram_buffer(54780) := X"1440FE0E";
        ram_buffer(54781) := X"00000000";
        ram_buffer(54782) := X"100001C7";
        ram_buffer(54783) := X"00000000";
        ram_buffer(54784) := X"8FC300C8";
        ram_buffer(54785) := X"3C027FF0";
        ram_buffer(54786) := X"00621824";
        ram_buffer(54787) := X"3C02FFF0";
        ram_buffer(54788) := X"00621021";
        ram_buffer(54789) := X"AFC20070";
        ram_buffer(54790) := X"8FC30070";
        ram_buffer(54791) := X"3C02000F";
        ram_buffer(54792) := X"3442FFFF";
        ram_buffer(54793) := X"00621025";
        ram_buffer(54794) := X"AFC200C8";
        ram_buffer(54795) := X"2402FFFF";
        ram_buffer(54796) := X"AFC200CC";
        ram_buffer(54797) := X"100001B8";
        ram_buffer(54798) := X"00000000";
        ram_buffer(54799) := X"8FC20090";
        ram_buffer(54800) := X"00000000";
        ram_buffer(54801) := X"10400009";
        ram_buffer(54802) := X"00000000";
        ram_buffer(54803) := X"8FC300C8";
        ram_buffer(54804) := X"8FC20090";
        ram_buffer(54805) := X"00000000";
        ram_buffer(54806) := X"00621024";
        ram_buffer(54807) := X"14400009";
        ram_buffer(54808) := X"00000000";
        ram_buffer(54809) := X"100001AC";
        ram_buffer(54810) := X"00000000";
        ram_buffer(54811) := X"8FC300CC";
        ram_buffer(54812) := X"8FC2008C";
        ram_buffer(54813) := X"00000000";
        ram_buffer(54814) := X"00621024";
        ram_buffer(54815) := X"104001A2";
        ram_buffer(54816) := X"00000000";
        ram_buffer(54817) := X"8FC200A0";
        ram_buffer(54818) := X"00000000";
        ram_buffer(54819) := X"10400014";
        ram_buffer(54820) := X"00000000";
        ram_buffer(54821) := X"8FC60018";
        ram_buffer(54822) := X"8FC500CC";
        ram_buffer(54823) := X"8FC400C8";
        ram_buffer(54824) := X"0C02CE35";
        ram_buffer(54825) := X"00000000";
        ram_buffer(54826) := X"00602821";
        ram_buffer(54827) := X"00402021";
        ram_buffer(54828) := X"8FC300CC";
        ram_buffer(54829) := X"8FC200C8";
        ram_buffer(54830) := X"00A03821";
        ram_buffer(54831) := X"00803021";
        ram_buffer(54832) := X"00602821";
        ram_buffer(54833) := X"00402021";
        ram_buffer(54834) := X"0C0311FC";
        ram_buffer(54835) := X"00000000";
        ram_buffer(54836) := X"AFC300CC";
        ram_buffer(54837) := X"AFC200C8";
        ram_buffer(54838) := X"1000001C";
        ram_buffer(54839) := X"00000000";
        ram_buffer(54840) := X"8FC60018";
        ram_buffer(54841) := X"8FC500CC";
        ram_buffer(54842) := X"8FC400C8";
        ram_buffer(54843) := X"0C02CE35";
        ram_buffer(54844) := X"00000000";
        ram_buffer(54845) := X"00602821";
        ram_buffer(54846) := X"00402021";
        ram_buffer(54847) := X"8FC300CC";
        ram_buffer(54848) := X"8FC200C8";
        ram_buffer(54849) := X"00A03821";
        ram_buffer(54850) := X"00803021";
        ram_buffer(54851) := X"00602821";
        ram_buffer(54852) := X"00402021";
        ram_buffer(54853) := X"0C0318D3";
        ram_buffer(54854) := X"00000000";
        ram_buffer(54855) := X"AFC300CC";
        ram_buffer(54856) := X"AFC200C8";
        ram_buffer(54857) := X"8FC300CC";
        ram_buffer(54858) := X"8FC200C8";
        ram_buffer(54859) := X"00003821";
        ram_buffer(54860) := X"00003021";
        ram_buffer(54861) := X"00602821";
        ram_buffer(54862) := X"00402021";
        ram_buffer(54863) := X"0C03167F";
        ram_buffer(54864) := X"00000000";
        ram_buffer(54865) := X"1040FDBC";
        ram_buffer(54866) := X"00000000";
        ram_buffer(54867) := X"24030001";
        ram_buffer(54868) := X"8FC200A0";
        ram_buffer(54869) := X"00000000";
        ram_buffer(54870) := X"00621023";
        ram_buffer(54871) := X"AFC200A0";
        ram_buffer(54872) := X"1000016D";
        ram_buffer(54873) := X"00000000";
        ram_buffer(54874) := X"8FC50084";
        ram_buffer(54875) := X"8FC40088";
        ram_buffer(54876) := X"0C02C55B";
        ram_buffer(54877) := X"00000000";
        ram_buffer(54878) := X"AFC3006C";
        ram_buffer(54879) := X"AFC20068";
        ram_buffer(54880) := X"8F87815C";
        ram_buffer(54881) := X"8F868158";
        ram_buffer(54882) := X"8FC5006C";
        ram_buffer(54883) := X"8FC40068";
        ram_buffer(54884) := X"0C0316F7";
        ram_buffer(54885) := X"00000000";
        ram_buffer(54886) := X"1C40004A";
        ram_buffer(54887) := X"00000000";
        ram_buffer(54888) := X"8FC200A0";
        ram_buffer(54889) := X"00000000";
        ram_buffer(54890) := X"1040000B";
        ram_buffer(54891) := X"00000000";
        ram_buffer(54892) := X"8F838164";
        ram_buffer(54893) := X"8F828160";
        ram_buffer(54894) := X"AFC300C4";
        ram_buffer(54895) := X"AFC200C0";
        ram_buffer(54896) := X"8FC300C4";
        ram_buffer(54897) := X"8FC200C0";
        ram_buffer(54898) := X"AFC3006C";
        ram_buffer(54899) := X"AFC20068";
        ram_buffer(54900) := X"10000052";
        ram_buffer(54901) := X"00000000";
        ram_buffer(54902) := X"8FC200CC";
        ram_buffer(54903) := X"00000000";
        ram_buffer(54904) := X"14400007";
        ram_buffer(54905) := X"00000000";
        ram_buffer(54906) := X"8FC300C8";
        ram_buffer(54907) := X"3C02000F";
        ram_buffer(54908) := X"3442FFFF";
        ram_buffer(54909) := X"00621024";
        ram_buffer(54910) := X"10400013";
        ram_buffer(54911) := X"00000000";
        ram_buffer(54912) := X"8FC300CC";
        ram_buffer(54913) := X"24020001";
        ram_buffer(54914) := X"14620005";
        ram_buffer(54915) := X"00000000";
        ram_buffer(54916) := X"8FC200C8";
        ram_buffer(54917) := X"00000000";
        ram_buffer(54918) := X"1040FD8A";
        ram_buffer(54919) := X"00000000";
        ram_buffer(54920) := X"8F838164";
        ram_buffer(54921) := X"8F828160";
        ram_buffer(54922) := X"AFC3006C";
        ram_buffer(54923) := X"AFC20068";
        ram_buffer(54924) := X"8F83816C";
        ram_buffer(54925) := X"8F828168";
        ram_buffer(54926) := X"AFC300C4";
        ram_buffer(54927) := X"AFC200C0";
        ram_buffer(54928) := X"10000036";
        ram_buffer(54929) := X"00000000";
        ram_buffer(54930) := X"8F878164";
        ram_buffer(54931) := X"8F868160";
        ram_buffer(54932) := X"8FC5006C";
        ram_buffer(54933) := X"8FC40068";
        ram_buffer(54934) := X"0C0316F7";
        ram_buffer(54935) := X"00000000";
        ram_buffer(54936) := X"04410007";
        ram_buffer(54937) := X"00000000";
        ram_buffer(54938) := X"8F838174";
        ram_buffer(54939) := X"8F828170";
        ram_buffer(54940) := X"AFC3006C";
        ram_buffer(54941) := X"AFC20068";
        ram_buffer(54942) := X"10000009";
        ram_buffer(54943) := X"00000000";
        ram_buffer(54944) := X"8F878174";
        ram_buffer(54945) := X"8F868170";
        ram_buffer(54946) := X"8FC5006C";
        ram_buffer(54947) := X"8FC40068";
        ram_buffer(54948) := X"0C03174A";
        ram_buffer(54949) := X"00000000";
        ram_buffer(54950) := X"AFC3006C";
        ram_buffer(54951) := X"AFC20068";
        ram_buffer(54952) := X"8FC30068";
        ram_buffer(54953) := X"3C028000";
        ram_buffer(54954) := X"0062B026";
        ram_buffer(54955) := X"8FD7006C";
        ram_buffer(54956) := X"00000000";
        ram_buffer(54957) := X"AFD700C4";
        ram_buffer(54958) := X"AFD600C0";
        ram_buffer(54959) := X"10000017";
        ram_buffer(54960) := X"00000000";
        ram_buffer(54961) := X"8F878174";
        ram_buffer(54962) := X"8F868170";
        ram_buffer(54963) := X"8FC5006C";
        ram_buffer(54964) := X"8FC40068";
        ram_buffer(54965) := X"0C03174A";
        ram_buffer(54966) := X"00000000";
        ram_buffer(54967) := X"AFC3006C";
        ram_buffer(54968) := X"AFC20068";
        ram_buffer(54969) := X"8FC200A0";
        ram_buffer(54970) := X"00000000";
        ram_buffer(54971) := X"14400007";
        ram_buffer(54972) := X"00000000";
        ram_buffer(54973) := X"8FC30068";
        ram_buffer(54974) := X"3C028000";
        ram_buffer(54975) := X"00628026";
        ram_buffer(54976) := X"8FD1006C";
        ram_buffer(54977) := X"10000003";
        ram_buffer(54978) := X"00000000";
        ram_buffer(54979) := X"8FD1006C";
        ram_buffer(54980) := X"8FD00068";
        ram_buffer(54981) := X"AFD100C4";
        ram_buffer(54982) := X"AFD000C0";
        ram_buffer(54983) := X"8FC300C8";
        ram_buffer(54984) := X"3C027FF0";
        ram_buffer(54985) := X"00621024";
        ram_buffer(54986) := X"AFC20074";
        ram_buffer(54987) := X"8FC30074";
        ram_buffer(54988) := X"3C027FE0";
        ram_buffer(54989) := X"14620042";
        ram_buffer(54990) := X"00000000";
        ram_buffer(54991) := X"8FC300CC";
        ram_buffer(54992) := X"8FC200C8";
        ram_buffer(54993) := X"AFC300D4";
        ram_buffer(54994) := X"AFC200D0";
        ram_buffer(54995) := X"8FC300C8";
        ram_buffer(54996) := X"3C02FCB0";
        ram_buffer(54997) := X"00621021";
        ram_buffer(54998) := X"AFC200C8";
        ram_buffer(54999) := X"8FC300C4";
        ram_buffer(55000) := X"8FC200C0";
        ram_buffer(55001) := X"AFC300F4";
        ram_buffer(55002) := X"AFC200F0";
        ram_buffer(55003) := X"8FC300CC";
        ram_buffer(55004) := X"8FC200C8";
        ram_buffer(55005) := X"00602821";
        ram_buffer(55006) := X"00402021";
        ram_buffer(55007) := X"0C02C3B7";
        ram_buffer(55008) := X"00000000";
        ram_buffer(55009) := X"00603821";
        ram_buffer(55010) := X"00403021";
        ram_buffer(55011) := X"8FC500F4";
        ram_buffer(55012) := X"8FC400F0";
        ram_buffer(55013) := X"0C03174A";
        ram_buffer(55014) := X"00000000";
        ram_buffer(55015) := X"AFC300AC";
        ram_buffer(55016) := X"AFC200A8";
        ram_buffer(55017) := X"8FC300CC";
        ram_buffer(55018) := X"8FC200C8";
        ram_buffer(55019) := X"8FC700AC";
        ram_buffer(55020) := X"8FC600A8";
        ram_buffer(55021) := X"00602821";
        ram_buffer(55022) := X"00402021";
        ram_buffer(55023) := X"0C0311FC";
        ram_buffer(55024) := X"00000000";
        ram_buffer(55025) := X"AFC300CC";
        ram_buffer(55026) := X"AFC200C8";
        ram_buffer(55027) := X"8FC300C8";
        ram_buffer(55028) := X"3C027FF0";
        ram_buffer(55029) := X"00621824";
        ram_buffer(55030) := X"3C027CA0";
        ram_buffer(55031) := X"0062102B";
        ram_buffer(55032) := X"14400011";
        ram_buffer(55033) := X"00000000";
        ram_buffer(55034) := X"8FC300D0";
        ram_buffer(55035) := X"3C027FEF";
        ram_buffer(55036) := X"3442FFFF";
        ram_buffer(55037) := X"14620005";
        ram_buffer(55038) := X"00000000";
        ram_buffer(55039) := X"8FC300D4";
        ram_buffer(55040) := X"2402FFFF";
        ram_buffer(55041) := X"1062FC04";
        ram_buffer(55042) := X"00000000";
        ram_buffer(55043) := X"3C027FEF";
        ram_buffer(55044) := X"3442FFFF";
        ram_buffer(55045) := X"AFC200C8";
        ram_buffer(55046) := X"2402FFFF";
        ram_buffer(55047) := X"AFC200CC";
        ram_buffer(55048) := X"1000009F";
        ram_buffer(55049) := X"00000000";
        ram_buffer(55050) := X"8FC300C8";
        ram_buffer(55051) := X"3C020350";
        ram_buffer(55052) := X"00621021";
        ram_buffer(55053) := X"AFC200C8";
        ram_buffer(55054) := X"10000054";
        ram_buffer(55055) := X"00000000";
        ram_buffer(55056) := X"8FC20018";
        ram_buffer(55057) := X"00000000";
        ram_buffer(55058) := X"10400034";
        ram_buffer(55059) := X"00000000";
        ram_buffer(55060) := X"8FC30074";
        ram_buffer(55061) := X"3C0206A0";
        ram_buffer(55062) := X"34420001";
        ram_buffer(55063) := X"0062102B";
        ram_buffer(55064) := X"1040002E";
        ram_buffer(55065) := X"00000000";
        ram_buffer(55066) := X"8F87817C";
        ram_buffer(55067) := X"8F868178";
        ram_buffer(55068) := X"8FC5006C";
        ram_buffer(55069) := X"8FC40068";
        ram_buffer(55070) := X"0C0316F7";
        ram_buffer(55071) := X"00000000";
        ram_buffer(55072) := X"1C40001F";
        ram_buffer(55073) := X"00000000";
        ram_buffer(55074) := X"8FC5006C";
        ram_buffer(55075) := X"8FC40068";
        ram_buffer(55076) := X"0C031B5A";
        ram_buffer(55077) := X"00000000";
        ram_buffer(55078) := X"AFC20078";
        ram_buffer(55079) := X"8FC20078";
        ram_buffer(55080) := X"00000000";
        ram_buffer(55081) := X"14400003";
        ram_buffer(55082) := X"00000000";
        ram_buffer(55083) := X"24020001";
        ram_buffer(55084) := X"AFC20078";
        ram_buffer(55085) := X"8FC40078";
        ram_buffer(55086) := X"0C031BBD";
        ram_buffer(55087) := X"00000000";
        ram_buffer(55088) := X"AFC3006C";
        ram_buffer(55089) := X"AFC20068";
        ram_buffer(55090) := X"8FC200A0";
        ram_buffer(55091) := X"00000000";
        ram_buffer(55092) := X"14400007";
        ram_buffer(55093) := X"00000000";
        ram_buffer(55094) := X"8FC30068";
        ram_buffer(55095) := X"3C028000";
        ram_buffer(55096) := X"00629026";
        ram_buffer(55097) := X"8FD3006C";
        ram_buffer(55098) := X"10000003";
        ram_buffer(55099) := X"00000000";
        ram_buffer(55100) := X"8FD3006C";
        ram_buffer(55101) := X"8FD20068";
        ram_buffer(55102) := X"AFD300C4";
        ram_buffer(55103) := X"AFD200C0";
        ram_buffer(55104) := X"8FC300C0";
        ram_buffer(55105) := X"8FC20074";
        ram_buffer(55106) := X"00000000";
        ram_buffer(55107) := X"00621823";
        ram_buffer(55108) := X"3C0206B0";
        ram_buffer(55109) := X"00621021";
        ram_buffer(55110) := X"AFC200C0";
        ram_buffer(55111) := X"8FC300C4";
        ram_buffer(55112) := X"8FC200C0";
        ram_buffer(55113) := X"AFC300F4";
        ram_buffer(55114) := X"AFC200F0";
        ram_buffer(55115) := X"8FC300CC";
        ram_buffer(55116) := X"8FC200C8";
        ram_buffer(55117) := X"00602821";
        ram_buffer(55118) := X"00402021";
        ram_buffer(55119) := X"0C02C3B7";
        ram_buffer(55120) := X"00000000";
        ram_buffer(55121) := X"00603821";
        ram_buffer(55122) := X"00403021";
        ram_buffer(55123) := X"8FC500F4";
        ram_buffer(55124) := X"8FC400F0";
        ram_buffer(55125) := X"0C03174A";
        ram_buffer(55126) := X"00000000";
        ram_buffer(55127) := X"AFC300AC";
        ram_buffer(55128) := X"AFC200A8";
        ram_buffer(55129) := X"8FC300CC";
        ram_buffer(55130) := X"8FC200C8";
        ram_buffer(55131) := X"8FC700AC";
        ram_buffer(55132) := X"8FC600A8";
        ram_buffer(55133) := X"00602821";
        ram_buffer(55134) := X"00402021";
        ram_buffer(55135) := X"0C0311FC";
        ram_buffer(55136) := X"00000000";
        ram_buffer(55137) := X"AFC300CC";
        ram_buffer(55138) := X"AFC200C8";
        ram_buffer(55139) := X"8FC300C8";
        ram_buffer(55140) := X"3C027FF0";
        ram_buffer(55141) := X"00621024";
        ram_buffer(55142) := X"AFC20078";
        ram_buffer(55143) := X"8FC20018";
        ram_buffer(55144) := X"00000000";
        ram_buffer(55145) := X"1440003E";
        ram_buffer(55146) := X"00000000";
        ram_buffer(55147) := X"8FC30074";
        ram_buffer(55148) := X"8FC20078";
        ram_buffer(55149) := X"00000000";
        ram_buffer(55150) := X"14620039";
        ram_buffer(55151) := X"00000000";
        ram_buffer(55152) := X"8FC5006C";
        ram_buffer(55153) := X"8FC40068";
        ram_buffer(55154) := X"0C031B37";
        ram_buffer(55155) := X"00000000";
        ram_buffer(55156) := X"AFC20070";
        ram_buffer(55157) := X"8FC40070";
        ram_buffer(55158) := X"0C031B7C";
        ram_buffer(55159) := X"00000000";
        ram_buffer(55160) := X"00603821";
        ram_buffer(55161) := X"00403021";
        ram_buffer(55162) := X"8FC5006C";
        ram_buffer(55163) := X"8FC40068";
        ram_buffer(55164) := X"0C0318D3";
        ram_buffer(55165) := X"00000000";
        ram_buffer(55166) := X"AFC3006C";
        ram_buffer(55167) := X"AFC20068";
        ram_buffer(55168) := X"8FC200A0";
        ram_buffer(55169) := X"00000000";
        ram_buffer(55170) := X"1440000B";
        ram_buffer(55171) := X"00000000";
        ram_buffer(55172) := X"8FC200CC";
        ram_buffer(55173) := X"00000000";
        ram_buffer(55174) := X"14400007";
        ram_buffer(55175) := X"00000000";
        ram_buffer(55176) := X"8FC300C8";
        ram_buffer(55177) := X"3C02000F";
        ram_buffer(55178) := X"3442FFFF";
        ram_buffer(55179) := X"00621024";
        ram_buffer(55180) := X"10400013";
        ram_buffer(55181) := X"00000000";
        ram_buffer(55182) := X"8F878184";
        ram_buffer(55183) := X"8F868180";
        ram_buffer(55184) := X"8FC5006C";
        ram_buffer(55185) := X"8FC40068";
        ram_buffer(55186) := X"0C0316F7";
        ram_buffer(55187) := X"00000000";
        ram_buffer(55188) := X"04400031";
        ram_buffer(55189) := X"00000000";
        ram_buffer(55190) := X"8F87818C";
        ram_buffer(55191) := X"8F868188";
        ram_buffer(55192) := X"8FC5006C";
        ram_buffer(55193) := X"8FC40068";
        ram_buffer(55194) := X"0C0316AB";
        ram_buffer(55195) := X"00000000";
        ram_buffer(55196) := X"1C400029";
        ram_buffer(55197) := X"00000000";
        ram_buffer(55198) := X"10000009";
        ram_buffer(55199) := X"00000000";
        ram_buffer(55200) := X"8F878194";
        ram_buffer(55201) := X"8F868190";
        ram_buffer(55202) := X"8FC5006C";
        ram_buffer(55203) := X"8FC40068";
        ram_buffer(55204) := X"0C0316F7";
        ram_buffer(55205) := X"00000000";
        ram_buffer(55206) := X"0440001E";
        ram_buffer(55207) := X"00000000";
        ram_buffer(55208) := X"8FC200D8";
        ram_buffer(55209) := X"00000000";
        ram_buffer(55210) := X"00402821";
        ram_buffer(55211) := X"8FC40128";
        ram_buffer(55212) := X"0C02BE10";
        ram_buffer(55213) := X"00000000";
        ram_buffer(55214) := X"8FC5007C";
        ram_buffer(55215) := X"8FC40128";
        ram_buffer(55216) := X"0C02BE10";
        ram_buffer(55217) := X"00000000";
        ram_buffer(55218) := X"8FC50084";
        ram_buffer(55219) := X"8FC40128";
        ram_buffer(55220) := X"0C02BE10";
        ram_buffer(55221) := X"00000000";
        ram_buffer(55222) := X"8FC50088";
        ram_buffer(55223) := X"8FC40128";
        ram_buffer(55224) := X"0C02BE10";
        ram_buffer(55225) := X"00000000";
        ram_buffer(55226) := X"1000FC70";
        ram_buffer(55227) := X"00000000";
        ram_buffer(55228) := X"00000000";
        ram_buffer(55229) := X"10000008";
        ram_buffer(55230) := X"00000000";
        ram_buffer(55231) := X"00000000";
        ram_buffer(55232) := X"10000005";
        ram_buffer(55233) := X"00000000";
        ram_buffer(55234) := X"00000000";
        ram_buffer(55235) := X"10000002";
        ram_buffer(55236) := X"00000000";
        ram_buffer(55237) := X"00000000";
        ram_buffer(55238) := X"8FC20018";
        ram_buffer(55239) := X"00000000";
        ram_buffer(55240) := X"1040001B";
        ram_buffer(55241) := X"00000000";
        ram_buffer(55242) := X"3C023950";
        ram_buffer(55243) := X"AFC200D0";
        ram_buffer(55244) := X"AFC000D4";
        ram_buffer(55245) := X"8FC300CC";
        ram_buffer(55246) := X"8FC200C8";
        ram_buffer(55247) := X"8FC500D4";
        ram_buffer(55248) := X"8FC400D0";
        ram_buffer(55249) := X"00A03821";
        ram_buffer(55250) := X"00803021";
        ram_buffer(55251) := X"00602821";
        ram_buffer(55252) := X"00402021";
        ram_buffer(55253) := X"0C03174A";
        ram_buffer(55254) := X"00000000";
        ram_buffer(55255) := X"AFC300CC";
        ram_buffer(55256) := X"AFC200C8";
        ram_buffer(55257) := X"8FC200C8";
        ram_buffer(55258) := X"00000000";
        ram_buffer(55259) := X"14400008";
        ram_buffer(55260) := X"00000000";
        ram_buffer(55261) := X"8FC200CC";
        ram_buffer(55262) := X"00000000";
        ram_buffer(55263) := X"14400004";
        ram_buffer(55264) := X"00000000";
        ram_buffer(55265) := X"8FC20128";
        ram_buffer(55266) := X"24030022";
        ram_buffer(55267) := X"AC430000";
        ram_buffer(55268) := X"8FC200D8";
        ram_buffer(55269) := X"00000000";
        ram_buffer(55270) := X"00402821";
        ram_buffer(55271) := X"8FC40128";
        ram_buffer(55272) := X"0C02BE10";
        ram_buffer(55273) := X"00000000";
        ram_buffer(55274) := X"8FC5007C";
        ram_buffer(55275) := X"8FC40128";
        ram_buffer(55276) := X"0C02BE10";
        ram_buffer(55277) := X"00000000";
        ram_buffer(55278) := X"8FC50084";
        ram_buffer(55279) := X"8FC40128";
        ram_buffer(55280) := X"0C02BE10";
        ram_buffer(55281) := X"00000000";
        ram_buffer(55282) := X"8FC50080";
        ram_buffer(55283) := X"8FC40128";
        ram_buffer(55284) := X"0C02BE10";
        ram_buffer(55285) := X"00000000";
        ram_buffer(55286) := X"8FC50088";
        ram_buffer(55287) := X"8FC40128";
        ram_buffer(55288) := X"0C02BE10";
        ram_buffer(55289) := X"00000000";
        ram_buffer(55290) := X"10000011";
        ram_buffer(55291) := X"00000000";
        ram_buffer(55292) := X"00000000";
        ram_buffer(55293) := X"1000000E";
        ram_buffer(55294) := X"00000000";
        ram_buffer(55295) := X"00000000";
        ram_buffer(55296) := X"1000000B";
        ram_buffer(55297) := X"00000000";
        ram_buffer(55298) := X"00000000";
        ram_buffer(55299) := X"10000008";
        ram_buffer(55300) := X"00000000";
        ram_buffer(55301) := X"00000000";
        ram_buffer(55302) := X"10000005";
        ram_buffer(55303) := X"00000000";
        ram_buffer(55304) := X"00000000";
        ram_buffer(55305) := X"10000002";
        ram_buffer(55306) := X"00000000";
        ram_buffer(55307) := X"00000000";
        ram_buffer(55308) := X"8FC20130";
        ram_buffer(55309) := X"00000000";
        ram_buffer(55310) := X"10400005";
        ram_buffer(55311) := X"00000000";
        ram_buffer(55312) := X"8FC300B8";
        ram_buffer(55313) := X"8FC20130";
        ram_buffer(55314) := X"00000000";
        ram_buffer(55315) := X"AC430000";
        ram_buffer(55316) := X"8FC20060";
        ram_buffer(55317) := X"00000000";
        ram_buffer(55318) := X"10400008";
        ram_buffer(55319) := X"00000000";
        ram_buffer(55320) := X"8FC300CC";
        ram_buffer(55321) := X"8FC200C8";
        ram_buffer(55322) := X"3C048000";
        ram_buffer(55323) := X"0044A026";
        ram_buffer(55324) := X"0060A821";
        ram_buffer(55325) := X"10000003";
        ram_buffer(55326) := X"00000000";
        ram_buffer(55327) := X"8FD500CC";
        ram_buffer(55328) := X"8FD400C8";
        ram_buffer(55329) := X"02A01821";
        ram_buffer(55330) := X"02801021";
        ram_buffer(55331) := X"03C0E821";
        ram_buffer(55332) := X"8FBF0124";
        ram_buffer(55333) := X"8FBE0120";
        ram_buffer(55334) := X"8FB7011C";
        ram_buffer(55335) := X"8FB60118";
        ram_buffer(55336) := X"8FB50114";
        ram_buffer(55337) := X"8FB40110";
        ram_buffer(55338) := X"8FB3010C";
        ram_buffer(55339) := X"8FB20108";
        ram_buffer(55340) := X"8FB10104";
        ram_buffer(55341) := X"8FB00100";
        ram_buffer(55342) := X"27BD0128";
        ram_buffer(55343) := X"03E00008";
        ram_buffer(55344) := X"00000000";
        ram_buffer(55345) := X"27BDFFE8";
        ram_buffer(55346) := X"AFBF0014";
        ram_buffer(55347) := X"AFBE0010";
        ram_buffer(55348) := X"03A0F021";
        ram_buffer(55349) := X"AFC40018";
        ram_buffer(55350) := X"AFC5001C";
        ram_buffer(55351) := X"8F828098";
        ram_buffer(55352) := X"8FC6001C";
        ram_buffer(55353) := X"8FC50018";
        ram_buffer(55354) := X"00402021";
        ram_buffer(55355) := X"0C02CF1C";
        ram_buffer(55356) := X"00000000";
        ram_buffer(55357) := X"03C0E821";
        ram_buffer(55358) := X"8FBF0014";
        ram_buffer(55359) := X"8FBE0010";
        ram_buffer(55360) := X"27BD0018";
        ram_buffer(55361) := X"03E00008";
        ram_buffer(55362) := X"00000000";
        ram_buffer(55363) := X"27BDFFE0";
        ram_buffer(55364) := X"AFBF001C";
        ram_buffer(55365) := X"AFBE0018";
        ram_buffer(55366) := X"03A0F021";
        ram_buffer(55367) := X"AFC40020";
        ram_buffer(55368) := X"AFC50024";
        ram_buffer(55369) := X"8F828098";
        ram_buffer(55370) := X"8FC60024";
        ram_buffer(55371) := X"8FC50020";
        ram_buffer(55372) := X"00402021";
        ram_buffer(55373) := X"0C02CF1C";
        ram_buffer(55374) := X"00000000";
        ram_buffer(55375) := X"AFC30014";
        ram_buffer(55376) := X"AFC20010";
        ram_buffer(55377) := X"8FC50014";
        ram_buffer(55378) := X"8FC40010";
        ram_buffer(55379) := X"0C02CAED";
        ram_buffer(55380) := X"00000000";
        ram_buffer(55381) := X"14400006";
        ram_buffer(55382) := X"00000000";
        ram_buffer(55383) := X"00002021";
        ram_buffer(55384) := X"0C02CC22";
        ram_buffer(55385) := X"00000000";
        ram_buffer(55386) := X"10000005";
        ram_buffer(55387) := X"00000000";
        ram_buffer(55388) := X"8FC50014";
        ram_buffer(55389) := X"8FC40010";
        ram_buffer(55390) := X"0C031C96";
        ram_buffer(55391) := X"00000000";
        ram_buffer(55392) := X"03C0E821";
        ram_buffer(55393) := X"8FBF001C";
        ram_buffer(55394) := X"8FBE0018";
        ram_buffer(55395) := X"27BD0020";
        ram_buffer(55396) := X"03E00008";
        ram_buffer(55397) := X"00000000";
        ram_buffer(55398) := X"27BDFFE0";
        ram_buffer(55399) := X"AFBE001C";
        ram_buffer(55400) := X"AFB60018";
        ram_buffer(55401) := X"AFB50014";
        ram_buffer(55402) := X"AFB40010";
        ram_buffer(55403) := X"AFB3000C";
        ram_buffer(55404) := X"AFB20008";
        ram_buffer(55405) := X"AFB10004";
        ram_buffer(55406) := X"AFB00000";
        ram_buffer(55407) := X"03A0F021";
        ram_buffer(55408) := X"AFC40020";
        ram_buffer(55409) := X"AFC50024";
        ram_buffer(55410) := X"AFC60028";
        ram_buffer(55411) := X"AFC7002C";
        ram_buffer(55412) := X"8FD10024";
        ram_buffer(55413) := X"0000A821";
        ram_buffer(55414) := X"02201021";
        ram_buffer(55415) := X"24510001";
        ram_buffer(55416) := X"90420000";
        ram_buffer(55417) := X"00000000";
        ram_buffer(55418) := X"00408021";
        ram_buffer(55419) := X"8F838090";
        ram_buffer(55420) := X"02001021";
        ram_buffer(55421) := X"24420001";
        ram_buffer(55422) := X"00621021";
        ram_buffer(55423) := X"80420000";
        ram_buffer(55424) := X"00000000";
        ram_buffer(55425) := X"304200FF";
        ram_buffer(55426) := X"30420008";
        ram_buffer(55427) := X"1440FFF2";
        ram_buffer(55428) := X"00000000";
        ram_buffer(55429) := X"2402002D";
        ram_buffer(55430) := X"16020009";
        ram_buffer(55431) := X"00000000";
        ram_buffer(55432) := X"24150001";
        ram_buffer(55433) := X"02201021";
        ram_buffer(55434) := X"24510001";
        ram_buffer(55435) := X"90420000";
        ram_buffer(55436) := X"00000000";
        ram_buffer(55437) := X"00408021";
        ram_buffer(55438) := X"10000009";
        ram_buffer(55439) := X"00000000";
        ram_buffer(55440) := X"2402002B";
        ram_buffer(55441) := X"16020006";
        ram_buffer(55442) := X"00000000";
        ram_buffer(55443) := X"02201021";
        ram_buffer(55444) := X"24510001";
        ram_buffer(55445) := X"90420000";
        ram_buffer(55446) := X"00000000";
        ram_buffer(55447) := X"00408021";
        ram_buffer(55448) := X"8FC2002C";
        ram_buffer(55449) := X"00000000";
        ram_buffer(55450) := X"10400005";
        ram_buffer(55451) := X"00000000";
        ram_buffer(55452) := X"8FC3002C";
        ram_buffer(55453) := X"24020010";
        ram_buffer(55454) := X"14620013";
        ram_buffer(55455) := X"00000000";
        ram_buffer(55456) := X"24020030";
        ram_buffer(55457) := X"16020010";
        ram_buffer(55458) := X"00000000";
        ram_buffer(55459) := X"92230000";
        ram_buffer(55460) := X"24020078";
        ram_buffer(55461) := X"10620005";
        ram_buffer(55462) := X"00000000";
        ram_buffer(55463) := X"92230000";
        ram_buffer(55464) := X"24020058";
        ram_buffer(55465) := X"14620008";
        ram_buffer(55466) := X"00000000";
        ram_buffer(55467) := X"26220001";
        ram_buffer(55468) := X"90420000";
        ram_buffer(55469) := X"00000000";
        ram_buffer(55470) := X"00408021";
        ram_buffer(55471) := X"26310002";
        ram_buffer(55472) := X"24020010";
        ram_buffer(55473) := X"AFC2002C";
        ram_buffer(55474) := X"8FC2002C";
        ram_buffer(55475) := X"00000000";
        ram_buffer(55476) := X"14400009";
        ram_buffer(55477) := X"00000000";
        ram_buffer(55478) := X"24020030";
        ram_buffer(55479) := X"16020004";
        ram_buffer(55480) := X"00000000";
        ram_buffer(55481) := X"24020008";
        ram_buffer(55482) := X"10000002";
        ram_buffer(55483) := X"00000000";
        ram_buffer(55484) := X"2402000A";
        ram_buffer(55485) := X"AFC2002C";
        ram_buffer(55486) := X"12A00004";
        ram_buffer(55487) := X"00000000";
        ram_buffer(55488) := X"3C028000";
        ram_buffer(55489) := X"10000003";
        ram_buffer(55490) := X"00000000";
        ram_buffer(55491) := X"3C027FFF";
        ram_buffer(55492) := X"3442FFFF";
        ram_buffer(55493) := X"00409821";
        ram_buffer(55494) := X"8FC2002C";
        ram_buffer(55495) := X"00000000";
        ram_buffer(55496) := X"14400002";
        ram_buffer(55497) := X"0262001B";
        ram_buffer(55498) := X"0007000D";
        ram_buffer(55499) := X"00001010";
        ram_buffer(55500) := X"0040B021";
        ram_buffer(55501) := X"8FC2002C";
        ram_buffer(55502) := X"00000000";
        ram_buffer(55503) := X"14400002";
        ram_buffer(55504) := X"0262001B";
        ram_buffer(55505) := X"0007000D";
        ram_buffer(55506) := X"00001010";
        ram_buffer(55507) := X"00009812";
        ram_buffer(55508) := X"00009021";
        ram_buffer(55509) := X"0000A021";
        ram_buffer(55510) := X"8F838090";
        ram_buffer(55511) := X"02001021";
        ram_buffer(55512) := X"24420001";
        ram_buffer(55513) := X"00621021";
        ram_buffer(55514) := X"80420000";
        ram_buffer(55515) := X"00000000";
        ram_buffer(55516) := X"304200FF";
        ram_buffer(55517) := X"30420004";
        ram_buffer(55518) := X"10400004";
        ram_buffer(55519) := X"00000000";
        ram_buffer(55520) := X"2610FFD0";
        ram_buffer(55521) := X"1000001B";
        ram_buffer(55522) := X"00000000";
        ram_buffer(55523) := X"8F838090";
        ram_buffer(55524) := X"02001021";
        ram_buffer(55525) := X"24420001";
        ram_buffer(55526) := X"00621021";
        ram_buffer(55527) := X"80420000";
        ram_buffer(55528) := X"00000000";
        ram_buffer(55529) := X"304200FF";
        ram_buffer(55530) := X"30420003";
        ram_buffer(55531) := X"10400031";
        ram_buffer(55532) := X"00000000";
        ram_buffer(55533) := X"8F838090";
        ram_buffer(55534) := X"02001021";
        ram_buffer(55535) := X"24420001";
        ram_buffer(55536) := X"00621021";
        ram_buffer(55537) := X"80420000";
        ram_buffer(55538) := X"00000000";
        ram_buffer(55539) := X"304200FF";
        ram_buffer(55540) := X"30430003";
        ram_buffer(55541) := X"24020001";
        ram_buffer(55542) := X"14620004";
        ram_buffer(55543) := X"00000000";
        ram_buffer(55544) := X"24020037";
        ram_buffer(55545) := X"10000002";
        ram_buffer(55546) := X"00000000";
        ram_buffer(55547) := X"24020057";
        ram_buffer(55548) := X"02028023";
        ram_buffer(55549) := X"8FC2002C";
        ram_buffer(55550) := X"00000000";
        ram_buffer(55551) := X"0202102A";
        ram_buffer(55552) := X"1040001F";
        ram_buffer(55553) := X"00000000";
        ram_buffer(55554) := X"06800009";
        ram_buffer(55555) := X"00000000";
        ram_buffer(55556) := X"0272102B";
        ram_buffer(55557) := X"14400006";
        ram_buffer(55558) := X"00000000";
        ram_buffer(55559) := X"16530007";
        ram_buffer(55560) := X"00000000";
        ram_buffer(55561) := X"02D0102A";
        ram_buffer(55562) := X"10400004";
        ram_buffer(55563) := X"00000000";
        ram_buffer(55564) := X"2414FFFF";
        ram_buffer(55565) := X"10000008";
        ram_buffer(55566) := X"00000000";
        ram_buffer(55567) := X"24140001";
        ram_buffer(55568) := X"8FC2002C";
        ram_buffer(55569) := X"00000000";
        ram_buffer(55570) := X"02420018";
        ram_buffer(55571) := X"00009012";
        ram_buffer(55572) := X"02001021";
        ram_buffer(55573) := X"02429021";
        ram_buffer(55574) := X"02201021";
        ram_buffer(55575) := X"24510001";
        ram_buffer(55576) := X"90420000";
        ram_buffer(55577) := X"00000000";
        ram_buffer(55578) := X"00408021";
        ram_buffer(55579) := X"1000FFBA";
        ram_buffer(55580) := X"00000000";
        ram_buffer(55581) := X"00000000";
        ram_buffer(55582) := X"10000002";
        ram_buffer(55583) := X"00000000";
        ram_buffer(55584) := X"00000000";
        ram_buffer(55585) := X"0681000E";
        ram_buffer(55586) := X"00000000";
        ram_buffer(55587) := X"12A00004";
        ram_buffer(55588) := X"00000000";
        ram_buffer(55589) := X"3C028000";
        ram_buffer(55590) := X"10000003";
        ram_buffer(55591) := X"00000000";
        ram_buffer(55592) := X"3C027FFF";
        ram_buffer(55593) := X"3442FFFF";
        ram_buffer(55594) := X"00409021";
        ram_buffer(55595) := X"8FC20020";
        ram_buffer(55596) := X"24030022";
        ram_buffer(55597) := X"AC430000";
        ram_buffer(55598) := X"10000004";
        ram_buffer(55599) := X"00000000";
        ram_buffer(55600) := X"12A00002";
        ram_buffer(55601) := X"00000000";
        ram_buffer(55602) := X"00129023";
        ram_buffer(55603) := X"8FC20028";
        ram_buffer(55604) := X"00000000";
        ram_buffer(55605) := X"1040000A";
        ram_buffer(55606) := X"00000000";
        ram_buffer(55607) := X"12800004";
        ram_buffer(55608) := X"00000000";
        ram_buffer(55609) := X"2622FFFF";
        ram_buffer(55610) := X"10000002";
        ram_buffer(55611) := X"00000000";
        ram_buffer(55612) := X"8FC20024";
        ram_buffer(55613) := X"8FC30028";
        ram_buffer(55614) := X"00000000";
        ram_buffer(55615) := X"AC620000";
        ram_buffer(55616) := X"02401021";
        ram_buffer(55617) := X"03C0E821";
        ram_buffer(55618) := X"8FBE001C";
        ram_buffer(55619) := X"8FB60018";
        ram_buffer(55620) := X"8FB50014";
        ram_buffer(55621) := X"8FB40010";
        ram_buffer(55622) := X"8FB3000C";
        ram_buffer(55623) := X"8FB20008";
        ram_buffer(55624) := X"8FB10004";
        ram_buffer(55625) := X"8FB00000";
        ram_buffer(55626) := X"27BD0020";
        ram_buffer(55627) := X"03E00008";
        ram_buffer(55628) := X"00000000";
        ram_buffer(55629) := X"27BDFFE8";
        ram_buffer(55630) := X"AFBF0014";
        ram_buffer(55631) := X"AFBE0010";
        ram_buffer(55632) := X"03A0F021";
        ram_buffer(55633) := X"AFC40018";
        ram_buffer(55634) := X"AFC5001C";
        ram_buffer(55635) := X"AFC60020";
        ram_buffer(55636) := X"8F828098";
        ram_buffer(55637) := X"8FC70020";
        ram_buffer(55638) := X"8FC6001C";
        ram_buffer(55639) := X"8FC50018";
        ram_buffer(55640) := X"00402021";
        ram_buffer(55641) := X"0C02D866";
        ram_buffer(55642) := X"00000000";
        ram_buffer(55643) := X"03C0E821";
        ram_buffer(55644) := X"8FBF0014";
        ram_buffer(55645) := X"8FBE0010";
        ram_buffer(55646) := X"27BD0018";
        ram_buffer(55647) := X"03E00008";
        ram_buffer(55648) := X"00000000";
        ram_buffer(55649) := X"27BDFFB8";
        ram_buffer(55650) := X"AFBF0044";
        ram_buffer(55651) := X"AFBE0040";
        ram_buffer(55652) := X"AFB7003C";
        ram_buffer(55653) := X"AFB60038";
        ram_buffer(55654) := X"AFB50034";
        ram_buffer(55655) := X"AFB40030";
        ram_buffer(55656) := X"AFB3002C";
        ram_buffer(55657) := X"AFB20028";
        ram_buffer(55658) := X"AFB10024";
        ram_buffer(55659) := X"AFB00020";
        ram_buffer(55660) := X"03A0F021";
        ram_buffer(55661) := X"AFC40048";
        ram_buffer(55662) := X"AFC5004C";
        ram_buffer(55663) := X"AFC60050";
        ram_buffer(55664) := X"AFC70054";
        ram_buffer(55665) := X"8FD3004C";
        ram_buffer(55666) := X"AFC00010";
        ram_buffer(55667) := X"02601021";
        ram_buffer(55668) := X"24530001";
        ram_buffer(55669) := X"90420000";
        ram_buffer(55670) := X"00000000";
        ram_buffer(55671) := X"00409021";
        ram_buffer(55672) := X"8F838090";
        ram_buffer(55673) := X"02401021";
        ram_buffer(55674) := X"24420001";
        ram_buffer(55675) := X"00621021";
        ram_buffer(55676) := X"80420000";
        ram_buffer(55677) := X"00000000";
        ram_buffer(55678) := X"304200FF";
        ram_buffer(55679) := X"30420008";
        ram_buffer(55680) := X"1440FFF2";
        ram_buffer(55681) := X"00000000";
        ram_buffer(55682) := X"2402002D";
        ram_buffer(55683) := X"1642000A";
        ram_buffer(55684) := X"00000000";
        ram_buffer(55685) := X"24020001";
        ram_buffer(55686) := X"AFC20010";
        ram_buffer(55687) := X"02601021";
        ram_buffer(55688) := X"24530001";
        ram_buffer(55689) := X"90420000";
        ram_buffer(55690) := X"00000000";
        ram_buffer(55691) := X"00409021";
        ram_buffer(55692) := X"10000009";
        ram_buffer(55693) := X"00000000";
        ram_buffer(55694) := X"2402002B";
        ram_buffer(55695) := X"16420006";
        ram_buffer(55696) := X"00000000";
        ram_buffer(55697) := X"02601021";
        ram_buffer(55698) := X"24530001";
        ram_buffer(55699) := X"90420000";
        ram_buffer(55700) := X"00000000";
        ram_buffer(55701) := X"00409021";
        ram_buffer(55702) := X"8FC20054";
        ram_buffer(55703) := X"00000000";
        ram_buffer(55704) := X"10400005";
        ram_buffer(55705) := X"00000000";
        ram_buffer(55706) := X"8FC30054";
        ram_buffer(55707) := X"24020010";
        ram_buffer(55708) := X"14620013";
        ram_buffer(55709) := X"00000000";
        ram_buffer(55710) := X"24020030";
        ram_buffer(55711) := X"16420010";
        ram_buffer(55712) := X"00000000";
        ram_buffer(55713) := X"92630000";
        ram_buffer(55714) := X"24020078";
        ram_buffer(55715) := X"10620005";
        ram_buffer(55716) := X"00000000";
        ram_buffer(55717) := X"92630000";
        ram_buffer(55718) := X"24020058";
        ram_buffer(55719) := X"14620008";
        ram_buffer(55720) := X"00000000";
        ram_buffer(55721) := X"26620001";
        ram_buffer(55722) := X"90420000";
        ram_buffer(55723) := X"00000000";
        ram_buffer(55724) := X"00409021";
        ram_buffer(55725) := X"26730002";
        ram_buffer(55726) := X"24020010";
        ram_buffer(55727) := X"AFC20054";
        ram_buffer(55728) := X"8FC20054";
        ram_buffer(55729) := X"00000000";
        ram_buffer(55730) := X"14400009";
        ram_buffer(55731) := X"00000000";
        ram_buffer(55732) := X"24020030";
        ram_buffer(55733) := X"16420004";
        ram_buffer(55734) := X"00000000";
        ram_buffer(55735) := X"24020008";
        ram_buffer(55736) := X"10000002";
        ram_buffer(55737) := X"00000000";
        ram_buffer(55738) := X"2402000A";
        ram_buffer(55739) := X"AFC20054";
        ram_buffer(55740) := X"8FC20010";
        ram_buffer(55741) := X"00000000";
        ram_buffer(55742) := X"10400005";
        ram_buffer(55743) := X"00000000";
        ram_buffer(55744) := X"00001821";
        ram_buffer(55745) := X"3C028000";
        ram_buffer(55746) := X"10000004";
        ram_buffer(55747) := X"00000000";
        ram_buffer(55748) := X"2403FFFF";
        ram_buffer(55749) := X"3C027FFF";
        ram_buffer(55750) := X"3442FFFF";
        ram_buffer(55751) := X"0060A821";
        ram_buffer(55752) := X"0040A021";
        ram_buffer(55753) := X"8FC20054";
        ram_buffer(55754) := X"00000000";
        ram_buffer(55755) := X"00404821";
        ram_buffer(55756) := X"000217C3";
        ram_buffer(55757) := X"00404021";
        ram_buffer(55758) := X"01203821";
        ram_buffer(55759) := X"01003021";
        ram_buffer(55760) := X"02A02821";
        ram_buffer(55761) := X"02802021";
        ram_buffer(55762) := X"0C030BFE";
        ram_buffer(55763) := X"00000000";
        ram_buffer(55764) := X"AFC30014";
        ram_buffer(55765) := X"8FC20054";
        ram_buffer(55766) := X"00000000";
        ram_buffer(55767) := X"00408821";
        ram_buffer(55768) := X"000217C3";
        ram_buffer(55769) := X"00408021";
        ram_buffer(55770) := X"02203821";
        ram_buffer(55771) := X"02003021";
        ram_buffer(55772) := X"02A02821";
        ram_buffer(55773) := X"02802021";
        ram_buffer(55774) := X"0C030A67";
        ram_buffer(55775) := X"00000000";
        ram_buffer(55776) := X"0060A821";
        ram_buffer(55777) := X"0040A021";
        ram_buffer(55778) := X"00008821";
        ram_buffer(55779) := X"00008021";
        ram_buffer(55780) := X"00004021";
        ram_buffer(55781) := X"8F838090";
        ram_buffer(55782) := X"02401021";
        ram_buffer(55783) := X"24420001";
        ram_buffer(55784) := X"00621021";
        ram_buffer(55785) := X"80420000";
        ram_buffer(55786) := X"00000000";
        ram_buffer(55787) := X"304200FF";
        ram_buffer(55788) := X"30420004";
        ram_buffer(55789) := X"10400004";
        ram_buffer(55790) := X"00000000";
        ram_buffer(55791) := X"2652FFD0";
        ram_buffer(55792) := X"1000001B";
        ram_buffer(55793) := X"00000000";
        ram_buffer(55794) := X"8F838090";
        ram_buffer(55795) := X"02401021";
        ram_buffer(55796) := X"24420001";
        ram_buffer(55797) := X"00621021";
        ram_buffer(55798) := X"80420000";
        ram_buffer(55799) := X"00000000";
        ram_buffer(55800) := X"304200FF";
        ram_buffer(55801) := X"30420003";
        ram_buffer(55802) := X"1040005A";
        ram_buffer(55803) := X"00000000";
        ram_buffer(55804) := X"8F838090";
        ram_buffer(55805) := X"02401021";
        ram_buffer(55806) := X"24420001";
        ram_buffer(55807) := X"00621021";
        ram_buffer(55808) := X"80420000";
        ram_buffer(55809) := X"00000000";
        ram_buffer(55810) := X"304200FF";
        ram_buffer(55811) := X"30430003";
        ram_buffer(55812) := X"24020001";
        ram_buffer(55813) := X"14620004";
        ram_buffer(55814) := X"00000000";
        ram_buffer(55815) := X"24020037";
        ram_buffer(55816) := X"10000002";
        ram_buffer(55817) := X"00000000";
        ram_buffer(55818) := X"24020057";
        ram_buffer(55819) := X"02429023";
        ram_buffer(55820) := X"8FC20054";
        ram_buffer(55821) := X"00000000";
        ram_buffer(55822) := X"0242102A";
        ram_buffer(55823) := X"10400048";
        ram_buffer(55824) := X"00000000";
        ram_buffer(55825) := X"01001021";
        ram_buffer(55826) := X"04400015";
        ram_buffer(55827) := X"00000000";
        ram_buffer(55828) := X"0290102B";
        ram_buffer(55829) := X"14400012";
        ram_buffer(55830) := X"00000000";
        ram_buffer(55831) := X"02801021";
        ram_buffer(55832) := X"16020004";
        ram_buffer(55833) := X"00000000";
        ram_buffer(55834) := X"02B1102B";
        ram_buffer(55835) := X"1440000C";
        ram_buffer(55836) := X"00000000";
        ram_buffer(55837) := X"02801021";
        ram_buffer(55838) := X"1602000D";
        ram_buffer(55839) := X"00000000";
        ram_buffer(55840) := X"02A01021";
        ram_buffer(55841) := X"1622000A";
        ram_buffer(55842) := X"00000000";
        ram_buffer(55843) := X"8FC20014";
        ram_buffer(55844) := X"00000000";
        ram_buffer(55845) := X"0052102A";
        ram_buffer(55846) := X"10400005";
        ram_buffer(55847) := X"00000000";
        ram_buffer(55848) := X"2402FFFF";
        ram_buffer(55849) := X"00404021";
        ram_buffer(55850) := X"10000023";
        ram_buffer(55851) := X"00000000";
        ram_buffer(55852) := X"24020001";
        ram_buffer(55853) := X"00404021";
        ram_buffer(55854) := X"8FC20054";
        ram_buffer(55855) := X"00000000";
        ram_buffer(55856) := X"0040B821";
        ram_buffer(55857) := X"000217C3";
        ram_buffer(55858) := X"0040B021";
        ram_buffer(55859) := X"02170018";
        ram_buffer(55860) := X"00001012";
        ram_buffer(55861) := X"00000000";
        ram_buffer(55862) := X"00000000";
        ram_buffer(55863) := X"02D10018";
        ram_buffer(55864) := X"00001812";
        ram_buffer(55865) := X"00431021";
        ram_buffer(55866) := X"00000000";
        ram_buffer(55867) := X"02370019";
        ram_buffer(55868) := X"00008812";
        ram_buffer(55869) := X"00008010";
        ram_buffer(55870) := X"00501021";
        ram_buffer(55871) := X"00408021";
        ram_buffer(55872) := X"AFD2001C";
        ram_buffer(55873) := X"001217C3";
        ram_buffer(55874) := X"AFC20018";
        ram_buffer(55875) := X"8FC7001C";
        ram_buffer(55876) := X"8FC60018";
        ram_buffer(55877) := X"00E02021";
        ram_buffer(55878) := X"02241821";
        ram_buffer(55879) := X"0071202B";
        ram_buffer(55880) := X"00C02821";
        ram_buffer(55881) := X"02051021";
        ram_buffer(55882) := X"00822021";
        ram_buffer(55883) := X"00801021";
        ram_buffer(55884) := X"00608821";
        ram_buffer(55885) := X"00408021";
        ram_buffer(55886) := X"02601021";
        ram_buffer(55887) := X"24530001";
        ram_buffer(55888) := X"90420000";
        ram_buffer(55889) := X"00000000";
        ram_buffer(55890) := X"00409021";
        ram_buffer(55891) := X"1000FF91";
        ram_buffer(55892) := X"00000000";
        ram_buffer(55893) := X"00000000";
        ram_buffer(55894) := X"10000002";
        ram_buffer(55895) := X"00000000";
        ram_buffer(55896) := X"00000000";
        ram_buffer(55897) := X"01001021";
        ram_buffer(55898) := X"04410013";
        ram_buffer(55899) := X"00000000";
        ram_buffer(55900) := X"8FC20010";
        ram_buffer(55901) := X"00000000";
        ram_buffer(55902) := X"10400005";
        ram_buffer(55903) := X"00000000";
        ram_buffer(55904) := X"00001821";
        ram_buffer(55905) := X"3C028000";
        ram_buffer(55906) := X"10000004";
        ram_buffer(55907) := X"00000000";
        ram_buffer(55908) := X"2403FFFF";
        ram_buffer(55909) := X"3C027FFF";
        ram_buffer(55910) := X"3442FFFF";
        ram_buffer(55911) := X"00608821";
        ram_buffer(55912) := X"00408021";
        ram_buffer(55913) := X"8FC20048";
        ram_buffer(55914) := X"24030022";
        ram_buffer(55915) := X"AC430000";
        ram_buffer(55916) := X"1000000E";
        ram_buffer(55917) := X"00000000";
        ram_buffer(55918) := X"8FC20010";
        ram_buffer(55919) := X"00000000";
        ram_buffer(55920) := X"1040000A";
        ram_buffer(55921) := X"00000000";
        ram_buffer(55922) := X"00002821";
        ram_buffer(55923) := X"00002021";
        ram_buffer(55924) := X"00B11823";
        ram_buffer(55925) := X"00A3302B";
        ram_buffer(55926) := X"00901023";
        ram_buffer(55927) := X"00462023";
        ram_buffer(55928) := X"00801021";
        ram_buffer(55929) := X"00608821";
        ram_buffer(55930) := X"00408021";
        ram_buffer(55931) := X"8FC20050";
        ram_buffer(55932) := X"00000000";
        ram_buffer(55933) := X"1040000B";
        ram_buffer(55934) := X"00000000";
        ram_buffer(55935) := X"01001021";
        ram_buffer(55936) := X"10400004";
        ram_buffer(55937) := X"00000000";
        ram_buffer(55938) := X"2662FFFF";
        ram_buffer(55939) := X"10000002";
        ram_buffer(55940) := X"00000000";
        ram_buffer(55941) := X"8FC2004C";
        ram_buffer(55942) := X"8FC30050";
        ram_buffer(55943) := X"00000000";
        ram_buffer(55944) := X"AC620000";
        ram_buffer(55945) := X"02201821";
        ram_buffer(55946) := X"02001021";
        ram_buffer(55947) := X"03C0E821";
        ram_buffer(55948) := X"8FBF0044";
        ram_buffer(55949) := X"8FBE0040";
        ram_buffer(55950) := X"8FB7003C";
        ram_buffer(55951) := X"8FB60038";
        ram_buffer(55952) := X"8FB50034";
        ram_buffer(55953) := X"8FB40030";
        ram_buffer(55954) := X"8FB3002C";
        ram_buffer(55955) := X"8FB20028";
        ram_buffer(55956) := X"8FB10024";
        ram_buffer(55957) := X"8FB00020";
        ram_buffer(55958) := X"27BD0048";
        ram_buffer(55959) := X"03E00008";
        ram_buffer(55960) := X"00000000";
        ram_buffer(55961) := X"27BDFFE0";
        ram_buffer(55962) := X"AFBE001C";
        ram_buffer(55963) := X"AFB60018";
        ram_buffer(55964) := X"AFB50014";
        ram_buffer(55965) := X"AFB40010";
        ram_buffer(55966) := X"AFB3000C";
        ram_buffer(55967) := X"AFB20008";
        ram_buffer(55968) := X"AFB10004";
        ram_buffer(55969) := X"AFB00000";
        ram_buffer(55970) := X"03A0F021";
        ram_buffer(55971) := X"AFC40020";
        ram_buffer(55972) := X"AFC50024";
        ram_buffer(55973) := X"AFC60028";
        ram_buffer(55974) := X"AFC7002C";
        ram_buffer(55975) := X"8FD10024";
        ram_buffer(55976) := X"0000A021";
        ram_buffer(55977) := X"02201021";
        ram_buffer(55978) := X"24510001";
        ram_buffer(55979) := X"90420000";
        ram_buffer(55980) := X"00000000";
        ram_buffer(55981) := X"00408021";
        ram_buffer(55982) := X"8F838090";
        ram_buffer(55983) := X"02001021";
        ram_buffer(55984) := X"24420001";
        ram_buffer(55985) := X"00621021";
        ram_buffer(55986) := X"80420000";
        ram_buffer(55987) := X"00000000";
        ram_buffer(55988) := X"304200FF";
        ram_buffer(55989) := X"30420008";
        ram_buffer(55990) := X"1440FFF2";
        ram_buffer(55991) := X"00000000";
        ram_buffer(55992) := X"2402002D";
        ram_buffer(55993) := X"16020009";
        ram_buffer(55994) := X"00000000";
        ram_buffer(55995) := X"24140001";
        ram_buffer(55996) := X"02201021";
        ram_buffer(55997) := X"24510001";
        ram_buffer(55998) := X"90420000";
        ram_buffer(55999) := X"00000000";
        ram_buffer(56000) := X"00408021";
        ram_buffer(56001) := X"10000009";
        ram_buffer(56002) := X"00000000";
        ram_buffer(56003) := X"2402002B";
        ram_buffer(56004) := X"16020006";
        ram_buffer(56005) := X"00000000";
        ram_buffer(56006) := X"02201021";
        ram_buffer(56007) := X"24510001";
        ram_buffer(56008) := X"90420000";
        ram_buffer(56009) := X"00000000";
        ram_buffer(56010) := X"00408021";
        ram_buffer(56011) := X"8FC2002C";
        ram_buffer(56012) := X"00000000";
        ram_buffer(56013) := X"10400005";
        ram_buffer(56014) := X"00000000";
        ram_buffer(56015) := X"8FC3002C";
        ram_buffer(56016) := X"24020010";
        ram_buffer(56017) := X"14620013";
        ram_buffer(56018) := X"00000000";
        ram_buffer(56019) := X"24020030";
        ram_buffer(56020) := X"16020010";
        ram_buffer(56021) := X"00000000";
        ram_buffer(56022) := X"92230000";
        ram_buffer(56023) := X"24020078";
        ram_buffer(56024) := X"10620005";
        ram_buffer(56025) := X"00000000";
        ram_buffer(56026) := X"92230000";
        ram_buffer(56027) := X"24020058";
        ram_buffer(56028) := X"14620008";
        ram_buffer(56029) := X"00000000";
        ram_buffer(56030) := X"26220001";
        ram_buffer(56031) := X"90420000";
        ram_buffer(56032) := X"00000000";
        ram_buffer(56033) := X"00408021";
        ram_buffer(56034) := X"26310002";
        ram_buffer(56035) := X"24020010";
        ram_buffer(56036) := X"AFC2002C";
        ram_buffer(56037) := X"8FC2002C";
        ram_buffer(56038) := X"00000000";
        ram_buffer(56039) := X"14400009";
        ram_buffer(56040) := X"00000000";
        ram_buffer(56041) := X"24020030";
        ram_buffer(56042) := X"16020004";
        ram_buffer(56043) := X"00000000";
        ram_buffer(56044) := X"24020008";
        ram_buffer(56045) := X"10000002";
        ram_buffer(56046) := X"00000000";
        ram_buffer(56047) := X"2402000A";
        ram_buffer(56048) := X"AFC2002C";
        ram_buffer(56049) := X"8FC2002C";
        ram_buffer(56050) := X"2403FFFF";
        ram_buffer(56051) := X"14400002";
        ram_buffer(56052) := X"0062001B";
        ram_buffer(56053) := X"0007000D";
        ram_buffer(56054) := X"00001010";
        ram_buffer(56055) := X"0000A812";
        ram_buffer(56056) := X"8FC2002C";
        ram_buffer(56057) := X"2403FFFF";
        ram_buffer(56058) := X"14400002";
        ram_buffer(56059) := X"0062001B";
        ram_buffer(56060) := X"0007000D";
        ram_buffer(56061) := X"00001010";
        ram_buffer(56062) := X"0040B021";
        ram_buffer(56063) := X"00009021";
        ram_buffer(56064) := X"00009821";
        ram_buffer(56065) := X"8F838090";
        ram_buffer(56066) := X"02001021";
        ram_buffer(56067) := X"24420001";
        ram_buffer(56068) := X"00621021";
        ram_buffer(56069) := X"80420000";
        ram_buffer(56070) := X"00000000";
        ram_buffer(56071) := X"304200FF";
        ram_buffer(56072) := X"30420004";
        ram_buffer(56073) := X"10400004";
        ram_buffer(56074) := X"00000000";
        ram_buffer(56075) := X"2610FFD0";
        ram_buffer(56076) := X"1000001B";
        ram_buffer(56077) := X"00000000";
        ram_buffer(56078) := X"8F838090";
        ram_buffer(56079) := X"02001021";
        ram_buffer(56080) := X"24420001";
        ram_buffer(56081) := X"00621021";
        ram_buffer(56082) := X"80420000";
        ram_buffer(56083) := X"00000000";
        ram_buffer(56084) := X"304200FF";
        ram_buffer(56085) := X"30420003";
        ram_buffer(56086) := X"10400031";
        ram_buffer(56087) := X"00000000";
        ram_buffer(56088) := X"8F838090";
        ram_buffer(56089) := X"02001021";
        ram_buffer(56090) := X"24420001";
        ram_buffer(56091) := X"00621021";
        ram_buffer(56092) := X"80420000";
        ram_buffer(56093) := X"00000000";
        ram_buffer(56094) := X"304200FF";
        ram_buffer(56095) := X"30430003";
        ram_buffer(56096) := X"24020001";
        ram_buffer(56097) := X"14620004";
        ram_buffer(56098) := X"00000000";
        ram_buffer(56099) := X"24020037";
        ram_buffer(56100) := X"10000002";
        ram_buffer(56101) := X"00000000";
        ram_buffer(56102) := X"24020057";
        ram_buffer(56103) := X"02028023";
        ram_buffer(56104) := X"8FC2002C";
        ram_buffer(56105) := X"00000000";
        ram_buffer(56106) := X"0202102A";
        ram_buffer(56107) := X"1040001F";
        ram_buffer(56108) := X"00000000";
        ram_buffer(56109) := X"06600009";
        ram_buffer(56110) := X"00000000";
        ram_buffer(56111) := X"02B2102B";
        ram_buffer(56112) := X"14400006";
        ram_buffer(56113) := X"00000000";
        ram_buffer(56114) := X"16550007";
        ram_buffer(56115) := X"00000000";
        ram_buffer(56116) := X"02D0102A";
        ram_buffer(56117) := X"10400004";
        ram_buffer(56118) := X"00000000";
        ram_buffer(56119) := X"2413FFFF";
        ram_buffer(56120) := X"10000008";
        ram_buffer(56121) := X"00000000";
        ram_buffer(56122) := X"24130001";
        ram_buffer(56123) := X"8FC2002C";
        ram_buffer(56124) := X"00000000";
        ram_buffer(56125) := X"02420018";
        ram_buffer(56126) := X"00009012";
        ram_buffer(56127) := X"02001021";
        ram_buffer(56128) := X"02429021";
        ram_buffer(56129) := X"02201021";
        ram_buffer(56130) := X"24510001";
        ram_buffer(56131) := X"90420000";
        ram_buffer(56132) := X"00000000";
        ram_buffer(56133) := X"00408021";
        ram_buffer(56134) := X"1000FFBA";
        ram_buffer(56135) := X"00000000";
        ram_buffer(56136) := X"00000000";
        ram_buffer(56137) := X"10000002";
        ram_buffer(56138) := X"00000000";
        ram_buffer(56139) := X"00000000";
        ram_buffer(56140) := X"06610007";
        ram_buffer(56141) := X"00000000";
        ram_buffer(56142) := X"2412FFFF";
        ram_buffer(56143) := X"8FC20020";
        ram_buffer(56144) := X"24030022";
        ram_buffer(56145) := X"AC430000";
        ram_buffer(56146) := X"10000004";
        ram_buffer(56147) := X"00000000";
        ram_buffer(56148) := X"12800002";
        ram_buffer(56149) := X"00000000";
        ram_buffer(56150) := X"00129023";
        ram_buffer(56151) := X"8FC20028";
        ram_buffer(56152) := X"00000000";
        ram_buffer(56153) := X"1040000A";
        ram_buffer(56154) := X"00000000";
        ram_buffer(56155) := X"12600004";
        ram_buffer(56156) := X"00000000";
        ram_buffer(56157) := X"2622FFFF";
        ram_buffer(56158) := X"10000002";
        ram_buffer(56159) := X"00000000";
        ram_buffer(56160) := X"8FC20024";
        ram_buffer(56161) := X"8FC30028";
        ram_buffer(56162) := X"00000000";
        ram_buffer(56163) := X"AC620000";
        ram_buffer(56164) := X"02401021";
        ram_buffer(56165) := X"03C0E821";
        ram_buffer(56166) := X"8FBE001C";
        ram_buffer(56167) := X"8FB60018";
        ram_buffer(56168) := X"8FB50014";
        ram_buffer(56169) := X"8FB40010";
        ram_buffer(56170) := X"8FB3000C";
        ram_buffer(56171) := X"8FB20008";
        ram_buffer(56172) := X"8FB10004";
        ram_buffer(56173) := X"8FB00000";
        ram_buffer(56174) := X"27BD0020";
        ram_buffer(56175) := X"03E00008";
        ram_buffer(56176) := X"00000000";
        ram_buffer(56177) := X"27BDFFE8";
        ram_buffer(56178) := X"AFBF0014";
        ram_buffer(56179) := X"AFBE0010";
        ram_buffer(56180) := X"03A0F021";
        ram_buffer(56181) := X"AFC40018";
        ram_buffer(56182) := X"AFC5001C";
        ram_buffer(56183) := X"AFC60020";
        ram_buffer(56184) := X"8F828098";
        ram_buffer(56185) := X"8FC70020";
        ram_buffer(56186) := X"8FC6001C";
        ram_buffer(56187) := X"8FC50018";
        ram_buffer(56188) := X"00402021";
        ram_buffer(56189) := X"0C02DA99";
        ram_buffer(56190) := X"00000000";
        ram_buffer(56191) := X"03C0E821";
        ram_buffer(56192) := X"8FBF0014";
        ram_buffer(56193) := X"8FBE0010";
        ram_buffer(56194) := X"27BD0018";
        ram_buffer(56195) := X"03E00008";
        ram_buffer(56196) := X"00000000";
        ram_buffer(56197) := X"27BDFFB8";
        ram_buffer(56198) := X"AFBF0044";
        ram_buffer(56199) := X"AFBE0040";
        ram_buffer(56200) := X"AFB7003C";
        ram_buffer(56201) := X"AFB60038";
        ram_buffer(56202) := X"AFB50034";
        ram_buffer(56203) := X"AFB40030";
        ram_buffer(56204) := X"AFB3002C";
        ram_buffer(56205) := X"AFB20028";
        ram_buffer(56206) := X"AFB10024";
        ram_buffer(56207) := X"AFB00020";
        ram_buffer(56208) := X"03A0F021";
        ram_buffer(56209) := X"AFC40048";
        ram_buffer(56210) := X"AFC5004C";
        ram_buffer(56211) := X"AFC60050";
        ram_buffer(56212) := X"AFC70054";
        ram_buffer(56213) := X"8FD3004C";
        ram_buffer(56214) := X"AFC00010";
        ram_buffer(56215) := X"02601021";
        ram_buffer(56216) := X"24530001";
        ram_buffer(56217) := X"90420000";
        ram_buffer(56218) := X"00000000";
        ram_buffer(56219) := X"00409021";
        ram_buffer(56220) := X"8F838090";
        ram_buffer(56221) := X"02401021";
        ram_buffer(56222) := X"24420001";
        ram_buffer(56223) := X"00621021";
        ram_buffer(56224) := X"80420000";
        ram_buffer(56225) := X"00000000";
        ram_buffer(56226) := X"304200FF";
        ram_buffer(56227) := X"30420008";
        ram_buffer(56228) := X"1440FFF2";
        ram_buffer(56229) := X"00000000";
        ram_buffer(56230) := X"2402002D";
        ram_buffer(56231) := X"1642000A";
        ram_buffer(56232) := X"00000000";
        ram_buffer(56233) := X"24020001";
        ram_buffer(56234) := X"AFC20010";
        ram_buffer(56235) := X"02601021";
        ram_buffer(56236) := X"24530001";
        ram_buffer(56237) := X"90420000";
        ram_buffer(56238) := X"00000000";
        ram_buffer(56239) := X"00409021";
        ram_buffer(56240) := X"10000009";
        ram_buffer(56241) := X"00000000";
        ram_buffer(56242) := X"2402002B";
        ram_buffer(56243) := X"16420006";
        ram_buffer(56244) := X"00000000";
        ram_buffer(56245) := X"02601021";
        ram_buffer(56246) := X"24530001";
        ram_buffer(56247) := X"90420000";
        ram_buffer(56248) := X"00000000";
        ram_buffer(56249) := X"00409021";
        ram_buffer(56250) := X"8FC20054";
        ram_buffer(56251) := X"00000000";
        ram_buffer(56252) := X"10400005";
        ram_buffer(56253) := X"00000000";
        ram_buffer(56254) := X"8FC30054";
        ram_buffer(56255) := X"24020010";
        ram_buffer(56256) := X"14620013";
        ram_buffer(56257) := X"00000000";
        ram_buffer(56258) := X"24020030";
        ram_buffer(56259) := X"16420010";
        ram_buffer(56260) := X"00000000";
        ram_buffer(56261) := X"92630000";
        ram_buffer(56262) := X"24020078";
        ram_buffer(56263) := X"10620005";
        ram_buffer(56264) := X"00000000";
        ram_buffer(56265) := X"92630000";
        ram_buffer(56266) := X"24020058";
        ram_buffer(56267) := X"14620008";
        ram_buffer(56268) := X"00000000";
        ram_buffer(56269) := X"26620001";
        ram_buffer(56270) := X"90420000";
        ram_buffer(56271) := X"00000000";
        ram_buffer(56272) := X"00409021";
        ram_buffer(56273) := X"26730002";
        ram_buffer(56274) := X"24020010";
        ram_buffer(56275) := X"AFC20054";
        ram_buffer(56276) := X"8FC20054";
        ram_buffer(56277) := X"00000000";
        ram_buffer(56278) := X"14400009";
        ram_buffer(56279) := X"00000000";
        ram_buffer(56280) := X"24020030";
        ram_buffer(56281) := X"16420004";
        ram_buffer(56282) := X"00000000";
        ram_buffer(56283) := X"24020008";
        ram_buffer(56284) := X"10000002";
        ram_buffer(56285) := X"00000000";
        ram_buffer(56286) := X"2402000A";
        ram_buffer(56287) := X"AFC20054";
        ram_buffer(56288) := X"8FC20054";
        ram_buffer(56289) := X"00000000";
        ram_buffer(56290) := X"00404821";
        ram_buffer(56291) := X"000217C3";
        ram_buffer(56292) := X"00404021";
        ram_buffer(56293) := X"01203821";
        ram_buffer(56294) := X"01003021";
        ram_buffer(56295) := X"2405FFFF";
        ram_buffer(56296) := X"2404FFFF";
        ram_buffer(56297) := X"0C030A67";
        ram_buffer(56298) := X"00000000";
        ram_buffer(56299) := X"0060B821";
        ram_buffer(56300) := X"0040B021";
        ram_buffer(56301) := X"8FC20054";
        ram_buffer(56302) := X"00000000";
        ram_buffer(56303) := X"00408821";
        ram_buffer(56304) := X"000217C3";
        ram_buffer(56305) := X"00408021";
        ram_buffer(56306) := X"2403FFFF";
        ram_buffer(56307) := X"2402FFFF";
        ram_buffer(56308) := X"02203821";
        ram_buffer(56309) := X"02003021";
        ram_buffer(56310) := X"00602821";
        ram_buffer(56311) := X"00402021";
        ram_buffer(56312) := X"0C030BFE";
        ram_buffer(56313) := X"00000000";
        ram_buffer(56314) := X"00604821";
        ram_buffer(56315) := X"00008821";
        ram_buffer(56316) := X"00008021";
        ram_buffer(56317) := X"00004021";
        ram_buffer(56318) := X"8F838090";
        ram_buffer(56319) := X"02401021";
        ram_buffer(56320) := X"24420001";
        ram_buffer(56321) := X"00621021";
        ram_buffer(56322) := X"80420000";
        ram_buffer(56323) := X"00000000";
        ram_buffer(56324) := X"304200FF";
        ram_buffer(56325) := X"30420004";
        ram_buffer(56326) := X"10400004";
        ram_buffer(56327) := X"00000000";
        ram_buffer(56328) := X"2652FFD0";
        ram_buffer(56329) := X"1000001B";
        ram_buffer(56330) := X"00000000";
        ram_buffer(56331) := X"8F838090";
        ram_buffer(56332) := X"02401021";
        ram_buffer(56333) := X"24420001";
        ram_buffer(56334) := X"00621021";
        ram_buffer(56335) := X"80420000";
        ram_buffer(56336) := X"00000000";
        ram_buffer(56337) := X"304200FF";
        ram_buffer(56338) := X"30420003";
        ram_buffer(56339) := X"10400059";
        ram_buffer(56340) := X"00000000";
        ram_buffer(56341) := X"8F838090";
        ram_buffer(56342) := X"02401021";
        ram_buffer(56343) := X"24420001";
        ram_buffer(56344) := X"00621021";
        ram_buffer(56345) := X"80420000";
        ram_buffer(56346) := X"00000000";
        ram_buffer(56347) := X"304200FF";
        ram_buffer(56348) := X"30430003";
        ram_buffer(56349) := X"24020001";
        ram_buffer(56350) := X"14620004";
        ram_buffer(56351) := X"00000000";
        ram_buffer(56352) := X"24020037";
        ram_buffer(56353) := X"10000002";
        ram_buffer(56354) := X"00000000";
        ram_buffer(56355) := X"24020057";
        ram_buffer(56356) := X"02429023";
        ram_buffer(56357) := X"8FC20054";
        ram_buffer(56358) := X"00000000";
        ram_buffer(56359) := X"0242102A";
        ram_buffer(56360) := X"10400047";
        ram_buffer(56361) := X"00000000";
        ram_buffer(56362) := X"01001021";
        ram_buffer(56363) := X"04400014";
        ram_buffer(56364) := X"00000000";
        ram_buffer(56365) := X"02D0102B";
        ram_buffer(56366) := X"14400011";
        ram_buffer(56367) := X"00000000";
        ram_buffer(56368) := X"02C01021";
        ram_buffer(56369) := X"16020004";
        ram_buffer(56370) := X"00000000";
        ram_buffer(56371) := X"02F1102B";
        ram_buffer(56372) := X"1440000B";
        ram_buffer(56373) := X"00000000";
        ram_buffer(56374) := X"02C01021";
        ram_buffer(56375) := X"1602000C";
        ram_buffer(56376) := X"00000000";
        ram_buffer(56377) := X"02E01021";
        ram_buffer(56378) := X"16220009";
        ram_buffer(56379) := X"00000000";
        ram_buffer(56380) := X"01201021";
        ram_buffer(56381) := X"0052102A";
        ram_buffer(56382) := X"10400005";
        ram_buffer(56383) := X"00000000";
        ram_buffer(56384) := X"2402FFFF";
        ram_buffer(56385) := X"00404021";
        ram_buffer(56386) := X"10000023";
        ram_buffer(56387) := X"00000000";
        ram_buffer(56388) := X"24020001";
        ram_buffer(56389) := X"00404021";
        ram_buffer(56390) := X"8FC20054";
        ram_buffer(56391) := X"00000000";
        ram_buffer(56392) := X"0040A821";
        ram_buffer(56393) := X"000217C3";
        ram_buffer(56394) := X"0040A021";
        ram_buffer(56395) := X"02150018";
        ram_buffer(56396) := X"00001012";
        ram_buffer(56397) := X"00000000";
        ram_buffer(56398) := X"00000000";
        ram_buffer(56399) := X"02910018";
        ram_buffer(56400) := X"00001812";
        ram_buffer(56401) := X"00431021";
        ram_buffer(56402) := X"00000000";
        ram_buffer(56403) := X"02350019";
        ram_buffer(56404) := X"00008812";
        ram_buffer(56405) := X"00008010";
        ram_buffer(56406) := X"00501021";
        ram_buffer(56407) := X"00408021";
        ram_buffer(56408) := X"AFD2001C";
        ram_buffer(56409) := X"001217C3";
        ram_buffer(56410) := X"AFC20018";
        ram_buffer(56411) := X"8FC7001C";
        ram_buffer(56412) := X"8FC60018";
        ram_buffer(56413) := X"00E02021";
        ram_buffer(56414) := X"02241821";
        ram_buffer(56415) := X"0071202B";
        ram_buffer(56416) := X"00C02821";
        ram_buffer(56417) := X"02051021";
        ram_buffer(56418) := X"00822021";
        ram_buffer(56419) := X"00801021";
        ram_buffer(56420) := X"00608821";
        ram_buffer(56421) := X"00408021";
        ram_buffer(56422) := X"02601021";
        ram_buffer(56423) := X"24530001";
        ram_buffer(56424) := X"90420000";
        ram_buffer(56425) := X"00000000";
        ram_buffer(56426) := X"00409021";
        ram_buffer(56427) := X"1000FF92";
        ram_buffer(56428) := X"00000000";
        ram_buffer(56429) := X"00000000";
        ram_buffer(56430) := X"10000002";
        ram_buffer(56431) := X"00000000";
        ram_buffer(56432) := X"00000000";
        ram_buffer(56433) := X"01001021";
        ram_buffer(56434) := X"04410008";
        ram_buffer(56435) := X"00000000";
        ram_buffer(56436) := X"2411FFFF";
        ram_buffer(56437) := X"2410FFFF";
        ram_buffer(56438) := X"8FC20048";
        ram_buffer(56439) := X"24030022";
        ram_buffer(56440) := X"AC430000";
        ram_buffer(56441) := X"1000000E";
        ram_buffer(56442) := X"00000000";
        ram_buffer(56443) := X"8FC20010";
        ram_buffer(56444) := X"00000000";
        ram_buffer(56445) := X"1040000A";
        ram_buffer(56446) := X"00000000";
        ram_buffer(56447) := X"00002821";
        ram_buffer(56448) := X"00002021";
        ram_buffer(56449) := X"00B11823";
        ram_buffer(56450) := X"00A3302B";
        ram_buffer(56451) := X"00901023";
        ram_buffer(56452) := X"00462023";
        ram_buffer(56453) := X"00801021";
        ram_buffer(56454) := X"00608821";
        ram_buffer(56455) := X"00408021";
        ram_buffer(56456) := X"8FC20050";
        ram_buffer(56457) := X"00000000";
        ram_buffer(56458) := X"1040000B";
        ram_buffer(56459) := X"00000000";
        ram_buffer(56460) := X"01001021";
        ram_buffer(56461) := X"10400004";
        ram_buffer(56462) := X"00000000";
        ram_buffer(56463) := X"2662FFFF";
        ram_buffer(56464) := X"10000002";
        ram_buffer(56465) := X"00000000";
        ram_buffer(56466) := X"8FC2004C";
        ram_buffer(56467) := X"8FC30050";
        ram_buffer(56468) := X"00000000";
        ram_buffer(56469) := X"AC620000";
        ram_buffer(56470) := X"02201821";
        ram_buffer(56471) := X"02001021";
        ram_buffer(56472) := X"03C0E821";
        ram_buffer(56473) := X"8FBF0044";
        ram_buffer(56474) := X"8FBE0040";
        ram_buffer(56475) := X"8FB7003C";
        ram_buffer(56476) := X"8FB60038";
        ram_buffer(56477) := X"8FB50034";
        ram_buffer(56478) := X"8FB40030";
        ram_buffer(56479) := X"8FB3002C";
        ram_buffer(56480) := X"8FB20028";
        ram_buffer(56481) := X"8FB10024";
        ram_buffer(56482) := X"8FB00020";
        ram_buffer(56483) := X"27BD0048";
        ram_buffer(56484) := X"03E00008";
        ram_buffer(56485) := X"00000000";
        ram_buffer(56486) := X"27BDFFC0";
        ram_buffer(56487) := X"AFBF003C";
        ram_buffer(56488) := X"AFBE0038";
        ram_buffer(56489) := X"AFB40034";
        ram_buffer(56490) := X"AFB30030";
        ram_buffer(56491) := X"AFB2002C";
        ram_buffer(56492) := X"AFB10028";
        ram_buffer(56493) := X"AFB00024";
        ram_buffer(56494) := X"03A0F021";
        ram_buffer(56495) := X"AFC40040";
        ram_buffer(56496) := X"AFC50044";
        ram_buffer(56497) := X"00C08021";
        ram_buffer(56498) := X"0000A021";
        ram_buffer(56499) := X"8E130000";
        ram_buffer(56500) := X"00008821";
        ram_buffer(56501) := X"8E020008";
        ram_buffer(56502) := X"00000000";
        ram_buffer(56503) := X"14400008";
        ram_buffer(56504) := X"00000000";
        ram_buffer(56505) := X"AE000004";
        ram_buffer(56506) := X"00001021";
        ram_buffer(56507) := X"100000DB";
        ram_buffer(56508) := X"00000000";
        ram_buffer(56509) := X"8E740000";
        ram_buffer(56510) := X"8E710004";
        ram_buffer(56511) := X"26730008";
        ram_buffer(56512) := X"1220FFFC";
        ram_buffer(56513) := X"00000000";
        ram_buffer(56514) := X"8FC20044";
        ram_buffer(56515) := X"00000000";
        ram_buffer(56516) := X"8C520008";
        ram_buffer(56517) := X"00000000";
        ram_buffer(56518) := X"02401021";
        ram_buffer(56519) := X"0222102B";
        ram_buffer(56520) := X"14400091";
        ram_buffer(56521) := X"00000000";
        ram_buffer(56522) := X"8FC20044";
        ram_buffer(56523) := X"00000000";
        ram_buffer(56524) := X"8442000C";
        ram_buffer(56525) := X"00000000";
        ram_buffer(56526) := X"3042FFFF";
        ram_buffer(56527) := X"30420480";
        ram_buffer(56528) := X"10400089";
        ram_buffer(56529) := X"00000000";
        ram_buffer(56530) := X"8FC20044";
        ram_buffer(56531) := X"00000000";
        ram_buffer(56532) := X"8C420000";
        ram_buffer(56533) := X"00000000";
        ram_buffer(56534) := X"00401821";
        ram_buffer(56535) := X"8FC20044";
        ram_buffer(56536) := X"00000000";
        ram_buffer(56537) := X"8C420010";
        ram_buffer(56538) := X"00000000";
        ram_buffer(56539) := X"00621023";
        ram_buffer(56540) := X"AFC20018";
        ram_buffer(56541) := X"8FC20044";
        ram_buffer(56542) := X"00000000";
        ram_buffer(56543) := X"8C430014";
        ram_buffer(56544) := X"00000000";
        ram_buffer(56545) := X"00601021";
        ram_buffer(56546) := X"00021040";
        ram_buffer(56547) := X"00431021";
        ram_buffer(56548) := X"00021FC2";
        ram_buffer(56549) := X"00621021";
        ram_buffer(56550) := X"00021043";
        ram_buffer(56551) := X"AFC20014";
        ram_buffer(56552) := X"8FC20018";
        ram_buffer(56553) := X"00000000";
        ram_buffer(56554) := X"00511021";
        ram_buffer(56555) := X"24430001";
        ram_buffer(56556) := X"8FC20014";
        ram_buffer(56557) := X"00000000";
        ram_buffer(56558) := X"0043102B";
        ram_buffer(56559) := X"10400006";
        ram_buffer(56560) := X"00000000";
        ram_buffer(56561) := X"8FC20018";
        ram_buffer(56562) := X"00000000";
        ram_buffer(56563) := X"00511021";
        ram_buffer(56564) := X"24420001";
        ram_buffer(56565) := X"AFC20014";
        ram_buffer(56566) := X"8FC20044";
        ram_buffer(56567) := X"00000000";
        ram_buffer(56568) := X"8442000C";
        ram_buffer(56569) := X"00000000";
        ram_buffer(56570) := X"3042FFFF";
        ram_buffer(56571) := X"30420400";
        ram_buffer(56572) := X"1040002A";
        ram_buffer(56573) := X"00000000";
        ram_buffer(56574) := X"8FC20014";
        ram_buffer(56575) := X"00000000";
        ram_buffer(56576) := X"00402821";
        ram_buffer(56577) := X"8FC40040";
        ram_buffer(56578) := X"0C027B8F";
        ram_buffer(56579) := X"00000000";
        ram_buffer(56580) := X"AFC20010";
        ram_buffer(56581) := X"8FC20010";
        ram_buffer(56582) := X"00000000";
        ram_buffer(56583) := X"14400006";
        ram_buffer(56584) := X"00000000";
        ram_buffer(56585) := X"8FC20040";
        ram_buffer(56586) := X"2403000C";
        ram_buffer(56587) := X"AC430000";
        ram_buffer(56588) := X"1000007D";
        ram_buffer(56589) := X"00000000";
        ram_buffer(56590) := X"8FC20044";
        ram_buffer(56591) := X"00000000";
        ram_buffer(56592) := X"8C420010";
        ram_buffer(56593) := X"8FC30018";
        ram_buffer(56594) := X"00000000";
        ram_buffer(56595) := X"00603021";
        ram_buffer(56596) := X"00402821";
        ram_buffer(56597) := X"8FC40010";
        ram_buffer(56598) := X"0C027F93";
        ram_buffer(56599) := X"00000000";
        ram_buffer(56600) := X"8FC20044";
        ram_buffer(56601) := X"00000000";
        ram_buffer(56602) := X"8443000C";
        ram_buffer(56603) := X"2402FB7F";
        ram_buffer(56604) := X"00621024";
        ram_buffer(56605) := X"00021400";
        ram_buffer(56606) := X"00021403";
        ram_buffer(56607) := X"34420080";
        ram_buffer(56608) := X"00021C00";
        ram_buffer(56609) := X"00031C03";
        ram_buffer(56610) := X"8FC20044";
        ram_buffer(56611) := X"00000000";
        ram_buffer(56612) := X"A443000C";
        ram_buffer(56613) := X"1000001D";
        ram_buffer(56614) := X"00000000";
        ram_buffer(56615) := X"8FC20044";
        ram_buffer(56616) := X"00000000";
        ram_buffer(56617) := X"8C420010";
        ram_buffer(56618) := X"8FC30014";
        ram_buffer(56619) := X"00000000";
        ram_buffer(56620) := X"00603021";
        ram_buffer(56621) := X"00402821";
        ram_buffer(56622) := X"8FC40040";
        ram_buffer(56623) := X"0C02C6A7";
        ram_buffer(56624) := X"00000000";
        ram_buffer(56625) := X"AFC20010";
        ram_buffer(56626) := X"8FC20010";
        ram_buffer(56627) := X"00000000";
        ram_buffer(56628) := X"1440000E";
        ram_buffer(56629) := X"00000000";
        ram_buffer(56630) := X"8FC20044";
        ram_buffer(56631) := X"00000000";
        ram_buffer(56632) := X"8C420010";
        ram_buffer(56633) := X"00000000";
        ram_buffer(56634) := X"00402821";
        ram_buffer(56635) := X"8FC40040";
        ram_buffer(56636) := X"0C027301";
        ram_buffer(56637) := X"00000000";
        ram_buffer(56638) := X"8FC20040";
        ram_buffer(56639) := X"2403000C";
        ram_buffer(56640) := X"AC430000";
        ram_buffer(56641) := X"10000048";
        ram_buffer(56642) := X"00000000";
        ram_buffer(56643) := X"8FC20044";
        ram_buffer(56644) := X"8FC30010";
        ram_buffer(56645) := X"00000000";
        ram_buffer(56646) := X"AC430010";
        ram_buffer(56647) := X"8FC20018";
        ram_buffer(56648) := X"8FC30010";
        ram_buffer(56649) := X"00000000";
        ram_buffer(56650) := X"00621821";
        ram_buffer(56651) := X"8FC20044";
        ram_buffer(56652) := X"00000000";
        ram_buffer(56653) := X"AC430000";
        ram_buffer(56654) := X"8FC20044";
        ram_buffer(56655) := X"8FC30014";
        ram_buffer(56656) := X"00000000";
        ram_buffer(56657) := X"AC430014";
        ram_buffer(56658) := X"02209021";
        ram_buffer(56659) := X"8FC30014";
        ram_buffer(56660) := X"8FC20018";
        ram_buffer(56661) := X"00000000";
        ram_buffer(56662) := X"00621823";
        ram_buffer(56663) := X"8FC20044";
        ram_buffer(56664) := X"00000000";
        ram_buffer(56665) := X"AC430008";
        ram_buffer(56666) := X"02401021";
        ram_buffer(56667) := X"0222102B";
        ram_buffer(56668) := X"10400002";
        ram_buffer(56669) := X"00000000";
        ram_buffer(56670) := X"02209021";
        ram_buffer(56671) := X"8FC20044";
        ram_buffer(56672) := X"00000000";
        ram_buffer(56673) := X"8C420000";
        ram_buffer(56674) := X"02401821";
        ram_buffer(56675) := X"00603021";
        ram_buffer(56676) := X"02802821";
        ram_buffer(56677) := X"00402021";
        ram_buffer(56678) := X"0C02BCED";
        ram_buffer(56679) := X"00000000";
        ram_buffer(56680) := X"8FC20044";
        ram_buffer(56681) := X"00000000";
        ram_buffer(56682) := X"8C420008";
        ram_buffer(56683) := X"00000000";
        ram_buffer(56684) := X"00521823";
        ram_buffer(56685) := X"8FC20044";
        ram_buffer(56686) := X"00000000";
        ram_buffer(56687) := X"AC430008";
        ram_buffer(56688) := X"8FC20044";
        ram_buffer(56689) := X"00000000";
        ram_buffer(56690) := X"8C420000";
        ram_buffer(56691) := X"02401821";
        ram_buffer(56692) := X"00431821";
        ram_buffer(56693) := X"8FC20044";
        ram_buffer(56694) := X"00000000";
        ram_buffer(56695) := X"AC430000";
        ram_buffer(56696) := X"02209021";
        ram_buffer(56697) := X"02401021";
        ram_buffer(56698) := X"0282A021";
        ram_buffer(56699) := X"02401021";
        ram_buffer(56700) := X"02228823";
        ram_buffer(56701) := X"8E020008";
        ram_buffer(56702) := X"02401821";
        ram_buffer(56703) := X"00431023";
        ram_buffer(56704) := X"AE020008";
        ram_buffer(56705) := X"8E020008";
        ram_buffer(56706) := X"00000000";
        ram_buffer(56707) := X"1440FF3C";
        ram_buffer(56708) := X"00000000";
        ram_buffer(56709) := X"AE000008";
        ram_buffer(56710) := X"AE000004";
        ram_buffer(56711) := X"00001021";
        ram_buffer(56712) := X"1000000E";
        ram_buffer(56713) := X"00000000";
        ram_buffer(56714) := X"8FC20044";
        ram_buffer(56715) := X"00000000";
        ram_buffer(56716) := X"8442000C";
        ram_buffer(56717) := X"00000000";
        ram_buffer(56718) := X"34420040";
        ram_buffer(56719) := X"00021C00";
        ram_buffer(56720) := X"00031C03";
        ram_buffer(56721) := X"8FC20044";
        ram_buffer(56722) := X"00000000";
        ram_buffer(56723) := X"A443000C";
        ram_buffer(56724) := X"AE000008";
        ram_buffer(56725) := X"AE000004";
        ram_buffer(56726) := X"2402FFFF";
        ram_buffer(56727) := X"03C0E821";
        ram_buffer(56728) := X"8FBF003C";
        ram_buffer(56729) := X"8FBE0038";
        ram_buffer(56730) := X"8FB40034";
        ram_buffer(56731) := X"8FB30030";
        ram_buffer(56732) := X"8FB2002C";
        ram_buffer(56733) := X"8FB10028";
        ram_buffer(56734) := X"8FB00024";
        ram_buffer(56735) := X"27BD0040";
        ram_buffer(56736) := X"03E00008";
        ram_buffer(56737) := X"00000000";
        ram_buffer(56738) := X"27BDFE78";
        ram_buffer(56739) := X"AFBF0184";
        ram_buffer(56740) := X"AFBE0180";
        ram_buffer(56741) := X"AFB7017C";
        ram_buffer(56742) := X"AFB60178";
        ram_buffer(56743) := X"AFB50174";
        ram_buffer(56744) := X"AFB40170";
        ram_buffer(56745) := X"AFB3016C";
        ram_buffer(56746) := X"AFB20168";
        ram_buffer(56747) := X"AFB10164";
        ram_buffer(56748) := X"AFB00160";
        ram_buffer(56749) := X"03A0F021";
        ram_buffer(56750) := X"AFC40188";
        ram_buffer(56751) := X"AFC5018C";
        ram_buffer(56752) := X"AFC60190";
        ram_buffer(56753) := X"AFC70194";
        ram_buffer(56754) := X"AFC0001C";
        ram_buffer(56755) := X"AFC00020";
        ram_buffer(56756) := X"AFC00024";
        ram_buffer(56757) := X"AFC00028";
        ram_buffer(56758) := X"AFC00048";
        ram_buffer(56759) := X"AFC0004C";
        ram_buffer(56760) := X"8FC2018C";
        ram_buffer(56761) := X"00000000";
        ram_buffer(56762) := X"8442000C";
        ram_buffer(56763) := X"00000000";
        ram_buffer(56764) := X"3042FFFF";
        ram_buffer(56765) := X"30420080";
        ram_buffer(56766) := X"10400024";
        ram_buffer(56767) := X"00000000";
        ram_buffer(56768) := X"8FC2018C";
        ram_buffer(56769) := X"00000000";
        ram_buffer(56770) := X"8C420010";
        ram_buffer(56771) := X"00000000";
        ram_buffer(56772) := X"1440001E";
        ram_buffer(56773) := X"00000000";
        ram_buffer(56774) := X"24050040";
        ram_buffer(56775) := X"8FC40188";
        ram_buffer(56776) := X"0C027B8F";
        ram_buffer(56777) := X"00000000";
        ram_buffer(56778) := X"00401821";
        ram_buffer(56779) := X"8FC2018C";
        ram_buffer(56780) := X"00000000";
        ram_buffer(56781) := X"AC430000";
        ram_buffer(56782) := X"8FC2018C";
        ram_buffer(56783) := X"00000000";
        ram_buffer(56784) := X"8C430000";
        ram_buffer(56785) := X"8FC2018C";
        ram_buffer(56786) := X"00000000";
        ram_buffer(56787) := X"AC430010";
        ram_buffer(56788) := X"8FC2018C";
        ram_buffer(56789) := X"00000000";
        ram_buffer(56790) := X"8C420000";
        ram_buffer(56791) := X"00000000";
        ram_buffer(56792) := X"14400007";
        ram_buffer(56793) := X"00000000";
        ram_buffer(56794) := X"8FC20188";
        ram_buffer(56795) := X"2403000C";
        ram_buffer(56796) := X"AC430000";
        ram_buffer(56797) := X"2402FFFF";
        ram_buffer(56798) := X"10000615";
        ram_buffer(56799) := X"00000000";
        ram_buffer(56800) := X"8FC2018C";
        ram_buffer(56801) := X"24030040";
        ram_buffer(56802) := X"AC430014";
        ram_buffer(56803) := X"8FD50190";
        ram_buffer(56804) := X"27D10068";
        ram_buffer(56805) := X"AFD1005C";
        ram_buffer(56806) := X"AFC00064";
        ram_buffer(56807) := X"AFC00060";
        ram_buffer(56808) := X"AFC00010";
        ram_buffer(56809) := X"02A09821";
        ram_buffer(56810) := X"10000002";
        ram_buffer(56811) := X"00000000";
        ram_buffer(56812) := X"26B50001";
        ram_buffer(56813) := X"82A20000";
        ram_buffer(56814) := X"00000000";
        ram_buffer(56815) := X"10400005";
        ram_buffer(56816) := X"00000000";
        ram_buffer(56817) := X"82A30000";
        ram_buffer(56818) := X"24020025";
        ram_buffer(56819) := X"1462FFF8";
        ram_buffer(56820) := X"00000000";
        ram_buffer(56821) := X"02A01821";
        ram_buffer(56822) := X"02601021";
        ram_buffer(56823) := X"00628023";
        ram_buffer(56824) := X"1200001F";
        ram_buffer(56825) := X"00000000";
        ram_buffer(56826) := X"AE330000";
        ram_buffer(56827) := X"02001021";
        ram_buffer(56828) := X"AE220004";
        ram_buffer(56829) := X"8FC20064";
        ram_buffer(56830) := X"02001821";
        ram_buffer(56831) := X"00431021";
        ram_buffer(56832) := X"AFC20064";
        ram_buffer(56833) := X"26310008";
        ram_buffer(56834) := X"8FC20060";
        ram_buffer(56835) := X"00000000";
        ram_buffer(56836) := X"24420001";
        ram_buffer(56837) := X"AFC20060";
        ram_buffer(56838) := X"8FC20060";
        ram_buffer(56839) := X"00000000";
        ram_buffer(56840) := X"28420008";
        ram_buffer(56841) := X"1440000A";
        ram_buffer(56842) := X"00000000";
        ram_buffer(56843) := X"27C2005C";
        ram_buffer(56844) := X"00403021";
        ram_buffer(56845) := X"8FC5018C";
        ram_buffer(56846) := X"8FC40188";
        ram_buffer(56847) := X"0C02DCA6";
        ram_buffer(56848) := X"00000000";
        ram_buffer(56849) := X"144005A5";
        ram_buffer(56850) := X"00000000";
        ram_buffer(56851) := X"27D10068";
        ram_buffer(56852) := X"8FC20010";
        ram_buffer(56853) := X"00000000";
        ram_buffer(56854) := X"00501021";
        ram_buffer(56855) := X"AFC20010";
        ram_buffer(56856) := X"82A20000";
        ram_buffer(56857) := X"00000000";
        ram_buffer(56858) := X"10400588";
        ram_buffer(56859) := X"00000000";
        ram_buffer(56860) := X"AFD50050";
        ram_buffer(56861) := X"26B50001";
        ram_buffer(56862) := X"00009021";
        ram_buffer(56863) := X"AFC0003C";
        ram_buffer(56864) := X"AFC00014";
        ram_buffer(56865) := X"2402FFFF";
        ram_buffer(56866) := X"AFC20018";
        ram_buffer(56867) := X"A3C00058";
        ram_buffer(56868) := X"02A01021";
        ram_buffer(56869) := X"24550001";
        ram_buffer(56870) := X"80420000";
        ram_buffer(56871) := X"00000000";
        ram_buffer(56872) := X"0040A021";
        ram_buffer(56873) := X"2683FFE0";
        ram_buffer(56874) := X"2C62005B";
        ram_buffer(56875) := X"104003BF";
        ram_buffer(56876) := X"00000000";
        ram_buffer(56877) := X"00031880";
        ram_buffer(56878) := X"3C02100D";
        ram_buffer(56879) := X"2442ABE4";
        ram_buffer(56880) := X"00621021";
        ram_buffer(56881) := X"8C420000";
        ram_buffer(56882) := X"00000000";
        ram_buffer(56883) := X"00400008";
        ram_buffer(56884) := X"00000000";
        ram_buffer(56885) := X"8FC40188";
        ram_buffer(56886) := X"0C02BB25";
        ram_buffer(56887) := X"00000000";
        ram_buffer(56888) := X"8C420004";
        ram_buffer(56889) := X"00000000";
        ram_buffer(56890) := X"AFC2001C";
        ram_buffer(56891) := X"8FC4001C";
        ram_buffer(56892) := X"0C02851E";
        ram_buffer(56893) := X"00000000";
        ram_buffer(56894) := X"AFC20020";
        ram_buffer(56895) := X"8FC40188";
        ram_buffer(56896) := X"0C02BB25";
        ram_buffer(56897) := X"00000000";
        ram_buffer(56898) := X"8C420008";
        ram_buffer(56899) := X"00000000";
        ram_buffer(56900) := X"AFC20024";
        ram_buffer(56901) := X"8FC20020";
        ram_buffer(56902) := X"00000000";
        ram_buffer(56903) := X"1040FFDC";
        ram_buffer(56904) := X"00000000";
        ram_buffer(56905) := X"8FC20024";
        ram_buffer(56906) := X"00000000";
        ram_buffer(56907) := X"1040FFD8";
        ram_buffer(56908) := X"00000000";
        ram_buffer(56909) := X"8FC20024";
        ram_buffer(56910) := X"00000000";
        ram_buffer(56911) := X"80420000";
        ram_buffer(56912) := X"00000000";
        ram_buffer(56913) := X"1040FFD2";
        ram_buffer(56914) := X"00000000";
        ram_buffer(56915) := X"36520400";
        ram_buffer(56916) := X"1000FFCF";
        ram_buffer(56917) := X"00000000";
        ram_buffer(56918) := X"83C20058";
        ram_buffer(56919) := X"00000000";
        ram_buffer(56920) := X"1440FFCB";
        ram_buffer(56921) := X"00000000";
        ram_buffer(56922) := X"24020020";
        ram_buffer(56923) := X"A3C20058";
        ram_buffer(56924) := X"1000FFC7";
        ram_buffer(56925) := X"00000000";
        ram_buffer(56926) := X"36520001";
        ram_buffer(56927) := X"1000FFC4";
        ram_buffer(56928) := X"00000000";
        ram_buffer(56929) := X"8FC20194";
        ram_buffer(56930) := X"00000000";
        ram_buffer(56931) := X"24430004";
        ram_buffer(56932) := X"AFC30194";
        ram_buffer(56933) := X"8C420000";
        ram_buffer(56934) := X"00000000";
        ram_buffer(56935) := X"AFC20014";
        ram_buffer(56936) := X"8FC20014";
        ram_buffer(56937) := X"00000000";
        ram_buffer(56938) := X"04400003";
        ram_buffer(56939) := X"00000000";
        ram_buffer(56940) := X"1000FFB7";
        ram_buffer(56941) := X"00000000";
        ram_buffer(56942) := X"8FC20014";
        ram_buffer(56943) := X"00000000";
        ram_buffer(56944) := X"00021023";
        ram_buffer(56945) := X"AFC20014";
        ram_buffer(56946) := X"36520004";
        ram_buffer(56947) := X"1000FFB0";
        ram_buffer(56948) := X"00000000";
        ram_buffer(56949) := X"2402002B";
        ram_buffer(56950) := X"A3C20058";
        ram_buffer(56951) := X"1000FFAC";
        ram_buffer(56952) := X"00000000";
        ram_buffer(56953) := X"02A01021";
        ram_buffer(56954) := X"24550001";
        ram_buffer(56955) := X"80420000";
        ram_buffer(56956) := X"00000000";
        ram_buffer(56957) := X"0040A021";
        ram_buffer(56958) := X"2402002A";
        ram_buffer(56959) := X"16820010";
        ram_buffer(56960) := X"00000000";
        ram_buffer(56961) := X"8FC20194";
        ram_buffer(56962) := X"00000000";
        ram_buffer(56963) := X"24430004";
        ram_buffer(56964) := X"AFC30194";
        ram_buffer(56965) := X"8C420000";
        ram_buffer(56966) := X"00000000";
        ram_buffer(56967) := X"AFC20018";
        ram_buffer(56968) := X"8FC20018";
        ram_buffer(56969) := X"00000000";
        ram_buffer(56970) := X"0441FF99";
        ram_buffer(56971) := X"00000000";
        ram_buffer(56972) := X"2402FFFF";
        ram_buffer(56973) := X"AFC20018";
        ram_buffer(56974) := X"1000FF95";
        ram_buffer(56975) := X"00000000";
        ram_buffer(56976) := X"00008021";
        ram_buffer(56977) := X"1000000D";
        ram_buffer(56978) := X"00000000";
        ram_buffer(56979) := X"02001821";
        ram_buffer(56980) := X"00031040";
        ram_buffer(56981) := X"00401821";
        ram_buffer(56982) := X"00031080";
        ram_buffer(56983) := X"00621821";
        ram_buffer(56984) := X"2682FFD0";
        ram_buffer(56985) := X"00628021";
        ram_buffer(56986) := X"02A01021";
        ram_buffer(56987) := X"24550001";
        ram_buffer(56988) := X"80420000";
        ram_buffer(56989) := X"00000000";
        ram_buffer(56990) := X"0040A021";
        ram_buffer(56991) := X"2682FFD0";
        ram_buffer(56992) := X"2C42000A";
        ram_buffer(56993) := X"1440FFF1";
        ram_buffer(56994) := X"00000000";
        ram_buffer(56995) := X"02001021";
        ram_buffer(56996) := X"04410002";
        ram_buffer(56997) := X"00000000";
        ram_buffer(56998) := X"2402FFFF";
        ram_buffer(56999) := X"AFC20018";
        ram_buffer(57000) := X"1000FF80";
        ram_buffer(57001) := X"00000000";
        ram_buffer(57002) := X"36520080";
        ram_buffer(57003) := X"1000FF78";
        ram_buffer(57004) := X"00000000";
        ram_buffer(57005) := X"00008021";
        ram_buffer(57006) := X"02001821";
        ram_buffer(57007) := X"00031040";
        ram_buffer(57008) := X"00401821";
        ram_buffer(57009) := X"00031080";
        ram_buffer(57010) := X"00621821";
        ram_buffer(57011) := X"2682FFD0";
        ram_buffer(57012) := X"00628021";
        ram_buffer(57013) := X"02A01021";
        ram_buffer(57014) := X"24550001";
        ram_buffer(57015) := X"80420000";
        ram_buffer(57016) := X"00000000";
        ram_buffer(57017) := X"0040A021";
        ram_buffer(57018) := X"2682FFD0";
        ram_buffer(57019) := X"2C42000A";
        ram_buffer(57020) := X"1440FFF1";
        ram_buffer(57021) := X"00000000";
        ram_buffer(57022) := X"AFD00014";
        ram_buffer(57023) := X"1000FF69";
        ram_buffer(57024) := X"00000000";
        ram_buffer(57025) := X"82A30000";
        ram_buffer(57026) := X"24020068";
        ram_buffer(57027) := X"14620005";
        ram_buffer(57028) := X"00000000";
        ram_buffer(57029) := X"26B50001";
        ram_buffer(57030) := X"36520200";
        ram_buffer(57031) := X"1000FF5C";
        ram_buffer(57032) := X"00000000";
        ram_buffer(57033) := X"36520040";
        ram_buffer(57034) := X"1000FF59";
        ram_buffer(57035) := X"00000000";
        ram_buffer(57036) := X"82A30000";
        ram_buffer(57037) := X"2402006C";
        ram_buffer(57038) := X"14620005";
        ram_buffer(57039) := X"00000000";
        ram_buffer(57040) := X"26B50001";
        ram_buffer(57041) := X"36520020";
        ram_buffer(57042) := X"1000FF51";
        ram_buffer(57043) := X"00000000";
        ram_buffer(57044) := X"36520010";
        ram_buffer(57045) := X"1000FF4E";
        ram_buffer(57046) := X"00000000";
        ram_buffer(57047) := X"36520020";
        ram_buffer(57048) := X"1000FF4B";
        ram_buffer(57049) := X"00000000";
        ram_buffer(57050) := X"36520020";
        ram_buffer(57051) := X"1000FF48";
        ram_buffer(57052) := X"00000000";
        ram_buffer(57053) := X"27D300A8";
        ram_buffer(57054) := X"8FC30194";
        ram_buffer(57055) := X"00000000";
        ram_buffer(57056) := X"24620004";
        ram_buffer(57057) := X"AFC20194";
        ram_buffer(57058) := X"8C620000";
        ram_buffer(57059) := X"00000000";
        ram_buffer(57060) := X"00021600";
        ram_buffer(57061) := X"00021603";
        ram_buffer(57062) := X"A2620000";
        ram_buffer(57063) := X"24020001";
        ram_buffer(57064) := X"AFC20044";
        ram_buffer(57065) := X"A3C00058";
        ram_buffer(57066) := X"1000030A";
        ram_buffer(57067) := X"00000000";
        ram_buffer(57068) := X"36520010";
        ram_buffer(57069) := X"32420020";
        ram_buffer(57070) := X"1040000E";
        ram_buffer(57071) := X"00000000";
        ram_buffer(57072) := X"8FC20194";
        ram_buffer(57073) := X"00000000";
        ram_buffer(57074) := X"24430007";
        ram_buffer(57075) := X"2402FFF8";
        ram_buffer(57076) := X"00621024";
        ram_buffer(57077) := X"24430008";
        ram_buffer(57078) := X"AFC30194";
        ram_buffer(57079) := X"8C430004";
        ram_buffer(57080) := X"8C420000";
        ram_buffer(57081) := X"AFC30114";
        ram_buffer(57082) := X"AFC20110";
        ram_buffer(57083) := X"10000038";
        ram_buffer(57084) := X"00000000";
        ram_buffer(57085) := X"32420010";
        ram_buffer(57086) := X"1040000C";
        ram_buffer(57087) := X"00000000";
        ram_buffer(57088) := X"8FC20194";
        ram_buffer(57089) := X"00000000";
        ram_buffer(57090) := X"24430004";
        ram_buffer(57091) := X"AFC30194";
        ram_buffer(57092) := X"8C420000";
        ram_buffer(57093) := X"00000000";
        ram_buffer(57094) := X"AFC20114";
        ram_buffer(57095) := X"000217C3";
        ram_buffer(57096) := X"AFC20110";
        ram_buffer(57097) := X"1000002A";
        ram_buffer(57098) := X"00000000";
        ram_buffer(57099) := X"32420040";
        ram_buffer(57100) := X"1040000E";
        ram_buffer(57101) := X"00000000";
        ram_buffer(57102) := X"8FC20194";
        ram_buffer(57103) := X"00000000";
        ram_buffer(57104) := X"24430004";
        ram_buffer(57105) := X"AFC30194";
        ram_buffer(57106) := X"8C420000";
        ram_buffer(57107) := X"00000000";
        ram_buffer(57108) := X"00021400";
        ram_buffer(57109) := X"00021403";
        ram_buffer(57110) := X"AFC20114";
        ram_buffer(57111) := X"000217C3";
        ram_buffer(57112) := X"AFC20110";
        ram_buffer(57113) := X"1000001A";
        ram_buffer(57114) := X"00000000";
        ram_buffer(57115) := X"32420200";
        ram_buffer(57116) := X"1040000E";
        ram_buffer(57117) := X"00000000";
        ram_buffer(57118) := X"8FC20194";
        ram_buffer(57119) := X"00000000";
        ram_buffer(57120) := X"24430004";
        ram_buffer(57121) := X"AFC30194";
        ram_buffer(57122) := X"8C420000";
        ram_buffer(57123) := X"00000000";
        ram_buffer(57124) := X"00021600";
        ram_buffer(57125) := X"00021603";
        ram_buffer(57126) := X"AFC20114";
        ram_buffer(57127) := X"000217C3";
        ram_buffer(57128) := X"AFC20110";
        ram_buffer(57129) := X"1000000A";
        ram_buffer(57130) := X"00000000";
        ram_buffer(57131) := X"8FC20194";
        ram_buffer(57132) := X"00000000";
        ram_buffer(57133) := X"24430004";
        ram_buffer(57134) := X"AFC30194";
        ram_buffer(57135) := X"8C420000";
        ram_buffer(57136) := X"00000000";
        ram_buffer(57137) := X"AFC20114";
        ram_buffer(57138) := X"000217C3";
        ram_buffer(57139) := X"AFC20110";
        ram_buffer(57140) := X"8FC30114";
        ram_buffer(57141) := X"8FC20110";
        ram_buffer(57142) := X"AFC30034";
        ram_buffer(57143) := X"AFC20030";
        ram_buffer(57144) := X"8FC30034";
        ram_buffer(57145) := X"8FC20030";
        ram_buffer(57146) := X"00000000";
        ram_buffer(57147) := X"0441000E";
        ram_buffer(57148) := X"00000000";
        ram_buffer(57149) := X"00001821";
        ram_buffer(57150) := X"00001021";
        ram_buffer(57151) := X"8FC50034";
        ram_buffer(57152) := X"8FC40030";
        ram_buffer(57153) := X"00653823";
        ram_buffer(57154) := X"0067402B";
        ram_buffer(57155) := X"00443023";
        ram_buffer(57156) := X"00C81023";
        ram_buffer(57157) := X"00403021";
        ram_buffer(57158) := X"AFC70034";
        ram_buffer(57159) := X"AFC60030";
        ram_buffer(57160) := X"2402002D";
        ram_buffer(57161) := X"A3C20058";
        ram_buffer(57162) := X"24020001";
        ram_buffer(57163) := X"A3C20038";
        ram_buffer(57164) := X"100001AB";
        ram_buffer(57165) := X"00000000";
        ram_buffer(57166) := X"32420020";
        ram_buffer(57167) := X"10400011";
        ram_buffer(57168) := X"00000000";
        ram_buffer(57169) := X"8FC20194";
        ram_buffer(57170) := X"00000000";
        ram_buffer(57171) := X"24430004";
        ram_buffer(57172) := X"AFC30194";
        ram_buffer(57173) := X"8C430000";
        ram_buffer(57174) := X"8FC20010";
        ram_buffer(57175) := X"00000000";
        ram_buffer(57176) := X"AFC2012C";
        ram_buffer(57177) := X"000217C3";
        ram_buffer(57178) := X"AFC20128";
        ram_buffer(57179) := X"8FC5012C";
        ram_buffer(57180) := X"8FC40128";
        ram_buffer(57181) := X"AC650004";
        ram_buffer(57182) := X"AC640000";
        ram_buffer(57183) := X"10000441";
        ram_buffer(57184) := X"00000000";
        ram_buffer(57185) := X"32420010";
        ram_buffer(57186) := X"1040000B";
        ram_buffer(57187) := X"00000000";
        ram_buffer(57188) := X"8FC20194";
        ram_buffer(57189) := X"00000000";
        ram_buffer(57190) := X"24430004";
        ram_buffer(57191) := X"AFC30194";
        ram_buffer(57192) := X"8C420000";
        ram_buffer(57193) := X"8FC30010";
        ram_buffer(57194) := X"00000000";
        ram_buffer(57195) := X"AC430000";
        ram_buffer(57196) := X"10000434";
        ram_buffer(57197) := X"00000000";
        ram_buffer(57198) := X"32420040";
        ram_buffer(57199) := X"1040000D";
        ram_buffer(57200) := X"00000000";
        ram_buffer(57201) := X"8FC20194";
        ram_buffer(57202) := X"00000000";
        ram_buffer(57203) := X"24430004";
        ram_buffer(57204) := X"AFC30194";
        ram_buffer(57205) := X"8C420000";
        ram_buffer(57206) := X"8FC30010";
        ram_buffer(57207) := X"00000000";
        ram_buffer(57208) := X"00031C00";
        ram_buffer(57209) := X"00031C03";
        ram_buffer(57210) := X"A4430000";
        ram_buffer(57211) := X"10000425";
        ram_buffer(57212) := X"00000000";
        ram_buffer(57213) := X"32420200";
        ram_buffer(57214) := X"1040000D";
        ram_buffer(57215) := X"00000000";
        ram_buffer(57216) := X"8FC20194";
        ram_buffer(57217) := X"00000000";
        ram_buffer(57218) := X"24430004";
        ram_buffer(57219) := X"AFC30194";
        ram_buffer(57220) := X"8C420000";
        ram_buffer(57221) := X"8FC30010";
        ram_buffer(57222) := X"00000000";
        ram_buffer(57223) := X"00031E00";
        ram_buffer(57224) := X"00031E03";
        ram_buffer(57225) := X"A0430000";
        ram_buffer(57226) := X"10000416";
        ram_buffer(57227) := X"00000000";
        ram_buffer(57228) := X"8FC20194";
        ram_buffer(57229) := X"00000000";
        ram_buffer(57230) := X"24430004";
        ram_buffer(57231) := X"AFC30194";
        ram_buffer(57232) := X"8C420000";
        ram_buffer(57233) := X"8FC30010";
        ram_buffer(57234) := X"00000000";
        ram_buffer(57235) := X"AC430000";
        ram_buffer(57236) := X"1000040C";
        ram_buffer(57237) := X"00000000";
        ram_buffer(57238) := X"36520010";
        ram_buffer(57239) := X"32420020";
        ram_buffer(57240) := X"1040000C";
        ram_buffer(57241) := X"00000000";
        ram_buffer(57242) := X"8FC20194";
        ram_buffer(57243) := X"00000000";
        ram_buffer(57244) := X"24430007";
        ram_buffer(57245) := X"2402FFF8";
        ram_buffer(57246) := X"00621024";
        ram_buffer(57247) := X"24430008";
        ram_buffer(57248) := X"AFC30194";
        ram_buffer(57249) := X"8C570004";
        ram_buffer(57250) := X"8C560000";
        ram_buffer(57251) := X"1000003C";
        ram_buffer(57252) := X"00000000";
        ram_buffer(57253) := X"32420010";
        ram_buffer(57254) := X"1040000B";
        ram_buffer(57255) := X"00000000";
        ram_buffer(57256) := X"8FC20194";
        ram_buffer(57257) := X"00000000";
        ram_buffer(57258) := X"24430004";
        ram_buffer(57259) := X"AFC30194";
        ram_buffer(57260) := X"8C420000";
        ram_buffer(57261) := X"00000000";
        ram_buffer(57262) := X"0040B821";
        ram_buffer(57263) := X"0000B021";
        ram_buffer(57264) := X"1000002F";
        ram_buffer(57265) := X"00000000";
        ram_buffer(57266) := X"32420040";
        ram_buffer(57267) := X"10400011";
        ram_buffer(57268) := X"00000000";
        ram_buffer(57269) := X"8FC20194";
        ram_buffer(57270) := X"00000000";
        ram_buffer(57271) := X"24430004";
        ram_buffer(57272) := X"AFC30194";
        ram_buffer(57273) := X"8C420000";
        ram_buffer(57274) := X"00000000";
        ram_buffer(57275) := X"AFC20134";
        ram_buffer(57276) := X"AFC00130";
        ram_buffer(57277) := X"8FC30134";
        ram_buffer(57278) := X"8FC20130";
        ram_buffer(57279) := X"00000000";
        ram_buffer(57280) := X"00402021";
        ram_buffer(57281) := X"30960000";
        ram_buffer(57282) := X"3077FFFF";
        ram_buffer(57283) := X"1000001C";
        ram_buffer(57284) := X"00000000";
        ram_buffer(57285) := X"32420200";
        ram_buffer(57286) := X"10400011";
        ram_buffer(57287) := X"00000000";
        ram_buffer(57288) := X"8FC20194";
        ram_buffer(57289) := X"00000000";
        ram_buffer(57290) := X"24430004";
        ram_buffer(57291) := X"AFC30194";
        ram_buffer(57292) := X"8C420000";
        ram_buffer(57293) := X"00000000";
        ram_buffer(57294) := X"AFC2013C";
        ram_buffer(57295) := X"AFC00138";
        ram_buffer(57296) := X"8FC3013C";
        ram_buffer(57297) := X"8FC20138";
        ram_buffer(57298) := X"00000000";
        ram_buffer(57299) := X"00402021";
        ram_buffer(57300) := X"30960000";
        ram_buffer(57301) := X"307700FF";
        ram_buffer(57302) := X"10000009";
        ram_buffer(57303) := X"00000000";
        ram_buffer(57304) := X"8FC20194";
        ram_buffer(57305) := X"00000000";
        ram_buffer(57306) := X"24430004";
        ram_buffer(57307) := X"AFC30194";
        ram_buffer(57308) := X"8C420000";
        ram_buffer(57309) := X"00000000";
        ram_buffer(57310) := X"0040B821";
        ram_buffer(57311) := X"0000B021";
        ram_buffer(57312) := X"AFD70034";
        ram_buffer(57313) := X"AFD60030";
        ram_buffer(57314) := X"A3C00038";
        ram_buffer(57315) := X"2402FBFF";
        ram_buffer(57316) := X"02429024";
        ram_buffer(57317) := X"10000111";
        ram_buffer(57318) := X"00000000";
        ram_buffer(57319) := X"8FC20194";
        ram_buffer(57320) := X"00000000";
        ram_buffer(57321) := X"24430004";
        ram_buffer(57322) := X"AFC30194";
        ram_buffer(57323) := X"8C420000";
        ram_buffer(57324) := X"00000000";
        ram_buffer(57325) := X"AFC20034";
        ram_buffer(57326) := X"AFC00030";
        ram_buffer(57327) := X"24020002";
        ram_buffer(57328) := X"A3C20038";
        ram_buffer(57329) := X"3C02100D";
        ram_buffer(57330) := X"2442AB98";
        ram_buffer(57331) := X"AFC20048";
        ram_buffer(57332) := X"36520002";
        ram_buffer(57333) := X"24020030";
        ram_buffer(57334) := X"A3C2010C";
        ram_buffer(57335) := X"24140078";
        ram_buffer(57336) := X"24020078";
        ram_buffer(57337) := X"A3C2010D";
        ram_buffer(57338) := X"100000FC";
        ram_buffer(57339) := X"00000000";
        ram_buffer(57340) := X"8FC20194";
        ram_buffer(57341) := X"00000000";
        ram_buffer(57342) := X"24430004";
        ram_buffer(57343) := X"AFC30194";
        ram_buffer(57344) := X"8C530000";
        ram_buffer(57345) := X"A3C00058";
        ram_buffer(57346) := X"1660000D";
        ram_buffer(57347) := X"00000000";
        ram_buffer(57348) := X"3C02100D";
        ram_buffer(57349) := X"2453ABAC";
        ram_buffer(57350) := X"8FC20018";
        ram_buffer(57351) := X"00000000";
        ram_buffer(57352) := X"00401821";
        ram_buffer(57353) := X"2C620007";
        ram_buffer(57354) := X"14400002";
        ram_buffer(57355) := X"00000000";
        ram_buffer(57356) := X"24030006";
        ram_buffer(57357) := X"AFC30044";
        ram_buffer(57358) := X"100001E6";
        ram_buffer(57359) := X"00000000";
        ram_buffer(57360) := X"8FC20018";
        ram_buffer(57361) := X"00000000";
        ram_buffer(57362) := X"04400018";
        ram_buffer(57363) := X"00000000";
        ram_buffer(57364) := X"8FC20018";
        ram_buffer(57365) := X"00000000";
        ram_buffer(57366) := X"00403021";
        ram_buffer(57367) := X"00002821";
        ram_buffer(57368) := X"02602021";
        ram_buffer(57369) := X"0C02BC51";
        ram_buffer(57370) := X"00000000";
        ram_buffer(57371) := X"AFC20054";
        ram_buffer(57372) := X"8FC20054";
        ram_buffer(57373) := X"00000000";
        ram_buffer(57374) := X"10400007";
        ram_buffer(57375) := X"00000000";
        ram_buffer(57376) := X"8FC30054";
        ram_buffer(57377) := X"02601021";
        ram_buffer(57378) := X"00621023";
        ram_buffer(57379) := X"AFC20044";
        ram_buffer(57380) := X"100001D0";
        ram_buffer(57381) := X"00000000";
        ram_buffer(57382) := X"8FC20018";
        ram_buffer(57383) := X"00000000";
        ram_buffer(57384) := X"AFC20044";
        ram_buffer(57385) := X"100001CB";
        ram_buffer(57386) := X"00000000";
        ram_buffer(57387) := X"02602021";
        ram_buffer(57388) := X"0C02851E";
        ram_buffer(57389) := X"00000000";
        ram_buffer(57390) := X"AFC20044";
        ram_buffer(57391) := X"100001C5";
        ram_buffer(57392) := X"00000000";
        ram_buffer(57393) := X"36520010";
        ram_buffer(57394) := X"32420020";
        ram_buffer(57395) := X"1040000E";
        ram_buffer(57396) := X"00000000";
        ram_buffer(57397) := X"8FC20194";
        ram_buffer(57398) := X"00000000";
        ram_buffer(57399) := X"24430007";
        ram_buffer(57400) := X"2402FFF8";
        ram_buffer(57401) := X"00621024";
        ram_buffer(57402) := X"24430008";
        ram_buffer(57403) := X"AFC30194";
        ram_buffer(57404) := X"8C430004";
        ram_buffer(57405) := X"8C420000";
        ram_buffer(57406) := X"AFC3011C";
        ram_buffer(57407) := X"AFC20118";
        ram_buffer(57408) := X"10000040";
        ram_buffer(57409) := X"00000000";
        ram_buffer(57410) := X"32420010";
        ram_buffer(57411) := X"1040000B";
        ram_buffer(57412) := X"00000000";
        ram_buffer(57413) := X"8FC20194";
        ram_buffer(57414) := X"00000000";
        ram_buffer(57415) := X"24430004";
        ram_buffer(57416) := X"AFC30194";
        ram_buffer(57417) := X"8C420000";
        ram_buffer(57418) := X"00000000";
        ram_buffer(57419) := X"AFC2011C";
        ram_buffer(57420) := X"AFC00118";
        ram_buffer(57421) := X"10000033";
        ram_buffer(57422) := X"00000000";
        ram_buffer(57423) := X"32420040";
        ram_buffer(57424) := X"10400013";
        ram_buffer(57425) := X"00000000";
        ram_buffer(57426) := X"8FC20194";
        ram_buffer(57427) := X"00000000";
        ram_buffer(57428) := X"24430004";
        ram_buffer(57429) := X"AFC30194";
        ram_buffer(57430) := X"8C420000";
        ram_buffer(57431) := X"00000000";
        ram_buffer(57432) := X"AFC20144";
        ram_buffer(57433) := X"AFC00140";
        ram_buffer(57434) := X"8FC30144";
        ram_buffer(57435) := X"8FC20140";
        ram_buffer(57436) := X"00000000";
        ram_buffer(57437) := X"00402021";
        ram_buffer(57438) := X"30840000";
        ram_buffer(57439) := X"AFC40118";
        ram_buffer(57440) := X"3062FFFF";
        ram_buffer(57441) := X"AFC2011C";
        ram_buffer(57442) := X"1000001E";
        ram_buffer(57443) := X"00000000";
        ram_buffer(57444) := X"32420200";
        ram_buffer(57445) := X"10400013";
        ram_buffer(57446) := X"00000000";
        ram_buffer(57447) := X"8FC20194";
        ram_buffer(57448) := X"00000000";
        ram_buffer(57449) := X"24430004";
        ram_buffer(57450) := X"AFC30194";
        ram_buffer(57451) := X"8C420000";
        ram_buffer(57452) := X"00000000";
        ram_buffer(57453) := X"AFC2014C";
        ram_buffer(57454) := X"AFC00148";
        ram_buffer(57455) := X"8FC3014C";
        ram_buffer(57456) := X"8FC20148";
        ram_buffer(57457) := X"00000000";
        ram_buffer(57458) := X"00402021";
        ram_buffer(57459) := X"30840000";
        ram_buffer(57460) := X"AFC40118";
        ram_buffer(57461) := X"306200FF";
        ram_buffer(57462) := X"AFC2011C";
        ram_buffer(57463) := X"10000009";
        ram_buffer(57464) := X"00000000";
        ram_buffer(57465) := X"8FC20194";
        ram_buffer(57466) := X"00000000";
        ram_buffer(57467) := X"24430004";
        ram_buffer(57468) := X"AFC30194";
        ram_buffer(57469) := X"8C420000";
        ram_buffer(57470) := X"00000000";
        ram_buffer(57471) := X"AFC2011C";
        ram_buffer(57472) := X"AFC00118";
        ram_buffer(57473) := X"8FC3011C";
        ram_buffer(57474) := X"8FC20118";
        ram_buffer(57475) := X"AFC30034";
        ram_buffer(57476) := X"AFC20030";
        ram_buffer(57477) := X"24020001";
        ram_buffer(57478) := X"A3C20038";
        ram_buffer(57479) := X"1000006F";
        ram_buffer(57480) := X"00000000";
        ram_buffer(57481) := X"3C02100D";
        ram_buffer(57482) := X"2442ABB4";
        ram_buffer(57483) := X"AFC20048";
        ram_buffer(57484) := X"10000004";
        ram_buffer(57485) := X"00000000";
        ram_buffer(57486) := X"3C02100D";
        ram_buffer(57487) := X"2442AB98";
        ram_buffer(57488) := X"AFC20048";
        ram_buffer(57489) := X"32420020";
        ram_buffer(57490) := X"1040000E";
        ram_buffer(57491) := X"00000000";
        ram_buffer(57492) := X"8FC20194";
        ram_buffer(57493) := X"00000000";
        ram_buffer(57494) := X"24430007";
        ram_buffer(57495) := X"2402FFF8";
        ram_buffer(57496) := X"00621024";
        ram_buffer(57497) := X"24430008";
        ram_buffer(57498) := X"AFC30194";
        ram_buffer(57499) := X"8C430004";
        ram_buffer(57500) := X"8C420000";
        ram_buffer(57501) := X"AFC30124";
        ram_buffer(57502) := X"AFC20120";
        ram_buffer(57503) := X"10000040";
        ram_buffer(57504) := X"00000000";
        ram_buffer(57505) := X"32420010";
        ram_buffer(57506) := X"1040000B";
        ram_buffer(57507) := X"00000000";
        ram_buffer(57508) := X"8FC30194";
        ram_buffer(57509) := X"00000000";
        ram_buffer(57510) := X"24620004";
        ram_buffer(57511) := X"AFC20194";
        ram_buffer(57512) := X"8C620000";
        ram_buffer(57513) := X"00000000";
        ram_buffer(57514) := X"AFC20124";
        ram_buffer(57515) := X"AFC00120";
        ram_buffer(57516) := X"10000033";
        ram_buffer(57517) := X"00000000";
        ram_buffer(57518) := X"32420040";
        ram_buffer(57519) := X"10400013";
        ram_buffer(57520) := X"00000000";
        ram_buffer(57521) := X"8FC30194";
        ram_buffer(57522) := X"00000000";
        ram_buffer(57523) := X"24620004";
        ram_buffer(57524) := X"AFC20194";
        ram_buffer(57525) := X"8C620000";
        ram_buffer(57526) := X"00000000";
        ram_buffer(57527) := X"AFC20154";
        ram_buffer(57528) := X"AFC00150";
        ram_buffer(57529) := X"8FC30154";
        ram_buffer(57530) := X"8FC20150";
        ram_buffer(57531) := X"00000000";
        ram_buffer(57532) := X"00402021";
        ram_buffer(57533) := X"30840000";
        ram_buffer(57534) := X"AFC40120";
        ram_buffer(57535) := X"3062FFFF";
        ram_buffer(57536) := X"AFC20124";
        ram_buffer(57537) := X"1000001E";
        ram_buffer(57538) := X"00000000";
        ram_buffer(57539) := X"32420200";
        ram_buffer(57540) := X"10400013";
        ram_buffer(57541) := X"00000000";
        ram_buffer(57542) := X"8FC30194";
        ram_buffer(57543) := X"00000000";
        ram_buffer(57544) := X"24620004";
        ram_buffer(57545) := X"AFC20194";
        ram_buffer(57546) := X"8C620000";
        ram_buffer(57547) := X"00000000";
        ram_buffer(57548) := X"AFC2015C";
        ram_buffer(57549) := X"AFC00158";
        ram_buffer(57550) := X"8FC3015C";
        ram_buffer(57551) := X"8FC20158";
        ram_buffer(57552) := X"00000000";
        ram_buffer(57553) := X"00402021";
        ram_buffer(57554) := X"30840000";
        ram_buffer(57555) := X"AFC40120";
        ram_buffer(57556) := X"306200FF";
        ram_buffer(57557) := X"AFC20124";
        ram_buffer(57558) := X"10000009";
        ram_buffer(57559) := X"00000000";
        ram_buffer(57560) := X"8FC30194";
        ram_buffer(57561) := X"00000000";
        ram_buffer(57562) := X"24620004";
        ram_buffer(57563) := X"AFC20194";
        ram_buffer(57564) := X"8C620000";
        ram_buffer(57565) := X"00000000";
        ram_buffer(57566) := X"AFC20124";
        ram_buffer(57567) := X"AFC00120";
        ram_buffer(57568) := X"8FC30124";
        ram_buffer(57569) := X"8FC20120";
        ram_buffer(57570) := X"AFC30034";
        ram_buffer(57571) := X"AFC20030";
        ram_buffer(57572) := X"24020002";
        ram_buffer(57573) := X"A3C20038";
        ram_buffer(57574) := X"32420001";
        ram_buffer(57575) := X"1040000D";
        ram_buffer(57576) := X"00000000";
        ram_buffer(57577) := X"8FC20030";
        ram_buffer(57578) := X"8FC30034";
        ram_buffer(57579) := X"00000000";
        ram_buffer(57580) := X"00431025";
        ram_buffer(57581) := X"10400007";
        ram_buffer(57582) := X"00000000";
        ram_buffer(57583) := X"24020030";
        ram_buffer(57584) := X"A3C2010C";
        ram_buffer(57585) := X"00141600";
        ram_buffer(57586) := X"00021603";
        ram_buffer(57587) := X"A3C2010D";
        ram_buffer(57588) := X"36520002";
        ram_buffer(57589) := X"2402FBFF";
        ram_buffer(57590) := X"02429024";
        ram_buffer(57591) := X"A3C00058";
        ram_buffer(57592) := X"8FC20018";
        ram_buffer(57593) := X"00000000";
        ram_buffer(57594) := X"AFC2003C";
        ram_buffer(57595) := X"8FC2003C";
        ram_buffer(57596) := X"00000000";
        ram_buffer(57597) := X"04400003";
        ram_buffer(57598) := X"00000000";
        ram_buffer(57599) := X"2402FF7F";
        ram_buffer(57600) := X"02429024";
        ram_buffer(57601) := X"27D300A8";
        ram_buffer(57602) := X"26730064";
        ram_buffer(57603) := X"8FC20030";
        ram_buffer(57604) := X"8FC30034";
        ram_buffer(57605) := X"00000000";
        ram_buffer(57606) := X"00431025";
        ram_buffer(57607) := X"14400005";
        ram_buffer(57608) := X"00000000";
        ram_buffer(57609) := X"8FC20018";
        ram_buffer(57610) := X"00000000";
        ram_buffer(57611) := X"104000CD";
        ram_buffer(57612) := X"00000000";
        ram_buffer(57613) := X"93C30038";
        ram_buffer(57614) := X"24020001";
        ram_buffer(57615) := X"1062002E";
        ram_buffer(57616) := X"00000000";
        ram_buffer(57617) := X"24020002";
        ram_buffer(57618) := X"1062009C";
        ram_buffer(57619) := X"00000000";
        ram_buffer(57620) := X"146000B8";
        ram_buffer(57621) := X"00000000";
        ram_buffer(57622) := X"2673FFFF";
        ram_buffer(57623) := X"93C20037";
        ram_buffer(57624) := X"00000000";
        ram_buffer(57625) := X"30420007";
        ram_buffer(57626) := X"304200FF";
        ram_buffer(57627) := X"24420030";
        ram_buffer(57628) := X"304200FF";
        ram_buffer(57629) := X"00021600";
        ram_buffer(57630) := X"00021603";
        ram_buffer(57631) := X"A2620000";
        ram_buffer(57632) := X"8FC20030";
        ram_buffer(57633) := X"00000000";
        ram_buffer(57634) := X"00021F40";
        ram_buffer(57635) := X"8FC20034";
        ram_buffer(57636) := X"00000000";
        ram_buffer(57637) := X"000210C2";
        ram_buffer(57638) := X"00431025";
        ram_buffer(57639) := X"AFC20034";
        ram_buffer(57640) := X"8FC20030";
        ram_buffer(57641) := X"00000000";
        ram_buffer(57642) := X"000210C2";
        ram_buffer(57643) := X"AFC20030";
        ram_buffer(57644) := X"8FC20030";
        ram_buffer(57645) := X"8FC30034";
        ram_buffer(57646) := X"00000000";
        ram_buffer(57647) := X"00431025";
        ram_buffer(57648) := X"1440FFE5";
        ram_buffer(57649) := X"00000000";
        ram_buffer(57650) := X"32420001";
        ram_buffer(57651) := X"104000A2";
        ram_buffer(57652) := X"00000000";
        ram_buffer(57653) := X"82630000";
        ram_buffer(57654) := X"24020030";
        ram_buffer(57655) := X"1062009E";
        ram_buffer(57656) := X"00000000";
        ram_buffer(57657) := X"2673FFFF";
        ram_buffer(57658) := X"24020030";
        ram_buffer(57659) := X"A2620000";
        ram_buffer(57660) := X"10000099";
        ram_buffer(57661) := X"00000000";
        ram_buffer(57662) := X"8FC20030";
        ram_buffer(57663) := X"00000000";
        ram_buffer(57664) := X"14400014";
        ram_buffer(57665) := X"00000000";
        ram_buffer(57666) := X"8FC20030";
        ram_buffer(57667) := X"00000000";
        ram_buffer(57668) := X"14400006";
        ram_buffer(57669) := X"00000000";
        ram_buffer(57670) := X"8FC20034";
        ram_buffer(57671) := X"00000000";
        ram_buffer(57672) := X"2C42000A";
        ram_buffer(57673) := X"1040000B";
        ram_buffer(57674) := X"00000000";
        ram_buffer(57675) := X"2673FFFF";
        ram_buffer(57676) := X"93C20037";
        ram_buffer(57677) := X"00000000";
        ram_buffer(57678) := X"24420030";
        ram_buffer(57679) := X"304200FF";
        ram_buffer(57680) := X"00021600";
        ram_buffer(57681) := X"00021603";
        ram_buffer(57682) := X"A2620000";
        ram_buffer(57683) := X"10000083";
        ram_buffer(57684) := X"00000000";
        ram_buffer(57685) := X"AFC00028";
        ram_buffer(57686) := X"2673FFFF";
        ram_buffer(57687) := X"8FC30034";
        ram_buffer(57688) := X"8FC20030";
        ram_buffer(57689) := X"2407000A";
        ram_buffer(57690) := X"00003021";
        ram_buffer(57691) := X"00602821";
        ram_buffer(57692) := X"00402021";
        ram_buffer(57693) := X"0C030BFE";
        ram_buffer(57694) := X"00000000";
        ram_buffer(57695) := X"306200FF";
        ram_buffer(57696) := X"24420030";
        ram_buffer(57697) := X"304200FF";
        ram_buffer(57698) := X"00021600";
        ram_buffer(57699) := X"00021603";
        ram_buffer(57700) := X"A2620000";
        ram_buffer(57701) := X"8FC20028";
        ram_buffer(57702) := X"00000000";
        ram_buffer(57703) := X"24420001";
        ram_buffer(57704) := X"AFC20028";
        ram_buffer(57705) := X"32420400";
        ram_buffer(57706) := X"10400032";
        ram_buffer(57707) := X"00000000";
        ram_buffer(57708) := X"8FC20024";
        ram_buffer(57709) := X"00000000";
        ram_buffer(57710) := X"80420000";
        ram_buffer(57711) := X"00000000";
        ram_buffer(57712) := X"00401821";
        ram_buffer(57713) := X"8FC20028";
        ram_buffer(57714) := X"00000000";
        ram_buffer(57715) := X"14620029";
        ram_buffer(57716) := X"00000000";
        ram_buffer(57717) := X"8FC20024";
        ram_buffer(57718) := X"00000000";
        ram_buffer(57719) := X"80430000";
        ram_buffer(57720) := X"2402007F";
        ram_buffer(57721) := X"10620023";
        ram_buffer(57722) := X"00000000";
        ram_buffer(57723) := X"8FC20030";
        ram_buffer(57724) := X"00000000";
        ram_buffer(57725) := X"1440000A";
        ram_buffer(57726) := X"00000000";
        ram_buffer(57727) := X"8FC20030";
        ram_buffer(57728) := X"00000000";
        ram_buffer(57729) := X"1440001B";
        ram_buffer(57730) := X"00000000";
        ram_buffer(57731) := X"8FC20034";
        ram_buffer(57732) := X"00000000";
        ram_buffer(57733) := X"2C42000A";
        ram_buffer(57734) := X"14400016";
        ram_buffer(57735) := X"00000000";
        ram_buffer(57736) := X"8FC20020";
        ram_buffer(57737) := X"00000000";
        ram_buffer(57738) := X"00021023";
        ram_buffer(57739) := X"02629821";
        ram_buffer(57740) := X"8FC60020";
        ram_buffer(57741) := X"8FC5001C";
        ram_buffer(57742) := X"02602021";
        ram_buffer(57743) := X"0C02CCBF";
        ram_buffer(57744) := X"00000000";
        ram_buffer(57745) := X"AFC00028";
        ram_buffer(57746) := X"8FC20024";
        ram_buffer(57747) := X"00000000";
        ram_buffer(57748) := X"24420001";
        ram_buffer(57749) := X"80420000";
        ram_buffer(57750) := X"00000000";
        ram_buffer(57751) := X"10400005";
        ram_buffer(57752) := X"00000000";
        ram_buffer(57753) := X"8FC20024";
        ram_buffer(57754) := X"00000000";
        ram_buffer(57755) := X"24420001";
        ram_buffer(57756) := X"AFC20024";
        ram_buffer(57757) := X"8FC30034";
        ram_buffer(57758) := X"8FC20030";
        ram_buffer(57759) := X"2407000A";
        ram_buffer(57760) := X"00003021";
        ram_buffer(57761) := X"00602821";
        ram_buffer(57762) := X"00402021";
        ram_buffer(57763) := X"0C030A67";
        ram_buffer(57764) := X"00000000";
        ram_buffer(57765) := X"AFC30034";
        ram_buffer(57766) := X"AFC20030";
        ram_buffer(57767) := X"8FC20030";
        ram_buffer(57768) := X"8FC30034";
        ram_buffer(57769) := X"00000000";
        ram_buffer(57770) := X"00431025";
        ram_buffer(57771) := X"1440FFAA";
        ram_buffer(57772) := X"00000000";
        ram_buffer(57773) := X"10000029";
        ram_buffer(57774) := X"00000000";
        ram_buffer(57775) := X"2673FFFF";
        ram_buffer(57776) := X"8FC20034";
        ram_buffer(57777) := X"00000000";
        ram_buffer(57778) := X"3043000F";
        ram_buffer(57779) := X"8FC20048";
        ram_buffer(57780) := X"00000000";
        ram_buffer(57781) := X"00431021";
        ram_buffer(57782) := X"80420000";
        ram_buffer(57783) := X"00000000";
        ram_buffer(57784) := X"A2620000";
        ram_buffer(57785) := X"8FC20030";
        ram_buffer(57786) := X"00000000";
        ram_buffer(57787) := X"00021F00";
        ram_buffer(57788) := X"8FC20034";
        ram_buffer(57789) := X"00000000";
        ram_buffer(57790) := X"00021102";
        ram_buffer(57791) := X"00431025";
        ram_buffer(57792) := X"AFC20034";
        ram_buffer(57793) := X"8FC20030";
        ram_buffer(57794) := X"00000000";
        ram_buffer(57795) := X"00021102";
        ram_buffer(57796) := X"AFC20030";
        ram_buffer(57797) := X"8FC20030";
        ram_buffer(57798) := X"8FC30034";
        ram_buffer(57799) := X"00000000";
        ram_buffer(57800) := X"00431025";
        ram_buffer(57801) := X"1440FFE5";
        ram_buffer(57802) := X"00000000";
        ram_buffer(57803) := X"1000000B";
        ram_buffer(57804) := X"00000000";
        ram_buffer(57805) := X"3C02100D";
        ram_buffer(57806) := X"2453ABC8";
        ram_buffer(57807) := X"02602021";
        ram_buffer(57808) := X"0C02851E";
        ram_buffer(57809) := X"00000000";
        ram_buffer(57810) := X"AFC20044";
        ram_buffer(57811) := X"00000000";
        ram_buffer(57812) := X"10000020";
        ram_buffer(57813) := X"00000000";
        ram_buffer(57814) := X"00000000";
        ram_buffer(57815) := X"1000000B";
        ram_buffer(57816) := X"00000000";
        ram_buffer(57817) := X"93C20038";
        ram_buffer(57818) := X"00000000";
        ram_buffer(57819) := X"14400007";
        ram_buffer(57820) := X"00000000";
        ram_buffer(57821) := X"32420001";
        ram_buffer(57822) := X"10400004";
        ram_buffer(57823) := X"00000000";
        ram_buffer(57824) := X"2673FFFF";
        ram_buffer(57825) := X"24020030";
        ram_buffer(57826) := X"A2620000";
        ram_buffer(57827) := X"27C200A8";
        ram_buffer(57828) := X"24420064";
        ram_buffer(57829) := X"00401821";
        ram_buffer(57830) := X"02601021";
        ram_buffer(57831) := X"00621023";
        ram_buffer(57832) := X"AFC20044";
        ram_buffer(57833) := X"1000000B";
        ram_buffer(57834) := X"00000000";
        ram_buffer(57835) := X"128001BA";
        ram_buffer(57836) := X"00000000";
        ram_buffer(57837) := X"27D300A8";
        ram_buffer(57838) := X"00141600";
        ram_buffer(57839) := X"00021603";
        ram_buffer(57840) := X"A2620000";
        ram_buffer(57841) := X"24020001";
        ram_buffer(57842) := X"AFC20044";
        ram_buffer(57843) := X"A3C00058";
        ram_buffer(57844) := X"00000000";
        ram_buffer(57845) := X"8FC4003C";
        ram_buffer(57846) := X"8FC30044";
        ram_buffer(57847) := X"00000000";
        ram_buffer(57848) := X"0064102A";
        ram_buffer(57849) := X"10400002";
        ram_buffer(57850) := X"00000000";
        ram_buffer(57851) := X"00801821";
        ram_buffer(57852) := X"AFC30040";
        ram_buffer(57853) := X"83C20058";
        ram_buffer(57854) := X"00000000";
        ram_buffer(57855) := X"10400005";
        ram_buffer(57856) := X"00000000";
        ram_buffer(57857) := X"8FC20040";
        ram_buffer(57858) := X"00000000";
        ram_buffer(57859) := X"24420001";
        ram_buffer(57860) := X"AFC20040";
        ram_buffer(57861) := X"32420002";
        ram_buffer(57862) := X"10400005";
        ram_buffer(57863) := X"00000000";
        ram_buffer(57864) := X"8FC20040";
        ram_buffer(57865) := X"00000000";
        ram_buffer(57866) := X"24420002";
        ram_buffer(57867) := X"AFC20040";
        ram_buffer(57868) := X"32420084";
        ram_buffer(57869) := X"14400045";
        ram_buffer(57870) := X"00000000";
        ram_buffer(57871) := X"8FC30014";
        ram_buffer(57872) := X"8FC20040";
        ram_buffer(57873) := X"00000000";
        ram_buffer(57874) := X"00628023";
        ram_buffer(57875) := X"1A00003F";
        ram_buffer(57876) := X"00000000";
        ram_buffer(57877) := X"1000001E";
        ram_buffer(57878) := X"00000000";
        ram_buffer(57879) := X"3C02100D";
        ram_buffer(57880) := X"2442AD50";
        ram_buffer(57881) := X"AE220000";
        ram_buffer(57882) := X"24020010";
        ram_buffer(57883) := X"AE220004";
        ram_buffer(57884) := X"8FC20064";
        ram_buffer(57885) := X"00000000";
        ram_buffer(57886) := X"24420010";
        ram_buffer(57887) := X"AFC20064";
        ram_buffer(57888) := X"26310008";
        ram_buffer(57889) := X"8FC20060";
        ram_buffer(57890) := X"00000000";
        ram_buffer(57891) := X"24420001";
        ram_buffer(57892) := X"AFC20060";
        ram_buffer(57893) := X"8FC20060";
        ram_buffer(57894) := X"00000000";
        ram_buffer(57895) := X"28420008";
        ram_buffer(57896) := X"1440000A";
        ram_buffer(57897) := X"00000000";
        ram_buffer(57898) := X"27C2005C";
        ram_buffer(57899) := X"00403021";
        ram_buffer(57900) := X"8FC5018C";
        ram_buffer(57901) := X"8FC40188";
        ram_buffer(57902) := X"0C02DCA6";
        ram_buffer(57903) := X"00000000";
        ram_buffer(57904) := X"14400189";
        ram_buffer(57905) := X"00000000";
        ram_buffer(57906) := X"27D10068";
        ram_buffer(57907) := X"2610FFF0";
        ram_buffer(57908) := X"2A020011";
        ram_buffer(57909) := X"1040FFE1";
        ram_buffer(57910) := X"00000000";
        ram_buffer(57911) := X"3C02100D";
        ram_buffer(57912) := X"2442AD50";
        ram_buffer(57913) := X"AE220000";
        ram_buffer(57914) := X"02001021";
        ram_buffer(57915) := X"AE220004";
        ram_buffer(57916) := X"8FC30064";
        ram_buffer(57917) := X"02001021";
        ram_buffer(57918) := X"00621021";
        ram_buffer(57919) := X"AFC20064";
        ram_buffer(57920) := X"26310008";
        ram_buffer(57921) := X"8FC20060";
        ram_buffer(57922) := X"00000000";
        ram_buffer(57923) := X"24420001";
        ram_buffer(57924) := X"AFC20060";
        ram_buffer(57925) := X"8FC20060";
        ram_buffer(57926) := X"00000000";
        ram_buffer(57927) := X"28420008";
        ram_buffer(57928) := X"1440000A";
        ram_buffer(57929) := X"00000000";
        ram_buffer(57930) := X"27C2005C";
        ram_buffer(57931) := X"00403021";
        ram_buffer(57932) := X"8FC5018C";
        ram_buffer(57933) := X"8FC40188";
        ram_buffer(57934) := X"0C02DCA6";
        ram_buffer(57935) := X"00000000";
        ram_buffer(57936) := X"1440016C";
        ram_buffer(57937) := X"00000000";
        ram_buffer(57938) := X"27D10068";
        ram_buffer(57939) := X"83C20058";
        ram_buffer(57940) := X"00000000";
        ram_buffer(57941) := X"1040001C";
        ram_buffer(57942) := X"00000000";
        ram_buffer(57943) := X"27C20058";
        ram_buffer(57944) := X"AE220000";
        ram_buffer(57945) := X"24020001";
        ram_buffer(57946) := X"AE220004";
        ram_buffer(57947) := X"8FC20064";
        ram_buffer(57948) := X"00000000";
        ram_buffer(57949) := X"24420001";
        ram_buffer(57950) := X"AFC20064";
        ram_buffer(57951) := X"26310008";
        ram_buffer(57952) := X"8FC20060";
        ram_buffer(57953) := X"00000000";
        ram_buffer(57954) := X"24420001";
        ram_buffer(57955) := X"AFC20060";
        ram_buffer(57956) := X"8FC20060";
        ram_buffer(57957) := X"00000000";
        ram_buffer(57958) := X"28420008";
        ram_buffer(57959) := X"1440000A";
        ram_buffer(57960) := X"00000000";
        ram_buffer(57961) := X"27C2005C";
        ram_buffer(57962) := X"00403021";
        ram_buffer(57963) := X"8FC5018C";
        ram_buffer(57964) := X"8FC40188";
        ram_buffer(57965) := X"0C02DCA6";
        ram_buffer(57966) := X"00000000";
        ram_buffer(57967) := X"14400150";
        ram_buffer(57968) := X"00000000";
        ram_buffer(57969) := X"27D10068";
        ram_buffer(57970) := X"32420002";
        ram_buffer(57971) := X"1040001C";
        ram_buffer(57972) := X"00000000";
        ram_buffer(57973) := X"27C2010C";
        ram_buffer(57974) := X"AE220000";
        ram_buffer(57975) := X"24020002";
        ram_buffer(57976) := X"AE220004";
        ram_buffer(57977) := X"8FC20064";
        ram_buffer(57978) := X"00000000";
        ram_buffer(57979) := X"24420002";
        ram_buffer(57980) := X"AFC20064";
        ram_buffer(57981) := X"26310008";
        ram_buffer(57982) := X"8FC20060";
        ram_buffer(57983) := X"00000000";
        ram_buffer(57984) := X"24420001";
        ram_buffer(57985) := X"AFC20060";
        ram_buffer(57986) := X"8FC20060";
        ram_buffer(57987) := X"00000000";
        ram_buffer(57988) := X"28420008";
        ram_buffer(57989) := X"1440000A";
        ram_buffer(57990) := X"00000000";
        ram_buffer(57991) := X"27C2005C";
        ram_buffer(57992) := X"00403021";
        ram_buffer(57993) := X"8FC5018C";
        ram_buffer(57994) := X"8FC40188";
        ram_buffer(57995) := X"0C02DCA6";
        ram_buffer(57996) := X"00000000";
        ram_buffer(57997) := X"14400135";
        ram_buffer(57998) := X"00000000";
        ram_buffer(57999) := X"27D10068";
        ram_buffer(58000) := X"32430084";
        ram_buffer(58001) := X"24020080";
        ram_buffer(58002) := X"14620045";
        ram_buffer(58003) := X"00000000";
        ram_buffer(58004) := X"8FC30014";
        ram_buffer(58005) := X"8FC20040";
        ram_buffer(58006) := X"00000000";
        ram_buffer(58007) := X"00628023";
        ram_buffer(58008) := X"1A00003F";
        ram_buffer(58009) := X"00000000";
        ram_buffer(58010) := X"1000001E";
        ram_buffer(58011) := X"00000000";
        ram_buffer(58012) := X"3C02100D";
        ram_buffer(58013) := X"2442AD60";
        ram_buffer(58014) := X"AE220000";
        ram_buffer(58015) := X"24020010";
        ram_buffer(58016) := X"AE220004";
        ram_buffer(58017) := X"8FC20064";
        ram_buffer(58018) := X"00000000";
        ram_buffer(58019) := X"24420010";
        ram_buffer(58020) := X"AFC20064";
        ram_buffer(58021) := X"26310008";
        ram_buffer(58022) := X"8FC20060";
        ram_buffer(58023) := X"00000000";
        ram_buffer(58024) := X"24420001";
        ram_buffer(58025) := X"AFC20060";
        ram_buffer(58026) := X"8FC20060";
        ram_buffer(58027) := X"00000000";
        ram_buffer(58028) := X"28420008";
        ram_buffer(58029) := X"1440000A";
        ram_buffer(58030) := X"00000000";
        ram_buffer(58031) := X"27C2005C";
        ram_buffer(58032) := X"00403021";
        ram_buffer(58033) := X"8FC5018C";
        ram_buffer(58034) := X"8FC40188";
        ram_buffer(58035) := X"0C02DCA6";
        ram_buffer(58036) := X"00000000";
        ram_buffer(58037) := X"14400110";
        ram_buffer(58038) := X"00000000";
        ram_buffer(58039) := X"27D10068";
        ram_buffer(58040) := X"2610FFF0";
        ram_buffer(58041) := X"2A020011";
        ram_buffer(58042) := X"1040FFE1";
        ram_buffer(58043) := X"00000000";
        ram_buffer(58044) := X"3C02100D";
        ram_buffer(58045) := X"2442AD60";
        ram_buffer(58046) := X"AE220000";
        ram_buffer(58047) := X"02001021";
        ram_buffer(58048) := X"AE220004";
        ram_buffer(58049) := X"8FC30064";
        ram_buffer(58050) := X"02001021";
        ram_buffer(58051) := X"00621021";
        ram_buffer(58052) := X"AFC20064";
        ram_buffer(58053) := X"26310008";
        ram_buffer(58054) := X"8FC20060";
        ram_buffer(58055) := X"00000000";
        ram_buffer(58056) := X"24420001";
        ram_buffer(58057) := X"AFC20060";
        ram_buffer(58058) := X"8FC20060";
        ram_buffer(58059) := X"00000000";
        ram_buffer(58060) := X"28420008";
        ram_buffer(58061) := X"1440000A";
        ram_buffer(58062) := X"00000000";
        ram_buffer(58063) := X"27C2005C";
        ram_buffer(58064) := X"00403021";
        ram_buffer(58065) := X"8FC5018C";
        ram_buffer(58066) := X"8FC40188";
        ram_buffer(58067) := X"0C02DCA6";
        ram_buffer(58068) := X"00000000";
        ram_buffer(58069) := X"144000F3";
        ram_buffer(58070) := X"00000000";
        ram_buffer(58071) := X"27D10068";
        ram_buffer(58072) := X"8FC3003C";
        ram_buffer(58073) := X"8FC20044";
        ram_buffer(58074) := X"00000000";
        ram_buffer(58075) := X"00628023";
        ram_buffer(58076) := X"1A00003F";
        ram_buffer(58077) := X"00000000";
        ram_buffer(58078) := X"1000001E";
        ram_buffer(58079) := X"00000000";
        ram_buffer(58080) := X"3C02100D";
        ram_buffer(58081) := X"2442AD60";
        ram_buffer(58082) := X"AE220000";
        ram_buffer(58083) := X"24020010";
        ram_buffer(58084) := X"AE220004";
        ram_buffer(58085) := X"8FC20064";
        ram_buffer(58086) := X"00000000";
        ram_buffer(58087) := X"24420010";
        ram_buffer(58088) := X"AFC20064";
        ram_buffer(58089) := X"26310008";
        ram_buffer(58090) := X"8FC20060";
        ram_buffer(58091) := X"00000000";
        ram_buffer(58092) := X"24420001";
        ram_buffer(58093) := X"AFC20060";
        ram_buffer(58094) := X"8FC20060";
        ram_buffer(58095) := X"00000000";
        ram_buffer(58096) := X"28420008";
        ram_buffer(58097) := X"1440000A";
        ram_buffer(58098) := X"00000000";
        ram_buffer(58099) := X"27C2005C";
        ram_buffer(58100) := X"00403021";
        ram_buffer(58101) := X"8FC5018C";
        ram_buffer(58102) := X"8FC40188";
        ram_buffer(58103) := X"0C02DCA6";
        ram_buffer(58104) := X"00000000";
        ram_buffer(58105) := X"144000D2";
        ram_buffer(58106) := X"00000000";
        ram_buffer(58107) := X"27D10068";
        ram_buffer(58108) := X"2610FFF0";
        ram_buffer(58109) := X"2A020011";
        ram_buffer(58110) := X"1040FFE1";
        ram_buffer(58111) := X"00000000";
        ram_buffer(58112) := X"3C02100D";
        ram_buffer(58113) := X"2442AD60";
        ram_buffer(58114) := X"AE220000";
        ram_buffer(58115) := X"02001021";
        ram_buffer(58116) := X"AE220004";
        ram_buffer(58117) := X"8FC30064";
        ram_buffer(58118) := X"02001021";
        ram_buffer(58119) := X"00621021";
        ram_buffer(58120) := X"AFC20064";
        ram_buffer(58121) := X"26310008";
        ram_buffer(58122) := X"8FC20060";
        ram_buffer(58123) := X"00000000";
        ram_buffer(58124) := X"24420001";
        ram_buffer(58125) := X"AFC20060";
        ram_buffer(58126) := X"8FC20060";
        ram_buffer(58127) := X"00000000";
        ram_buffer(58128) := X"28420008";
        ram_buffer(58129) := X"1440000A";
        ram_buffer(58130) := X"00000000";
        ram_buffer(58131) := X"27C2005C";
        ram_buffer(58132) := X"00403021";
        ram_buffer(58133) := X"8FC5018C";
        ram_buffer(58134) := X"8FC40188";
        ram_buffer(58135) := X"0C02DCA6";
        ram_buffer(58136) := X"00000000";
        ram_buffer(58137) := X"144000B5";
        ram_buffer(58138) := X"00000000";
        ram_buffer(58139) := X"27D10068";
        ram_buffer(58140) := X"AE330000";
        ram_buffer(58141) := X"8FC20044";
        ram_buffer(58142) := X"00000000";
        ram_buffer(58143) := X"AE220004";
        ram_buffer(58144) := X"8FC30064";
        ram_buffer(58145) := X"8FC20044";
        ram_buffer(58146) := X"00000000";
        ram_buffer(58147) := X"00621021";
        ram_buffer(58148) := X"AFC20064";
        ram_buffer(58149) := X"26310008";
        ram_buffer(58150) := X"8FC20060";
        ram_buffer(58151) := X"00000000";
        ram_buffer(58152) := X"24420001";
        ram_buffer(58153) := X"AFC20060";
        ram_buffer(58154) := X"8FC20060";
        ram_buffer(58155) := X"00000000";
        ram_buffer(58156) := X"28420008";
        ram_buffer(58157) := X"1440000A";
        ram_buffer(58158) := X"00000000";
        ram_buffer(58159) := X"27C2005C";
        ram_buffer(58160) := X"00403021";
        ram_buffer(58161) := X"8FC5018C";
        ram_buffer(58162) := X"8FC40188";
        ram_buffer(58163) := X"0C02DCA6";
        ram_buffer(58164) := X"00000000";
        ram_buffer(58165) := X"1440009C";
        ram_buffer(58166) := X"00000000";
        ram_buffer(58167) := X"27D10068";
        ram_buffer(58168) := X"32420004";
        ram_buffer(58169) := X"10400045";
        ram_buffer(58170) := X"00000000";
        ram_buffer(58171) := X"8FC30014";
        ram_buffer(58172) := X"8FC20040";
        ram_buffer(58173) := X"00000000";
        ram_buffer(58174) := X"00628023";
        ram_buffer(58175) := X"1A00003F";
        ram_buffer(58176) := X"00000000";
        ram_buffer(58177) := X"1000001E";
        ram_buffer(58178) := X"00000000";
        ram_buffer(58179) := X"3C02100D";
        ram_buffer(58180) := X"2442AD50";
        ram_buffer(58181) := X"AE220000";
        ram_buffer(58182) := X"24020010";
        ram_buffer(58183) := X"AE220004";
        ram_buffer(58184) := X"8FC20064";
        ram_buffer(58185) := X"00000000";
        ram_buffer(58186) := X"24420010";
        ram_buffer(58187) := X"AFC20064";
        ram_buffer(58188) := X"26310008";
        ram_buffer(58189) := X"8FC20060";
        ram_buffer(58190) := X"00000000";
        ram_buffer(58191) := X"24420001";
        ram_buffer(58192) := X"AFC20060";
        ram_buffer(58193) := X"8FC20060";
        ram_buffer(58194) := X"00000000";
        ram_buffer(58195) := X"28420008";
        ram_buffer(58196) := X"1440000A";
        ram_buffer(58197) := X"00000000";
        ram_buffer(58198) := X"27C2005C";
        ram_buffer(58199) := X"00403021";
        ram_buffer(58200) := X"8FC5018C";
        ram_buffer(58201) := X"8FC40188";
        ram_buffer(58202) := X"0C02DCA6";
        ram_buffer(58203) := X"00000000";
        ram_buffer(58204) := X"14400078";
        ram_buffer(58205) := X"00000000";
        ram_buffer(58206) := X"27D10068";
        ram_buffer(58207) := X"2610FFF0";
        ram_buffer(58208) := X"2A020011";
        ram_buffer(58209) := X"1040FFE1";
        ram_buffer(58210) := X"00000000";
        ram_buffer(58211) := X"3C02100D";
        ram_buffer(58212) := X"2442AD50";
        ram_buffer(58213) := X"AE220000";
        ram_buffer(58214) := X"02001021";
        ram_buffer(58215) := X"AE220004";
        ram_buffer(58216) := X"8FC20064";
        ram_buffer(58217) := X"02001821";
        ram_buffer(58218) := X"00431021";
        ram_buffer(58219) := X"AFC20064";
        ram_buffer(58220) := X"26310008";
        ram_buffer(58221) := X"8FC20060";
        ram_buffer(58222) := X"00000000";
        ram_buffer(58223) := X"24420001";
        ram_buffer(58224) := X"AFC20060";
        ram_buffer(58225) := X"8FC20060";
        ram_buffer(58226) := X"00000000";
        ram_buffer(58227) := X"28420008";
        ram_buffer(58228) := X"1440000A";
        ram_buffer(58229) := X"00000000";
        ram_buffer(58230) := X"27C2005C";
        ram_buffer(58231) := X"00403021";
        ram_buffer(58232) := X"8FC5018C";
        ram_buffer(58233) := X"8FC40188";
        ram_buffer(58234) := X"0C02DCA6";
        ram_buffer(58235) := X"00000000";
        ram_buffer(58236) := X"1440005B";
        ram_buffer(58237) := X"00000000";
        ram_buffer(58238) := X"27D10068";
        ram_buffer(58239) := X"8FC30014";
        ram_buffer(58240) := X"8FC20040";
        ram_buffer(58241) := X"00000000";
        ram_buffer(58242) := X"0043202A";
        ram_buffer(58243) := X"10800002";
        ram_buffer(58244) := X"00000000";
        ram_buffer(58245) := X"00601021";
        ram_buffer(58246) := X"8FC30010";
        ram_buffer(58247) := X"00000000";
        ram_buffer(58248) := X"00621021";
        ram_buffer(58249) := X"AFC20010";
        ram_buffer(58250) := X"8FC20064";
        ram_buffer(58251) := X"00000000";
        ram_buffer(58252) := X"10400009";
        ram_buffer(58253) := X"00000000";
        ram_buffer(58254) := X"27C2005C";
        ram_buffer(58255) := X"00403021";
        ram_buffer(58256) := X"8FC5018C";
        ram_buffer(58257) := X"8FC40188";
        ram_buffer(58258) := X"0C02DCA6";
        ram_buffer(58259) := X"00000000";
        ram_buffer(58260) := X"14400046";
        ram_buffer(58261) := X"00000000";
        ram_buffer(58262) := X"AFC00060";
        ram_buffer(58263) := X"27D10068";
        ram_buffer(58264) := X"8FC2004C";
        ram_buffer(58265) := X"00000000";
        ram_buffer(58266) := X"1040FA4E";
        ram_buffer(58267) := X"00000000";
        ram_buffer(58268) := X"8FC5004C";
        ram_buffer(58269) := X"8FC40188";
        ram_buffer(58270) := X"0C027301";
        ram_buffer(58271) := X"00000000";
        ram_buffer(58272) := X"AFC0004C";
        ram_buffer(58273) := X"1000FA47";
        ram_buffer(58274) := X"00000000";
        ram_buffer(58275) := X"00000000";
        ram_buffer(58276) := X"10000002";
        ram_buffer(58277) := X"00000000";
        ram_buffer(58278) := X"00000000";
        ram_buffer(58279) := X"8FC20064";
        ram_buffer(58280) := X"00000000";
        ram_buffer(58281) := X"10400009";
        ram_buffer(58282) := X"00000000";
        ram_buffer(58283) := X"27C2005C";
        ram_buffer(58284) := X"00403021";
        ram_buffer(58285) := X"8FC5018C";
        ram_buffer(58286) := X"8FC40188";
        ram_buffer(58287) := X"0C02DCA6";
        ram_buffer(58288) := X"00000000";
        ram_buffer(58289) := X"1440002C";
        ram_buffer(58290) := X"00000000";
        ram_buffer(58291) := X"AFC00060";
        ram_buffer(58292) := X"27D10068";
        ram_buffer(58293) := X"10000029";
        ram_buffer(58294) := X"00000000";
        ram_buffer(58295) := X"00000000";
        ram_buffer(58296) := X"10000026";
        ram_buffer(58297) := X"00000000";
        ram_buffer(58298) := X"00000000";
        ram_buffer(58299) := X"10000023";
        ram_buffer(58300) := X"00000000";
        ram_buffer(58301) := X"00000000";
        ram_buffer(58302) := X"10000020";
        ram_buffer(58303) := X"00000000";
        ram_buffer(58304) := X"00000000";
        ram_buffer(58305) := X"1000001D";
        ram_buffer(58306) := X"00000000";
        ram_buffer(58307) := X"00000000";
        ram_buffer(58308) := X"1000001A";
        ram_buffer(58309) := X"00000000";
        ram_buffer(58310) := X"00000000";
        ram_buffer(58311) := X"10000017";
        ram_buffer(58312) := X"00000000";
        ram_buffer(58313) := X"00000000";
        ram_buffer(58314) := X"10000014";
        ram_buffer(58315) := X"00000000";
        ram_buffer(58316) := X"00000000";
        ram_buffer(58317) := X"10000011";
        ram_buffer(58318) := X"00000000";
        ram_buffer(58319) := X"00000000";
        ram_buffer(58320) := X"1000000E";
        ram_buffer(58321) := X"00000000";
        ram_buffer(58322) := X"00000000";
        ram_buffer(58323) := X"1000000B";
        ram_buffer(58324) := X"00000000";
        ram_buffer(58325) := X"00000000";
        ram_buffer(58326) := X"10000008";
        ram_buffer(58327) := X"00000000";
        ram_buffer(58328) := X"00000000";
        ram_buffer(58329) := X"10000005";
        ram_buffer(58330) := X"00000000";
        ram_buffer(58331) := X"00000000";
        ram_buffer(58332) := X"10000002";
        ram_buffer(58333) := X"00000000";
        ram_buffer(58334) := X"00000000";
        ram_buffer(58335) := X"8FC2004C";
        ram_buffer(58336) := X"00000000";
        ram_buffer(58337) := X"10400005";
        ram_buffer(58338) := X"00000000";
        ram_buffer(58339) := X"8FC5004C";
        ram_buffer(58340) := X"8FC40188";
        ram_buffer(58341) := X"0C027301";
        ram_buffer(58342) := X"00000000";
        ram_buffer(58343) := X"8FC2018C";
        ram_buffer(58344) := X"00000000";
        ram_buffer(58345) := X"8442000C";
        ram_buffer(58346) := X"00000000";
        ram_buffer(58347) := X"3042FFFF";
        ram_buffer(58348) := X"30420040";
        ram_buffer(58349) := X"14400004";
        ram_buffer(58350) := X"00000000";
        ram_buffer(58351) := X"8FC20010";
        ram_buffer(58352) := X"10000003";
        ram_buffer(58353) := X"00000000";
        ram_buffer(58354) := X"2402FFFF";
        ram_buffer(58355) := X"00000000";
        ram_buffer(58356) := X"03C0E821";
        ram_buffer(58357) := X"8FBF0184";
        ram_buffer(58358) := X"8FBE0180";
        ram_buffer(58359) := X"8FB7017C";
        ram_buffer(58360) := X"8FB60178";
        ram_buffer(58361) := X"8FB50174";
        ram_buffer(58362) := X"8FB40170";
        ram_buffer(58363) := X"8FB3016C";
        ram_buffer(58364) := X"8FB20168";
        ram_buffer(58365) := X"8FB10164";
        ram_buffer(58366) := X"8FB00160";
        ram_buffer(58367) := X"27BD0188";
        ram_buffer(58368) := X"03E00008";
        ram_buffer(58369) := X"00000000";
        ram_buffer(58370) := X"27BDFFE0";
        ram_buffer(58371) := X"AFBF001C";
        ram_buffer(58372) := X"AFBE0018";
        ram_buffer(58373) := X"AFB00014";
        ram_buffer(58374) := X"03A0F021";
        ram_buffer(58375) := X"AFC40020";
        ram_buffer(58376) := X"AFC50024";
        ram_buffer(58377) := X"00C08021";
        ram_buffer(58378) := X"8FC30024";
        ram_buffer(58379) := X"2402FFFF";
        ram_buffer(58380) := X"14620004";
        ram_buffer(58381) := X"00000000";
        ram_buffer(58382) := X"2402FFFF";
        ram_buffer(58383) := X"10000060";
        ram_buffer(58384) := X"00000000";
        ram_buffer(58385) := X"8603000C";
        ram_buffer(58386) := X"2402FFDF";
        ram_buffer(58387) := X"00621024";
        ram_buffer(58388) := X"00021400";
        ram_buffer(58389) := X"00021403";
        ram_buffer(58390) := X"A602000C";
        ram_buffer(58391) := X"8FC20024";
        ram_buffer(58392) := X"00000000";
        ram_buffer(58393) := X"304200FF";
        ram_buffer(58394) := X"AFC20024";
        ram_buffer(58395) := X"8E020030";
        ram_buffer(58396) := X"00000000";
        ram_buffer(58397) := X"10400020";
        ram_buffer(58398) := X"00000000";
        ram_buffer(58399) := X"8E030004";
        ram_buffer(58400) := X"8E020034";
        ram_buffer(58401) := X"00000000";
        ram_buffer(58402) := X"0062102A";
        ram_buffer(58403) := X"1440000A";
        ram_buffer(58404) := X"00000000";
        ram_buffer(58405) := X"02002821";
        ram_buffer(58406) := X"8FC40020";
        ram_buffer(58407) := X"0C029C71";
        ram_buffer(58408) := X"00000000";
        ram_buffer(58409) := X"10400004";
        ram_buffer(58410) := X"00000000";
        ram_buffer(58411) := X"2402FFFF";
        ram_buffer(58412) := X"10000043";
        ram_buffer(58413) := X"00000000";
        ram_buffer(58414) := X"8E020000";
        ram_buffer(58415) := X"00000000";
        ram_buffer(58416) := X"2442FFFF";
        ram_buffer(58417) := X"AE020000";
        ram_buffer(58418) := X"8E020000";
        ram_buffer(58419) := X"8FC30024";
        ram_buffer(58420) := X"00000000";
        ram_buffer(58421) := X"306300FF";
        ram_buffer(58422) := X"A0430000";
        ram_buffer(58423) := X"8E020004";
        ram_buffer(58424) := X"00000000";
        ram_buffer(58425) := X"24420001";
        ram_buffer(58426) := X"AE020004";
        ram_buffer(58427) := X"8FC20024";
        ram_buffer(58428) := X"10000033";
        ram_buffer(58429) := X"00000000";
        ram_buffer(58430) := X"8E020010";
        ram_buffer(58431) := X"00000000";
        ram_buffer(58432) := X"1040001C";
        ram_buffer(58433) := X"00000000";
        ram_buffer(58434) := X"8E030000";
        ram_buffer(58435) := X"8E020010";
        ram_buffer(58436) := X"00000000";
        ram_buffer(58437) := X"0043102B";
        ram_buffer(58438) := X"10400016";
        ram_buffer(58439) := X"00000000";
        ram_buffer(58440) := X"8E020000";
        ram_buffer(58441) := X"00000000";
        ram_buffer(58442) := X"2442FFFF";
        ram_buffer(58443) := X"90420000";
        ram_buffer(58444) := X"00000000";
        ram_buffer(58445) := X"00401821";
        ram_buffer(58446) := X"8FC20024";
        ram_buffer(58447) := X"00000000";
        ram_buffer(58448) := X"1462000C";
        ram_buffer(58449) := X"00000000";
        ram_buffer(58450) := X"8E020000";
        ram_buffer(58451) := X"00000000";
        ram_buffer(58452) := X"2442FFFF";
        ram_buffer(58453) := X"AE020000";
        ram_buffer(58454) := X"8E020004";
        ram_buffer(58455) := X"00000000";
        ram_buffer(58456) := X"24420001";
        ram_buffer(58457) := X"AE020004";
        ram_buffer(58458) := X"8FC20024";
        ram_buffer(58459) := X"10000014";
        ram_buffer(58460) := X"00000000";
        ram_buffer(58461) := X"8E020004";
        ram_buffer(58462) := X"00000000";
        ram_buffer(58463) := X"AE02003C";
        ram_buffer(58464) := X"8E020000";
        ram_buffer(58465) := X"00000000";
        ram_buffer(58466) := X"AE020038";
        ram_buffer(58467) := X"26020040";
        ram_buffer(58468) := X"AE020030";
        ram_buffer(58469) := X"24020003";
        ram_buffer(58470) := X"AE020034";
        ram_buffer(58471) := X"8FC20024";
        ram_buffer(58472) := X"00000000";
        ram_buffer(58473) := X"304200FF";
        ram_buffer(58474) := X"A2020042";
        ram_buffer(58475) := X"26020042";
        ram_buffer(58476) := X"AE020000";
        ram_buffer(58477) := X"24020001";
        ram_buffer(58478) := X"AE020004";
        ram_buffer(58479) := X"8FC20024";
        ram_buffer(58480) := X"03C0E821";
        ram_buffer(58481) := X"8FBF001C";
        ram_buffer(58482) := X"8FBE0018";
        ram_buffer(58483) := X"8FB00014";
        ram_buffer(58484) := X"27BD0020";
        ram_buffer(58485) := X"03E00008";
        ram_buffer(58486) := X"00000000";
        ram_buffer(58487) := X"27BDFFE0";
        ram_buffer(58488) := X"AFBF001C";
        ram_buffer(58489) := X"AFBE0018";
        ram_buffer(58490) := X"AFB00014";
        ram_buffer(58491) := X"03A0F021";
        ram_buffer(58492) := X"AFC40020";
        ram_buffer(58493) := X"00A08021";
        ram_buffer(58494) := X"8E020030";
        ram_buffer(58495) := X"00000000";
        ram_buffer(58496) := X"10400019";
        ram_buffer(58497) := X"00000000";
        ram_buffer(58498) := X"8E030030";
        ram_buffer(58499) := X"26020040";
        ram_buffer(58500) := X"10620007";
        ram_buffer(58501) := X"00000000";
        ram_buffer(58502) := X"8E020030";
        ram_buffer(58503) := X"00000000";
        ram_buffer(58504) := X"00402821";
        ram_buffer(58505) := X"8FC40020";
        ram_buffer(58506) := X"0C027301";
        ram_buffer(58507) := X"00000000";
        ram_buffer(58508) := X"AE000030";
        ram_buffer(58509) := X"8E02003C";
        ram_buffer(58510) := X"00000000";
        ram_buffer(58511) := X"AE020004";
        ram_buffer(58512) := X"8E020004";
        ram_buffer(58513) := X"00000000";
        ram_buffer(58514) := X"10400007";
        ram_buffer(58515) := X"00000000";
        ram_buffer(58516) := X"8E020038";
        ram_buffer(58517) := X"00000000";
        ram_buffer(58518) := X"AE020000";
        ram_buffer(58519) := X"00001021";
        ram_buffer(58520) := X"1000000C";
        ram_buffer(58521) := X"00000000";
        ram_buffer(58522) := X"8E020010";
        ram_buffer(58523) := X"00000000";
        ram_buffer(58524) := X"AE020000";
        ram_buffer(58525) := X"AE000004";
        ram_buffer(58526) := X"8602000C";
        ram_buffer(58527) := X"00000000";
        ram_buffer(58528) := X"34420020";
        ram_buffer(58529) := X"00021400";
        ram_buffer(58530) := X"00021403";
        ram_buffer(58531) := X"A602000C";
        ram_buffer(58532) := X"2402FFFF";
        ram_buffer(58533) := X"03C0E821";
        ram_buffer(58534) := X"8FBF001C";
        ram_buffer(58535) := X"8FBE0018";
        ram_buffer(58536) := X"8FB00014";
        ram_buffer(58537) := X"27BD0020";
        ram_buffer(58538) := X"03E00008";
        ram_buffer(58539) := X"00000000";
        ram_buffer(58540) := X"27BDFFD0";
        ram_buffer(58541) := X"AFBF002C";
        ram_buffer(58542) := X"AFBE0028";
        ram_buffer(58543) := X"AFB20024";
        ram_buffer(58544) := X"AFB10020";
        ram_buffer(58545) := X"AFB0001C";
        ram_buffer(58546) := X"03A0F021";
        ram_buffer(58547) := X"AFC40030";
        ram_buffer(58548) := X"AFC50034";
        ram_buffer(58549) := X"AFC60038";
        ram_buffer(58550) := X"AFC7003C";
        ram_buffer(58551) := X"8FC3003C";
        ram_buffer(58552) := X"8FC20038";
        ram_buffer(58553) := X"00000000";
        ram_buffer(58554) := X"00620018";
        ram_buffer(58555) := X"00008012";
        ram_buffer(58556) := X"16000004";
        ram_buffer(58557) := X"00000000";
        ram_buffer(58558) := X"00001021";
        ram_buffer(58559) := X"10000051";
        ram_buffer(58560) := X"00000000";
        ram_buffer(58561) := X"AFD00010";
        ram_buffer(58562) := X"8FD10034";
        ram_buffer(58563) := X"1000002B";
        ram_buffer(58564) := X"00000000";
        ram_buffer(58565) := X"8FC20040";
        ram_buffer(58566) := X"00000000";
        ram_buffer(58567) := X"8C420000";
        ram_buffer(58568) := X"02401821";
        ram_buffer(58569) := X"00603021";
        ram_buffer(58570) := X"00402821";
        ram_buffer(58571) := X"02202021";
        ram_buffer(58572) := X"0C027F93";
        ram_buffer(58573) := X"00000000";
        ram_buffer(58574) := X"8FC20040";
        ram_buffer(58575) := X"00000000";
        ram_buffer(58576) := X"8C420000";
        ram_buffer(58577) := X"02401821";
        ram_buffer(58578) := X"00431821";
        ram_buffer(58579) := X"8FC20040";
        ram_buffer(58580) := X"00000000";
        ram_buffer(58581) := X"AC430000";
        ram_buffer(58582) := X"8FC20040";
        ram_buffer(58583) := X"00000000";
        ram_buffer(58584) := X"AC400004";
        ram_buffer(58585) := X"02401021";
        ram_buffer(58586) := X"02228821";
        ram_buffer(58587) := X"02401021";
        ram_buffer(58588) := X"02028023";
        ram_buffer(58589) := X"8FC50040";
        ram_buffer(58590) := X"8FC40030";
        ram_buffer(58591) := X"0C02E477";
        ram_buffer(58592) := X"00000000";
        ram_buffer(58593) := X"1040000D";
        ram_buffer(58594) := X"00000000";
        ram_buffer(58595) := X"8FC20010";
        ram_buffer(58596) := X"00000000";
        ram_buffer(58597) := X"00501823";
        ram_buffer(58598) := X"8FC20038";
        ram_buffer(58599) := X"00000000";
        ram_buffer(58600) := X"14400002";
        ram_buffer(58601) := X"0062001B";
        ram_buffer(58602) := X"0007000D";
        ram_buffer(58603) := X"00001010";
        ram_buffer(58604) := X"00001012";
        ram_buffer(58605) := X"10000023";
        ram_buffer(58606) := X"00000000";
        ram_buffer(58607) := X"8FC20040";
        ram_buffer(58608) := X"00000000";
        ram_buffer(58609) := X"8C520004";
        ram_buffer(58610) := X"00000000";
        ram_buffer(58611) := X"02401021";
        ram_buffer(58612) := X"0050102B";
        ram_buffer(58613) := X"1440FFCF";
        ram_buffer(58614) := X"00000000";
        ram_buffer(58615) := X"8FC20040";
        ram_buffer(58616) := X"00000000";
        ram_buffer(58617) := X"8C420000";
        ram_buffer(58618) := X"02003021";
        ram_buffer(58619) := X"00402821";
        ram_buffer(58620) := X"02202021";
        ram_buffer(58621) := X"0C027F93";
        ram_buffer(58622) := X"00000000";
        ram_buffer(58623) := X"8FC20040";
        ram_buffer(58624) := X"00000000";
        ram_buffer(58625) := X"8C420004";
        ram_buffer(58626) := X"00000000";
        ram_buffer(58627) := X"00501023";
        ram_buffer(58628) := X"00401821";
        ram_buffer(58629) := X"8FC20040";
        ram_buffer(58630) := X"00000000";
        ram_buffer(58631) := X"AC430004";
        ram_buffer(58632) := X"8FC20040";
        ram_buffer(58633) := X"00000000";
        ram_buffer(58634) := X"8C420000";
        ram_buffer(58635) := X"00000000";
        ram_buffer(58636) := X"00501821";
        ram_buffer(58637) := X"8FC20040";
        ram_buffer(58638) := X"00000000";
        ram_buffer(58639) := X"AC430000";
        ram_buffer(58640) := X"8FC2003C";
        ram_buffer(58641) := X"03C0E821";
        ram_buffer(58642) := X"8FBF002C";
        ram_buffer(58643) := X"8FBE0028";
        ram_buffer(58644) := X"8FB20024";
        ram_buffer(58645) := X"8FB10020";
        ram_buffer(58646) := X"8FB0001C";
        ram_buffer(58647) := X"27BD0030";
        ram_buffer(58648) := X"03E00008";
        ram_buffer(58649) := X"00000000";
        ram_buffer(58650) := X"27BDFE28";
        ram_buffer(58651) := X"AFBF01D4";
        ram_buffer(58652) := X"AFBE01D0";
        ram_buffer(58653) := X"AFB701CC";
        ram_buffer(58654) := X"AFB601C8";
        ram_buffer(58655) := X"AFB501C4";
        ram_buffer(58656) := X"AFB401C0";
        ram_buffer(58657) := X"AFB301BC";
        ram_buffer(58658) := X"AFB201B8";
        ram_buffer(58659) := X"AFB101B4";
        ram_buffer(58660) := X"AFB001B0";
        ram_buffer(58661) := X"03A0F021";
        ram_buffer(58662) := X"AFC401D8";
        ram_buffer(58663) := X"00A08821";
        ram_buffer(58664) := X"AFC601E0";
        ram_buffer(58665) := X"AFC701E4";
        ram_buffer(58666) := X"8FD501E0";
        ram_buffer(58667) := X"AFC00020";
        ram_buffer(58668) := X"24020001";
        ram_buffer(58669) := X"AFC20048";
        ram_buffer(58670) := X"AFC00028";
        ram_buffer(58671) := X"8622000C";
        ram_buffer(58672) := X"00000000";
        ram_buffer(58673) := X"3042FFFF";
        ram_buffer(58674) := X"30422000";
        ram_buffer(58675) := X"1440000B";
        ram_buffer(58676) := X"00000000";
        ram_buffer(58677) := X"8622000C";
        ram_buffer(58678) := X"00000000";
        ram_buffer(58679) := X"34422000";
        ram_buffer(58680) := X"00021400";
        ram_buffer(58681) := X"00021403";
        ram_buffer(58682) := X"A622000C";
        ram_buffer(58683) := X"8E230064";
        ram_buffer(58684) := X"2402DFFF";
        ram_buffer(58685) := X"00621024";
        ram_buffer(58686) := X"AE220064";
        ram_buffer(58687) := X"AFC00018";
        ram_buffer(58688) := X"AFC0001C";
        ram_buffer(58689) := X"92A20000";
        ram_buffer(58690) := X"00000000";
        ram_buffer(58691) := X"AFC20070";
        ram_buffer(58692) := X"8FC20048";
        ram_buffer(58693) := X"00000000";
        ram_buffer(58694) := X"02A2A821";
        ram_buffer(58695) := X"8FC20070";
        ram_buffer(58696) := X"00000000";
        ram_buffer(58697) := X"10400592";
        ram_buffer(58698) := X"00000000";
        ram_buffer(58699) := X"8FC30048";
        ram_buffer(58700) := X"24020001";
        ram_buffer(58701) := X"14620031";
        ram_buffer(58702) := X"00000000";
        ram_buffer(58703) := X"8F838090";
        ram_buffer(58704) := X"8FC20070";
        ram_buffer(58705) := X"00000000";
        ram_buffer(58706) := X"24420001";
        ram_buffer(58707) := X"00621021";
        ram_buffer(58708) := X"80420000";
        ram_buffer(58709) := X"00000000";
        ram_buffer(58710) := X"304200FF";
        ram_buffer(58711) := X"30420008";
        ram_buffer(58712) := X"10400026";
        ram_buffer(58713) := X"00000000";
        ram_buffer(58714) := X"8E220004";
        ram_buffer(58715) := X"00000000";
        ram_buffer(58716) := X"1C400007";
        ram_buffer(58717) := X"00000000";
        ram_buffer(58718) := X"02202821";
        ram_buffer(58719) := X"8FC401D8";
        ram_buffer(58720) := X"0C02E477";
        ram_buffer(58721) := X"00000000";
        ram_buffer(58722) := X"14400547";
        ram_buffer(58723) := X"00000000";
        ram_buffer(58724) := X"8F838090";
        ram_buffer(58725) := X"8E220000";
        ram_buffer(58726) := X"00000000";
        ram_buffer(58727) := X"90420000";
        ram_buffer(58728) := X"00000000";
        ram_buffer(58729) := X"24420001";
        ram_buffer(58730) := X"00621021";
        ram_buffer(58731) := X"80420000";
        ram_buffer(58732) := X"00000000";
        ram_buffer(58733) := X"304200FF";
        ram_buffer(58734) := X"30420008";
        ram_buffer(58735) := X"1040053A";
        ram_buffer(58736) := X"00000000";
        ram_buffer(58737) := X"8FC2001C";
        ram_buffer(58738) := X"00000000";
        ram_buffer(58739) := X"24420001";
        ram_buffer(58740) := X"AFC2001C";
        ram_buffer(58741) := X"8E220004";
        ram_buffer(58742) := X"00000000";
        ram_buffer(58743) := X"2442FFFF";
        ram_buffer(58744) := X"AE220004";
        ram_buffer(58745) := X"8E220000";
        ram_buffer(58746) := X"00000000";
        ram_buffer(58747) := X"24420001";
        ram_buffer(58748) := X"AE220000";
        ram_buffer(58749) := X"1000FFDC";
        ram_buffer(58750) := X"00000000";
        ram_buffer(58751) := X"8FC30070";
        ram_buffer(58752) := X"24020025";
        ram_buffer(58753) := X"14620013";
        ram_buffer(58754) := X"00000000";
        ram_buffer(58755) := X"00009021";
        ram_buffer(58756) := X"00008021";
        ram_buffer(58757) := X"02A01021";
        ram_buffer(58758) := X"24550001";
        ram_buffer(58759) := X"90420000";
        ram_buffer(58760) := X"00000000";
        ram_buffer(58761) := X"00409821";
        ram_buffer(58762) := X"2E62007B";
        ram_buffer(58763) := X"10400109";
        ram_buffer(58764) := X"00000000";
        ram_buffer(58765) := X"00131880";
        ram_buffer(58766) := X"3C02100D";
        ram_buffer(58767) := X"2442AD70";
        ram_buffer(58768) := X"00621021";
        ram_buffer(58769) := X"8C420000";
        ram_buffer(58770) := X"00000000";
        ram_buffer(58771) := X"00400008";
        ram_buffer(58772) := X"00000000";
        ram_buffer(58773) := X"00000000";
        ram_buffer(58774) := X"8FC20048";
        ram_buffer(58775) := X"00000000";
        ram_buffer(58776) := X"00021023";
        ram_buffer(58777) := X"02A21021";
        ram_buffer(58778) := X"AFC2002C";
        ram_buffer(58779) := X"00009821";
        ram_buffer(58780) := X"10000025";
        ram_buffer(58781) := X"00000000";
        ram_buffer(58782) := X"8E220004";
        ram_buffer(58783) := X"00000000";
        ram_buffer(58784) := X"1C400007";
        ram_buffer(58785) := X"00000000";
        ram_buffer(58786) := X"02202821";
        ram_buffer(58787) := X"8FC401D8";
        ram_buffer(58788) := X"0C02E477";
        ram_buffer(58789) := X"00000000";
        ram_buffer(58790) := X"1440050F";
        ram_buffer(58791) := X"00000000";
        ram_buffer(58792) := X"8E220000";
        ram_buffer(58793) := X"00000000";
        ram_buffer(58794) := X"90430000";
        ram_buffer(58795) := X"8FC2002C";
        ram_buffer(58796) := X"00000000";
        ram_buffer(58797) := X"90420000";
        ram_buffer(58798) := X"00000000";
        ram_buffer(58799) := X"1462052F";
        ram_buffer(58800) := X"00000000";
        ram_buffer(58801) := X"8E220004";
        ram_buffer(58802) := X"00000000";
        ram_buffer(58803) := X"2442FFFF";
        ram_buffer(58804) := X"AE220004";
        ram_buffer(58805) := X"8E220000";
        ram_buffer(58806) := X"00000000";
        ram_buffer(58807) := X"24420001";
        ram_buffer(58808) := X"AE220000";
        ram_buffer(58809) := X"8FC2001C";
        ram_buffer(58810) := X"00000000";
        ram_buffer(58811) := X"24420001";
        ram_buffer(58812) := X"AFC2001C";
        ram_buffer(58813) := X"8FC2002C";
        ram_buffer(58814) := X"00000000";
        ram_buffer(58815) := X"24420001";
        ram_buffer(58816) := X"AFC2002C";
        ram_buffer(58817) := X"26730001";
        ram_buffer(58818) := X"8FC20048";
        ram_buffer(58819) := X"00000000";
        ram_buffer(58820) := X"0262102A";
        ram_buffer(58821) := X"1440FFD8";
        ram_buffer(58822) := X"00000000";
        ram_buffer(58823) := X"100004EC";
        ram_buffer(58824) := X"00000000";
        ram_buffer(58825) := X"36100010";
        ram_buffer(58826) := X"1000FFBA";
        ram_buffer(58827) := X"00000000";
        ram_buffer(58828) := X"92A30000";
        ram_buffer(58829) := X"2402006C";
        ram_buffer(58830) := X"14620005";
        ram_buffer(58831) := X"00000000";
        ram_buffer(58832) := X"26B50001";
        ram_buffer(58833) := X"36100002";
        ram_buffer(58834) := X"1000FFB2";
        ram_buffer(58835) := X"00000000";
        ram_buffer(58836) := X"36100001";
        ram_buffer(58837) := X"1000FFAF";
        ram_buffer(58838) := X"00000000";
        ram_buffer(58839) := X"36100002";
        ram_buffer(58840) := X"1000FFAC";
        ram_buffer(58841) := X"00000000";
        ram_buffer(58842) := X"92A30000";
        ram_buffer(58843) := X"24020068";
        ram_buffer(58844) := X"14620005";
        ram_buffer(58845) := X"00000000";
        ram_buffer(58846) := X"26B50001";
        ram_buffer(58847) := X"36100008";
        ram_buffer(58848) := X"1000FFA4";
        ram_buffer(58849) := X"00000000";
        ram_buffer(58850) := X"36100004";
        ram_buffer(58851) := X"1000FFA1";
        ram_buffer(58852) := X"00000000";
        ram_buffer(58853) := X"36100002";
        ram_buffer(58854) := X"1000FF9E";
        ram_buffer(58855) := X"00000000";
        ram_buffer(58856) := X"02401021";
        ram_buffer(58857) := X"00021040";
        ram_buffer(58858) := X"00021880";
        ram_buffer(58859) := X"00431021";
        ram_buffer(58860) := X"02601821";
        ram_buffer(58861) := X"00431021";
        ram_buffer(58862) := X"2452FFD0";
        ram_buffer(58863) := X"1000FF95";
        ram_buffer(58864) := X"00000000";
        ram_buffer(58865) := X"36100001";
        ram_buffer(58866) := X"24130003";
        ram_buffer(58867) := X"3C02100B";
        ram_buffer(58868) := X"24426198";
        ram_buffer(58869) := X"AFC20028";
        ram_buffer(58870) := X"2402000A";
        ram_buffer(58871) := X"AFC20020";
        ram_buffer(58872) := X"100000AF";
        ram_buffer(58873) := X"00000000";
        ram_buffer(58874) := X"24130003";
        ram_buffer(58875) := X"3C02100B";
        ram_buffer(58876) := X"24426198";
        ram_buffer(58877) := X"AFC20028";
        ram_buffer(58878) := X"AFC00020";
        ram_buffer(58879) := X"100000A8";
        ram_buffer(58880) := X"00000000";
        ram_buffer(58881) := X"36100001";
        ram_buffer(58882) := X"24130003";
        ram_buffer(58883) := X"3C02100B";
        ram_buffer(58884) := X"24426A64";
        ram_buffer(58885) := X"AFC20028";
        ram_buffer(58886) := X"24020008";
        ram_buffer(58887) := X"AFC20020";
        ram_buffer(58888) := X"1000009F";
        ram_buffer(58889) := X"00000000";
        ram_buffer(58890) := X"24130003";
        ram_buffer(58891) := X"3C02100B";
        ram_buffer(58892) := X"24426A64";
        ram_buffer(58893) := X"AFC20028";
        ram_buffer(58894) := X"2402000A";
        ram_buffer(58895) := X"AFC20020";
        ram_buffer(58896) := X"10000097";
        ram_buffer(58897) := X"00000000";
        ram_buffer(58898) := X"36100200";
        ram_buffer(58899) := X"24130003";
        ram_buffer(58900) := X"3C02100B";
        ram_buffer(58901) := X"24426A64";
        ram_buffer(58902) := X"AFC20028";
        ram_buffer(58903) := X"24020010";
        ram_buffer(58904) := X"AFC20020";
        ram_buffer(58905) := X"1000008E";
        ram_buffer(58906) := X"00000000";
        ram_buffer(58907) := X"36100001";
        ram_buffer(58908) := X"24130002";
        ram_buffer(58909) := X"1000008A";
        ram_buffer(58910) := X"00000000";
        ram_buffer(58911) := X"27C20074";
        ram_buffer(58912) := X"02A02821";
        ram_buffer(58913) := X"00402021";
        ram_buffer(58914) := X"0C02CBBB";
        ram_buffer(58915) := X"00000000";
        ram_buffer(58916) := X"0040A821";
        ram_buffer(58917) := X"36100040";
        ram_buffer(58918) := X"24130001";
        ram_buffer(58919) := X"10000080";
        ram_buffer(58920) := X"00000000";
        ram_buffer(58921) := X"36100001";
        ram_buffer(58922) := X"36100040";
        ram_buffer(58923) := X"00009821";
        ram_buffer(58924) := X"1000007B";
        ram_buffer(58925) := X"00000000";
        ram_buffer(58926) := X"36100220";
        ram_buffer(58927) := X"24130003";
        ram_buffer(58928) := X"3C02100B";
        ram_buffer(58929) := X"24426A64";
        ram_buffer(58930) := X"AFC20028";
        ram_buffer(58931) := X"24020010";
        ram_buffer(58932) := X"AFC20020";
        ram_buffer(58933) := X"10000072";
        ram_buffer(58934) := X"00000000";
        ram_buffer(58935) := X"32020010";
        ram_buffer(58936) := X"14400474";
        ram_buffer(58937) := X"00000000";
        ram_buffer(58938) := X"32020008";
        ram_buffer(58939) := X"10400011";
        ram_buffer(58940) := X"00000000";
        ram_buffer(58941) := X"8FC201E4";
        ram_buffer(58942) := X"00000000";
        ram_buffer(58943) := X"24430004";
        ram_buffer(58944) := X"AFC301E4";
        ram_buffer(58945) := X"8C420000";
        ram_buffer(58946) := X"00000000";
        ram_buffer(58947) := X"AFC2004C";
        ram_buffer(58948) := X"8FC2001C";
        ram_buffer(58949) := X"00000000";
        ram_buffer(58950) := X"00021E00";
        ram_buffer(58951) := X"00031E03";
        ram_buffer(58952) := X"8FC2004C";
        ram_buffer(58953) := X"00000000";
        ram_buffer(58954) := X"A0430000";
        ram_buffer(58955) := X"10000468";
        ram_buffer(58956) := X"00000000";
        ram_buffer(58957) := X"32020004";
        ram_buffer(58958) := X"10400011";
        ram_buffer(58959) := X"00000000";
        ram_buffer(58960) := X"8FC201E4";
        ram_buffer(58961) := X"00000000";
        ram_buffer(58962) := X"24430004";
        ram_buffer(58963) := X"AFC301E4";
        ram_buffer(58964) := X"8C420000";
        ram_buffer(58965) := X"00000000";
        ram_buffer(58966) := X"AFC20050";
        ram_buffer(58967) := X"8FC2001C";
        ram_buffer(58968) := X"00000000";
        ram_buffer(58969) := X"00021C00";
        ram_buffer(58970) := X"00031C03";
        ram_buffer(58971) := X"8FC20050";
        ram_buffer(58972) := X"00000000";
        ram_buffer(58973) := X"A4430000";
        ram_buffer(58974) := X"10000455";
        ram_buffer(58975) := X"00000000";
        ram_buffer(58976) := X"32020001";
        ram_buffer(58977) := X"1040000E";
        ram_buffer(58978) := X"00000000";
        ram_buffer(58979) := X"8FC201E4";
        ram_buffer(58980) := X"00000000";
        ram_buffer(58981) := X"24430004";
        ram_buffer(58982) := X"AFC301E4";
        ram_buffer(58983) := X"8C420000";
        ram_buffer(58984) := X"00000000";
        ram_buffer(58985) := X"AFC20054";
        ram_buffer(58986) := X"8FC20054";
        ram_buffer(58987) := X"8FC3001C";
        ram_buffer(58988) := X"00000000";
        ram_buffer(58989) := X"AC430000";
        ram_buffer(58990) := X"10000445";
        ram_buffer(58991) := X"00000000";
        ram_buffer(58992) := X"32020002";
        ram_buffer(58993) := X"10400013";
        ram_buffer(58994) := X"00000000";
        ram_buffer(58995) := X"8FC201E4";
        ram_buffer(58996) := X"00000000";
        ram_buffer(58997) := X"24430004";
        ram_buffer(58998) := X"AFC301E4";
        ram_buffer(58999) := X"8C420000";
        ram_buffer(59000) := X"00000000";
        ram_buffer(59001) := X"AFC20058";
        ram_buffer(59002) := X"8FC2001C";
        ram_buffer(59003) := X"00000000";
        ram_buffer(59004) := X"0040B821";
        ram_buffer(59005) := X"000217C3";
        ram_buffer(59006) := X"0040B021";
        ram_buffer(59007) := X"8FC20058";
        ram_buffer(59008) := X"00000000";
        ram_buffer(59009) := X"AC570004";
        ram_buffer(59010) := X"AC560000";
        ram_buffer(59011) := X"10000430";
        ram_buffer(59012) := X"00000000";
        ram_buffer(59013) := X"8FC201E4";
        ram_buffer(59014) := X"00000000";
        ram_buffer(59015) := X"24430004";
        ram_buffer(59016) := X"AFC301E4";
        ram_buffer(59017) := X"8C420000";
        ram_buffer(59018) := X"00000000";
        ram_buffer(59019) := X"AFC2005C";
        ram_buffer(59020) := X"8FC2005C";
        ram_buffer(59021) := X"8FC3001C";
        ram_buffer(59022) := X"00000000";
        ram_buffer(59023) := X"AC430000";
        ram_buffer(59024) := X"10000423";
        ram_buffer(59025) := X"00000000";
        ram_buffer(59026) := X"2402FFFF";
        ram_buffer(59027) := X"10000453";
        ram_buffer(59028) := X"00000000";
        ram_buffer(59029) := X"8F838090";
        ram_buffer(59030) := X"02601021";
        ram_buffer(59031) := X"24420001";
        ram_buffer(59032) := X"00621021";
        ram_buffer(59033) := X"80420000";
        ram_buffer(59034) := X"00000000";
        ram_buffer(59035) := X"304200FF";
        ram_buffer(59036) := X"30430003";
        ram_buffer(59037) := X"24020001";
        ram_buffer(59038) := X"14620002";
        ram_buffer(59039) := X"00000000";
        ram_buffer(59040) := X"36100001";
        ram_buffer(59041) := X"24130003";
        ram_buffer(59042) := X"3C02100B";
        ram_buffer(59043) := X"24426198";
        ram_buffer(59044) := X"AFC20028";
        ram_buffer(59045) := X"2402000A";
        ram_buffer(59046) := X"AFC20020";
        ram_buffer(59047) := X"00000000";
        ram_buffer(59048) := X"8E220004";
        ram_buffer(59049) := X"00000000";
        ram_buffer(59050) := X"1C400007";
        ram_buffer(59051) := X"00000000";
        ram_buffer(59052) := X"02202821";
        ram_buffer(59053) := X"8FC401D8";
        ram_buffer(59054) := X"0C02E477";
        ram_buffer(59055) := X"00000000";
        ram_buffer(59056) := X"14400408";
        ram_buffer(59057) := X"00000000";
        ram_buffer(59058) := X"32020040";
        ram_buffer(59059) := X"14400028";
        ram_buffer(59060) := X"00000000";
        ram_buffer(59061) := X"10000019";
        ram_buffer(59062) := X"00000000";
        ram_buffer(59063) := X"8FC2001C";
        ram_buffer(59064) := X"00000000";
        ram_buffer(59065) := X"24420001";
        ram_buffer(59066) := X"AFC2001C";
        ram_buffer(59067) := X"8E220004";
        ram_buffer(59068) := X"00000000";
        ram_buffer(59069) := X"2442FFFF";
        ram_buffer(59070) := X"AE220004";
        ram_buffer(59071) := X"8E220004";
        ram_buffer(59072) := X"00000000";
        ram_buffer(59073) := X"18400007";
        ram_buffer(59074) := X"00000000";
        ram_buffer(59075) := X"8E220000";
        ram_buffer(59076) := X"00000000";
        ram_buffer(59077) := X"24420001";
        ram_buffer(59078) := X"AE220000";
        ram_buffer(59079) := X"10000007";
        ram_buffer(59080) := X"00000000";
        ram_buffer(59081) := X"02202821";
        ram_buffer(59082) := X"8FC401D8";
        ram_buffer(59083) := X"0C02E477";
        ram_buffer(59084) := X"00000000";
        ram_buffer(59085) := X"144003EE";
        ram_buffer(59086) := X"00000000";
        ram_buffer(59087) := X"8F838090";
        ram_buffer(59088) := X"8E220000";
        ram_buffer(59089) := X"00000000";
        ram_buffer(59090) := X"90420000";
        ram_buffer(59091) := X"00000000";
        ram_buffer(59092) := X"24420001";
        ram_buffer(59093) := X"00621021";
        ram_buffer(59094) := X"80420000";
        ram_buffer(59095) := X"00000000";
        ram_buffer(59096) := X"304200FF";
        ram_buffer(59097) := X"30420008";
        ram_buffer(59098) := X"1440FFDC";
        ram_buffer(59099) := X"00000000";
        ram_buffer(59100) := X"24020001";
        ram_buffer(59101) := X"126200DB";
        ram_buffer(59102) := X"00000000";
        ram_buffer(59103) := X"2A620002";
        ram_buffer(59104) := X"10400005";
        ram_buffer(59105) := X"00000000";
        ram_buffer(59106) := X"1260000B";
        ram_buffer(59107) := X"00000000";
        ram_buffer(59108) := X"100003CF";
        ram_buffer(59109) := X"00000000";
        ram_buffer(59110) := X"24020002";
        ram_buffer(59111) := X"12620153";
        ram_buffer(59112) := X"00000000";
        ram_buffer(59113) := X"24020003";
        ram_buffer(59114) := X"1262026C";
        ram_buffer(59115) := X"00000000";
        ram_buffer(59116) := X"100003C7";
        ram_buffer(59117) := X"00000000";
        ram_buffer(59118) := X"16400002";
        ram_buffer(59119) := X"00000000";
        ram_buffer(59120) := X"24120001";
        ram_buffer(59121) := X"32020001";
        ram_buffer(59122) := X"10400074";
        ram_buffer(59123) := X"00000000";
        ram_buffer(59124) := X"27C2019C";
        ram_buffer(59125) := X"24060008";
        ram_buffer(59126) := X"00002821";
        ram_buffer(59127) := X"00402021";
        ram_buffer(59128) := X"0C02801D";
        ram_buffer(59129) := X"00000000";
        ram_buffer(59130) := X"32020010";
        ram_buffer(59131) := X"1440000A";
        ram_buffer(59132) := X"00000000";
        ram_buffer(59133) := X"8FC201E4";
        ram_buffer(59134) := X"00000000";
        ram_buffer(59135) := X"24430004";
        ram_buffer(59136) := X"AFC301E4";
        ram_buffer(59137) := X"8C420000";
        ram_buffer(59138) := X"00000000";
        ram_buffer(59139) := X"AFC20024";
        ram_buffer(59140) := X"10000002";
        ram_buffer(59141) := X"00000000";
        ram_buffer(59142) := X"AFC00024";
        ram_buffer(59143) := X"00009821";
        ram_buffer(59144) := X"10000050";
        ram_buffer(59145) := X"00000000";
        ram_buffer(59146) := X"0C02BB09";
        ram_buffer(59147) := X"00000000";
        ram_buffer(59148) := X"105303B2";
        ram_buffer(59149) := X"00000000";
        ram_buffer(59150) := X"02601021";
        ram_buffer(59151) := X"24530001";
        ram_buffer(59152) := X"8E230000";
        ram_buffer(59153) := X"00000000";
        ram_buffer(59154) := X"90630000";
        ram_buffer(59155) := X"00000000";
        ram_buffer(59156) := X"00031E00";
        ram_buffer(59157) := X"00031E03";
        ram_buffer(59158) := X"27C40018";
        ram_buffer(59159) := X"00821021";
        ram_buffer(59160) := X"A043015C";
        ram_buffer(59161) := X"8E220004";
        ram_buffer(59162) := X"00000000";
        ram_buffer(59163) := X"2442FFFF";
        ram_buffer(59164) := X"AE220004";
        ram_buffer(59165) := X"8E220000";
        ram_buffer(59166) := X"00000000";
        ram_buffer(59167) := X"24420001";
        ram_buffer(59168) := X"AE220000";
        ram_buffer(59169) := X"02602021";
        ram_buffer(59170) := X"27C30174";
        ram_buffer(59171) := X"27C2019C";
        ram_buffer(59172) := X"AFA20010";
        ram_buffer(59173) := X"00803821";
        ram_buffer(59174) := X"00603021";
        ram_buffer(59175) := X"8FC50024";
        ram_buffer(59176) := X"8FC401D8";
        ram_buffer(59177) := X"0C02BB73";
        ram_buffer(59178) := X"00000000";
        ram_buffer(59179) := X"AFC20060";
        ram_buffer(59180) := X"8FC30060";
        ram_buffer(59181) := X"2402FFFF";
        ram_buffer(59182) := X"10620393";
        ram_buffer(59183) := X"00000000";
        ram_buffer(59184) := X"8FC20060";
        ram_buffer(59185) := X"00000000";
        ram_buffer(59186) := X"14400007";
        ram_buffer(59187) := X"00000000";
        ram_buffer(59188) := X"32020010";
        ram_buffer(59189) := X"14400004";
        ram_buffer(59190) := X"00000000";
        ram_buffer(59191) := X"8FC20024";
        ram_buffer(59192) := X"00000000";
        ram_buffer(59193) := X"AC400000";
        ram_buffer(59194) := X"8FC30060";
        ram_buffer(59195) := X"2402FFFE";
        ram_buffer(59196) := X"1062000E";
        ram_buffer(59197) := X"00000000";
        ram_buffer(59198) := X"8FC2001C";
        ram_buffer(59199) := X"00000000";
        ram_buffer(59200) := X"00531021";
        ram_buffer(59201) := X"AFC2001C";
        ram_buffer(59202) := X"2652FFFF";
        ram_buffer(59203) := X"32020010";
        ram_buffer(59204) := X"14400005";
        ram_buffer(59205) := X"00000000";
        ram_buffer(59206) := X"8FC20024";
        ram_buffer(59207) := X"00000000";
        ram_buffer(59208) := X"24420004";
        ram_buffer(59209) := X"AFC20024";
        ram_buffer(59210) := X"00009821";
        ram_buffer(59211) := X"8E220004";
        ram_buffer(59212) := X"00000000";
        ram_buffer(59213) := X"1C40000B";
        ram_buffer(59214) := X"00000000";
        ram_buffer(59215) := X"02202821";
        ram_buffer(59216) := X"8FC401D8";
        ram_buffer(59217) := X"0C02E477";
        ram_buffer(59218) := X"00000000";
        ram_buffer(59219) := X"10400005";
        ram_buffer(59220) := X"00000000";
        ram_buffer(59221) := X"12600007";
        ram_buffer(59222) := X"00000000";
        ram_buffer(59223) := X"10000374";
        ram_buffer(59224) := X"00000000";
        ram_buffer(59225) := X"1640FFB0";
        ram_buffer(59226) := X"00000000";
        ram_buffer(59227) := X"10000002";
        ram_buffer(59228) := X"00000000";
        ram_buffer(59229) := X"00000000";
        ram_buffer(59230) := X"32020010";
        ram_buffer(59231) := X"14400350";
        ram_buffer(59232) := X"00000000";
        ram_buffer(59233) := X"8FC20018";
        ram_buffer(59234) := X"00000000";
        ram_buffer(59235) := X"24420001";
        ram_buffer(59236) := X"AFC20018";
        ram_buffer(59237) := X"1000034A";
        ram_buffer(59238) := X"00000000";
        ram_buffer(59239) := X"32020010";
        ram_buffer(59240) := X"10400034";
        ram_buffer(59241) := X"00000000";
        ram_buffer(59242) := X"AFC00030";
        ram_buffer(59243) := X"8E330004";
        ram_buffer(59244) := X"02401021";
        ram_buffer(59245) := X"0262102A";
        ram_buffer(59246) := X"10400018";
        ram_buffer(59247) := X"00000000";
        ram_buffer(59248) := X"02601821";
        ram_buffer(59249) := X"8FC20030";
        ram_buffer(59250) := X"00000000";
        ram_buffer(59251) := X"00431021";
        ram_buffer(59252) := X"AFC20030";
        ram_buffer(59253) := X"02601021";
        ram_buffer(59254) := X"02429023";
        ram_buffer(59255) := X"8E220000";
        ram_buffer(59256) := X"02601821";
        ram_buffer(59257) := X"00431021";
        ram_buffer(59258) := X"AE220000";
        ram_buffer(59259) := X"02202821";
        ram_buffer(59260) := X"8FC401D8";
        ram_buffer(59261) := X"0C02E477";
        ram_buffer(59262) := X"00000000";
        ram_buffer(59263) := X"1040FFEB";
        ram_buffer(59264) := X"00000000";
        ram_buffer(59265) := X"8FC20030";
        ram_buffer(59266) := X"00000000";
        ram_buffer(59267) := X"14400011";
        ram_buffer(59268) := X"00000000";
        ram_buffer(59269) := X"10000346";
        ram_buffer(59270) := X"00000000";
        ram_buffer(59271) := X"8FC20030";
        ram_buffer(59272) := X"00000000";
        ram_buffer(59273) := X"00521021";
        ram_buffer(59274) := X"AFC20030";
        ram_buffer(59275) := X"8E220004";
        ram_buffer(59276) := X"00000000";
        ram_buffer(59277) := X"00521023";
        ram_buffer(59278) := X"AE220004";
        ram_buffer(59279) := X"8E220000";
        ram_buffer(59280) := X"00000000";
        ram_buffer(59281) := X"00521021";
        ram_buffer(59282) := X"AE220000";
        ram_buffer(59283) := X"10000002";
        ram_buffer(59284) := X"00000000";
        ram_buffer(59285) := X"00000000";
        ram_buffer(59286) := X"8FC3001C";
        ram_buffer(59287) := X"8FC20030";
        ram_buffer(59288) := X"00000000";
        ram_buffer(59289) := X"00621021";
        ram_buffer(59290) := X"AFC2001C";
        ram_buffer(59291) := X"10000314";
        ram_buffer(59292) := X"00000000";
        ram_buffer(59293) := X"8FC201E4";
        ram_buffer(59294) := X"00000000";
        ram_buffer(59295) := X"24430004";
        ram_buffer(59296) := X"AFC301E4";
        ram_buffer(59297) := X"8C420000";
        ram_buffer(59298) := X"AFB10010";
        ram_buffer(59299) := X"02403821";
        ram_buffer(59300) := X"24060001";
        ram_buffer(59301) := X"00402821";
        ram_buffer(59302) := X"8FC401D8";
        ram_buffer(59303) := X"0C02E4AC";
        ram_buffer(59304) := X"00000000";
        ram_buffer(59305) := X"AFC20064";
        ram_buffer(59306) := X"8FC20064";
        ram_buffer(59307) := X"00000000";
        ram_buffer(59308) := X"10400318";
        ram_buffer(59309) := X"00000000";
        ram_buffer(59310) := X"8FC3001C";
        ram_buffer(59311) := X"8FC20064";
        ram_buffer(59312) := X"00000000";
        ram_buffer(59313) := X"00621021";
        ram_buffer(59314) := X"AFC2001C";
        ram_buffer(59315) := X"8FC20018";
        ram_buffer(59316) := X"00000000";
        ram_buffer(59317) := X"24420001";
        ram_buffer(59318) := X"AFC20018";
        ram_buffer(59319) := X"100002F8";
        ram_buffer(59320) := X"00000000";
        ram_buffer(59321) := X"16400002";
        ram_buffer(59322) := X"00000000";
        ram_buffer(59323) := X"2412FFFF";
        ram_buffer(59324) := X"32020010";
        ram_buffer(59325) := X"10400033";
        ram_buffer(59326) := X"00000000";
        ram_buffer(59327) := X"00009821";
        ram_buffer(59328) := X"1000001B";
        ram_buffer(59329) := X"00000000";
        ram_buffer(59330) := X"26730001";
        ram_buffer(59331) := X"8E220004";
        ram_buffer(59332) := X"00000000";
        ram_buffer(59333) := X"2442FFFF";
        ram_buffer(59334) := X"AE220004";
        ram_buffer(59335) := X"8E220000";
        ram_buffer(59336) := X"00000000";
        ram_buffer(59337) := X"24420001";
        ram_buffer(59338) := X"AE220000";
        ram_buffer(59339) := X"2652FFFF";
        ram_buffer(59340) := X"1240001C";
        ram_buffer(59341) := X"00000000";
        ram_buffer(59342) := X"8E220004";
        ram_buffer(59343) := X"00000000";
        ram_buffer(59344) := X"1C40000B";
        ram_buffer(59345) := X"00000000";
        ram_buffer(59346) := X"02202821";
        ram_buffer(59347) := X"8FC401D8";
        ram_buffer(59348) := X"0C02E477";
        ram_buffer(59349) := X"00000000";
        ram_buffer(59350) := X"10400005";
        ram_buffer(59351) := X"00000000";
        ram_buffer(59352) := X"16600013";
        ram_buffer(59353) := X"00000000";
        ram_buffer(59354) := X"100002F1";
        ram_buffer(59355) := X"00000000";
        ram_buffer(59356) := X"8E220000";
        ram_buffer(59357) := X"00000000";
        ram_buffer(59358) := X"90420000";
        ram_buffer(59359) := X"00000000";
        ram_buffer(59360) := X"00401821";
        ram_buffer(59361) := X"27C20018";
        ram_buffer(59362) := X"00431021";
        ram_buffer(59363) := X"8042005C";
        ram_buffer(59364) := X"00000000";
        ram_buffer(59365) := X"1440FFDC";
        ram_buffer(59366) := X"00000000";
        ram_buffer(59367) := X"10000005";
        ram_buffer(59368) := X"00000000";
        ram_buffer(59369) := X"00000000";
        ram_buffer(59370) := X"10000002";
        ram_buffer(59371) := X"00000000";
        ram_buffer(59372) := X"00000000";
        ram_buffer(59373) := X"16600047";
        ram_buffer(59374) := X"00000000";
        ram_buffer(59375) := X"100002F6";
        ram_buffer(59376) := X"00000000";
        ram_buffer(59377) := X"8FC201E4";
        ram_buffer(59378) := X"00000000";
        ram_buffer(59379) := X"24430004";
        ram_buffer(59380) := X"AFC301E4";
        ram_buffer(59381) := X"8C540000";
        ram_buffer(59382) := X"00000000";
        ram_buffer(59383) := X"02808021";
        ram_buffer(59384) := X"10000021";
        ram_buffer(59385) := X"00000000";
        ram_buffer(59386) := X"8E220004";
        ram_buffer(59387) := X"00000000";
        ram_buffer(59388) := X"2442FFFF";
        ram_buffer(59389) := X"AE220004";
        ram_buffer(59390) := X"02801821";
        ram_buffer(59391) := X"24740001";
        ram_buffer(59392) := X"8E220000";
        ram_buffer(59393) := X"00000000";
        ram_buffer(59394) := X"24440001";
        ram_buffer(59395) := X"AE240000";
        ram_buffer(59396) := X"90420000";
        ram_buffer(59397) := X"00000000";
        ram_buffer(59398) := X"00021600";
        ram_buffer(59399) := X"00021603";
        ram_buffer(59400) := X"A0620000";
        ram_buffer(59401) := X"2652FFFF";
        ram_buffer(59402) := X"1240001C";
        ram_buffer(59403) := X"00000000";
        ram_buffer(59404) := X"8E220004";
        ram_buffer(59405) := X"00000000";
        ram_buffer(59406) := X"1C40000B";
        ram_buffer(59407) := X"00000000";
        ram_buffer(59408) := X"02202821";
        ram_buffer(59409) := X"8FC401D8";
        ram_buffer(59410) := X"0C02E477";
        ram_buffer(59411) := X"00000000";
        ram_buffer(59412) := X"10400005";
        ram_buffer(59413) := X"00000000";
        ram_buffer(59414) := X"16900013";
        ram_buffer(59415) := X"00000000";
        ram_buffer(59416) := X"100002B3";
        ram_buffer(59417) := X"00000000";
        ram_buffer(59418) := X"8E220000";
        ram_buffer(59419) := X"00000000";
        ram_buffer(59420) := X"90420000";
        ram_buffer(59421) := X"00000000";
        ram_buffer(59422) := X"00401821";
        ram_buffer(59423) := X"27C20018";
        ram_buffer(59424) := X"00431021";
        ram_buffer(59425) := X"8042005C";
        ram_buffer(59426) := X"00000000";
        ram_buffer(59427) := X"1440FFD6";
        ram_buffer(59428) := X"00000000";
        ram_buffer(59429) := X"10000005";
        ram_buffer(59430) := X"00000000";
        ram_buffer(59431) := X"00000000";
        ram_buffer(59432) := X"10000002";
        ram_buffer(59433) := X"00000000";
        ram_buffer(59434) := X"00000000";
        ram_buffer(59435) := X"02801821";
        ram_buffer(59436) := X"02001021";
        ram_buffer(59437) := X"00629823";
        ram_buffer(59438) := X"126002B3";
        ram_buffer(59439) := X"00000000";
        ram_buffer(59440) := X"A2800000";
        ram_buffer(59441) := X"8FC20018";
        ram_buffer(59442) := X"00000000";
        ram_buffer(59443) := X"24420001";
        ram_buffer(59444) := X"AFC20018";
        ram_buffer(59445) := X"8FC2001C";
        ram_buffer(59446) := X"00000000";
        ram_buffer(59447) := X"00531021";
        ram_buffer(59448) := X"AFC2001C";
        ram_buffer(59449) := X"1000027A";
        ram_buffer(59450) := X"00000000";
        ram_buffer(59451) := X"16400002";
        ram_buffer(59452) := X"00000000";
        ram_buffer(59453) := X"2412FFFF";
        ram_buffer(59454) := X"32020001";
        ram_buffer(59455) := X"1040009C";
        ram_buffer(59456) := X"00000000";
        ram_buffer(59457) := X"27C201A4";
        ram_buffer(59458) := X"24060008";
        ram_buffer(59459) := X"00002821";
        ram_buffer(59460) := X"00402021";
        ram_buffer(59461) := X"0C02801D";
        ram_buffer(59462) := X"00000000";
        ram_buffer(59463) := X"32020010";
        ram_buffer(59464) := X"1440000A";
        ram_buffer(59465) := X"00000000";
        ram_buffer(59466) := X"8FC201E4";
        ram_buffer(59467) := X"00000000";
        ram_buffer(59468) := X"24430004";
        ram_buffer(59469) := X"AFC301E4";
        ram_buffer(59470) := X"8C420000";
        ram_buffer(59471) := X"00000000";
        ram_buffer(59472) := X"AFC20024";
        ram_buffer(59473) := X"10000003";
        ram_buffer(59474) := X"00000000";
        ram_buffer(59475) := X"27C20070";
        ram_buffer(59476) := X"AFC20024";
        ram_buffer(59477) := X"00009821";
        ram_buffer(59478) := X"10000067";
        ram_buffer(59479) := X"00000000";
        ram_buffer(59480) := X"0C02BB09";
        ram_buffer(59481) := X"00000000";
        ram_buffer(59482) := X"1053026D";
        ram_buffer(59483) := X"00000000";
        ram_buffer(59484) := X"02601021";
        ram_buffer(59485) := X"24530001";
        ram_buffer(59486) := X"8E230000";
        ram_buffer(59487) := X"00000000";
        ram_buffer(59488) := X"90630000";
        ram_buffer(59489) := X"00000000";
        ram_buffer(59490) := X"00031E00";
        ram_buffer(59491) := X"00031E03";
        ram_buffer(59492) := X"27C40018";
        ram_buffer(59493) := X"00821021";
        ram_buffer(59494) := X"A043015C";
        ram_buffer(59495) := X"8E220004";
        ram_buffer(59496) := X"00000000";
        ram_buffer(59497) := X"2442FFFF";
        ram_buffer(59498) := X"AE220004";
        ram_buffer(59499) := X"8E220000";
        ram_buffer(59500) := X"00000000";
        ram_buffer(59501) := X"24420001";
        ram_buffer(59502) := X"AE220000";
        ram_buffer(59503) := X"02602021";
        ram_buffer(59504) := X"27C30174";
        ram_buffer(59505) := X"27C201A4";
        ram_buffer(59506) := X"AFA20010";
        ram_buffer(59507) := X"00803821";
        ram_buffer(59508) := X"00603021";
        ram_buffer(59509) := X"8FC50024";
        ram_buffer(59510) := X"8FC401D8";
        ram_buffer(59511) := X"0C02BB73";
        ram_buffer(59512) := X"00000000";
        ram_buffer(59513) := X"AFC20060";
        ram_buffer(59514) := X"8FC30060";
        ram_buffer(59515) := X"2402FFFF";
        ram_buffer(59516) := X"1062024E";
        ram_buffer(59517) := X"00000000";
        ram_buffer(59518) := X"8FC20060";
        ram_buffer(59519) := X"00000000";
        ram_buffer(59520) := X"14400004";
        ram_buffer(59521) := X"00000000";
        ram_buffer(59522) := X"8FC20024";
        ram_buffer(59523) := X"00000000";
        ram_buffer(59524) := X"AC400000";
        ram_buffer(59525) := X"8FC30060";
        ram_buffer(59526) := X"2402FFFE";
        ram_buffer(59527) := X"10620028";
        ram_buffer(59528) := X"00000000";
        ram_buffer(59529) := X"8FC20024";
        ram_buffer(59530) := X"00000000";
        ram_buffer(59531) := X"8C420000";
        ram_buffer(59532) := X"00000000";
        ram_buffer(59533) := X"00402021";
        ram_buffer(59534) := X"0C02BABA";
        ram_buffer(59535) := X"00000000";
        ram_buffer(59536) := X"10400012";
        ram_buffer(59537) := X"00000000";
        ram_buffer(59538) := X"1000000C";
        ram_buffer(59539) := X"00000000";
        ram_buffer(59540) := X"2673FFFF";
        ram_buffer(59541) := X"27C20018";
        ram_buffer(59542) := X"00531021";
        ram_buffer(59543) := X"8042015C";
        ram_buffer(59544) := X"00000000";
        ram_buffer(59545) := X"304200FF";
        ram_buffer(59546) := X"02203021";
        ram_buffer(59547) := X"00402821";
        ram_buffer(59548) := X"8FC401D8";
        ram_buffer(59549) := X"0C02E402";
        ram_buffer(59550) := X"00000000";
        ram_buffer(59551) := X"1660FFF4";
        ram_buffer(59552) := X"00000000";
        ram_buffer(59553) := X"1000002E";
        ram_buffer(59554) := X"00000000";
        ram_buffer(59555) := X"8FC2001C";
        ram_buffer(59556) := X"00000000";
        ram_buffer(59557) := X"00531021";
        ram_buffer(59558) := X"AFC2001C";
        ram_buffer(59559) := X"2652FFFF";
        ram_buffer(59560) := X"32020010";
        ram_buffer(59561) := X"14400005";
        ram_buffer(59562) := X"00000000";
        ram_buffer(59563) := X"8FC20024";
        ram_buffer(59564) := X"00000000";
        ram_buffer(59565) := X"24420004";
        ram_buffer(59566) := X"AFC20024";
        ram_buffer(59567) := X"00009821";
        ram_buffer(59568) := X"8E220004";
        ram_buffer(59569) := X"00000000";
        ram_buffer(59570) := X"1C40000B";
        ram_buffer(59571) := X"00000000";
        ram_buffer(59572) := X"02202821";
        ram_buffer(59573) := X"8FC401D8";
        ram_buffer(59574) := X"0C02E477";
        ram_buffer(59575) := X"00000000";
        ram_buffer(59576) := X"10400005";
        ram_buffer(59577) := X"00000000";
        ram_buffer(59578) := X"12600014";
        ram_buffer(59579) := X"00000000";
        ram_buffer(59580) := X"1000020F";
        ram_buffer(59581) := X"00000000";
        ram_buffer(59582) := X"8F838090";
        ram_buffer(59583) := X"8E220000";
        ram_buffer(59584) := X"00000000";
        ram_buffer(59585) := X"90420000";
        ram_buffer(59586) := X"00000000";
        ram_buffer(59587) := X"24420001";
        ram_buffer(59588) := X"00621021";
        ram_buffer(59589) := X"80420000";
        ram_buffer(59590) := X"00000000";
        ram_buffer(59591) := X"304200FF";
        ram_buffer(59592) := X"30420008";
        ram_buffer(59593) := X"14400006";
        ram_buffer(59594) := X"00000000";
        ram_buffer(59595) := X"1640FF8C";
        ram_buffer(59596) := X"00000000";
        ram_buffer(59597) := X"10000002";
        ram_buffer(59598) := X"00000000";
        ram_buffer(59599) := X"00000000";
        ram_buffer(59600) := X"32020010";
        ram_buffer(59601) := X"144001E1";
        ram_buffer(59602) := X"00000000";
        ram_buffer(59603) := X"8FC20024";
        ram_buffer(59604) := X"00000000";
        ram_buffer(59605) := X"AC400000";
        ram_buffer(59606) := X"8FC20018";
        ram_buffer(59607) := X"00000000";
        ram_buffer(59608) := X"24420001";
        ram_buffer(59609) := X"AFC20018";
        ram_buffer(59610) := X"100001D8";
        ram_buffer(59611) := X"00000000";
        ram_buffer(59612) := X"32020010";
        ram_buffer(59613) := X"10400033";
        ram_buffer(59614) := X"00000000";
        ram_buffer(59615) := X"00009821";
        ram_buffer(59616) := X"10000017";
        ram_buffer(59617) := X"00000000";
        ram_buffer(59618) := X"26730001";
        ram_buffer(59619) := X"8E220004";
        ram_buffer(59620) := X"00000000";
        ram_buffer(59621) := X"2442FFFF";
        ram_buffer(59622) := X"AE220004";
        ram_buffer(59623) := X"8E220000";
        ram_buffer(59624) := X"00000000";
        ram_buffer(59625) := X"24420001";
        ram_buffer(59626) := X"AE220000";
        ram_buffer(59627) := X"2652FFFF";
        ram_buffer(59628) := X"1240001A";
        ram_buffer(59629) := X"00000000";
        ram_buffer(59630) := X"8E220004";
        ram_buffer(59631) := X"00000000";
        ram_buffer(59632) := X"1C400007";
        ram_buffer(59633) := X"00000000";
        ram_buffer(59634) := X"02202821";
        ram_buffer(59635) := X"8FC401D8";
        ram_buffer(59636) := X"0C02E477";
        ram_buffer(59637) := X"00000000";
        ram_buffer(59638) := X"14400013";
        ram_buffer(59639) := X"00000000";
        ram_buffer(59640) := X"8F838090";
        ram_buffer(59641) := X"8E220000";
        ram_buffer(59642) := X"00000000";
        ram_buffer(59643) := X"90420000";
        ram_buffer(59644) := X"00000000";
        ram_buffer(59645) := X"24420001";
        ram_buffer(59646) := X"00621021";
        ram_buffer(59647) := X"80420000";
        ram_buffer(59648) := X"00000000";
        ram_buffer(59649) := X"304200FF";
        ram_buffer(59650) := X"30420008";
        ram_buffer(59651) := X"1040FFDE";
        ram_buffer(59652) := X"00000000";
        ram_buffer(59653) := X"10000005";
        ram_buffer(59654) := X"00000000";
        ram_buffer(59655) := X"00000000";
        ram_buffer(59656) := X"10000002";
        ram_buffer(59657) := X"00000000";
        ram_buffer(59658) := X"00000000";
        ram_buffer(59659) := X"8FC2001C";
        ram_buffer(59660) := X"00000000";
        ram_buffer(59661) := X"00531021";
        ram_buffer(59662) := X"AFC2001C";
        ram_buffer(59663) := X"100001A3";
        ram_buffer(59664) := X"00000000";
        ram_buffer(59665) := X"8FC201E4";
        ram_buffer(59666) := X"00000000";
        ram_buffer(59667) := X"24430004";
        ram_buffer(59668) := X"AFC301E4";
        ram_buffer(59669) := X"8C540000";
        ram_buffer(59670) := X"00000000";
        ram_buffer(59671) := X"02808021";
        ram_buffer(59672) := X"1000001D";
        ram_buffer(59673) := X"00000000";
        ram_buffer(59674) := X"8E220004";
        ram_buffer(59675) := X"00000000";
        ram_buffer(59676) := X"2442FFFF";
        ram_buffer(59677) := X"AE220004";
        ram_buffer(59678) := X"02801821";
        ram_buffer(59679) := X"24740001";
        ram_buffer(59680) := X"8E220000";
        ram_buffer(59681) := X"00000000";
        ram_buffer(59682) := X"24440001";
        ram_buffer(59683) := X"AE240000";
        ram_buffer(59684) := X"90420000";
        ram_buffer(59685) := X"00000000";
        ram_buffer(59686) := X"00021600";
        ram_buffer(59687) := X"00021603";
        ram_buffer(59688) := X"A0620000";
        ram_buffer(59689) := X"2652FFFF";
        ram_buffer(59690) := X"1240001A";
        ram_buffer(59691) := X"00000000";
        ram_buffer(59692) := X"8E220004";
        ram_buffer(59693) := X"00000000";
        ram_buffer(59694) := X"1C400007";
        ram_buffer(59695) := X"00000000";
        ram_buffer(59696) := X"02202821";
        ram_buffer(59697) := X"8FC401D8";
        ram_buffer(59698) := X"0C02E477";
        ram_buffer(59699) := X"00000000";
        ram_buffer(59700) := X"14400013";
        ram_buffer(59701) := X"00000000";
        ram_buffer(59702) := X"8F838090";
        ram_buffer(59703) := X"8E220000";
        ram_buffer(59704) := X"00000000";
        ram_buffer(59705) := X"90420000";
        ram_buffer(59706) := X"00000000";
        ram_buffer(59707) := X"24420001";
        ram_buffer(59708) := X"00621021";
        ram_buffer(59709) := X"80420000";
        ram_buffer(59710) := X"00000000";
        ram_buffer(59711) := X"304200FF";
        ram_buffer(59712) := X"30420008";
        ram_buffer(59713) := X"1040FFD8";
        ram_buffer(59714) := X"00000000";
        ram_buffer(59715) := X"10000005";
        ram_buffer(59716) := X"00000000";
        ram_buffer(59717) := X"00000000";
        ram_buffer(59718) := X"10000002";
        ram_buffer(59719) := X"00000000";
        ram_buffer(59720) := X"00000000";
        ram_buffer(59721) := X"A2800000";
        ram_buffer(59722) := X"02801821";
        ram_buffer(59723) := X"02001021";
        ram_buffer(59724) := X"00621023";
        ram_buffer(59725) := X"8FC3001C";
        ram_buffer(59726) := X"00000000";
        ram_buffer(59727) := X"00621021";
        ram_buffer(59728) := X"AFC2001C";
        ram_buffer(59729) := X"8FC20018";
        ram_buffer(59730) := X"00000000";
        ram_buffer(59731) := X"24420001";
        ram_buffer(59732) := X"AFC20018";
        ram_buffer(59733) := X"1000015D";
        ram_buffer(59734) := X"00000000";
        ram_buffer(59735) := X"AFC00034";
        ram_buffer(59736) := X"AFC00038";
        ram_buffer(59737) := X"2642FFFF";
        ram_buffer(59738) := X"2C420027";
        ram_buffer(59739) := X"14400004";
        ram_buffer(59740) := X"00000000";
        ram_buffer(59741) := X"2642FFD9";
        ram_buffer(59742) := X"AFC20034";
        ram_buffer(59743) := X"24120027";
        ram_buffer(59744) := X"36100D80";
        ram_buffer(59745) := X"27D40174";
        ram_buffer(59746) := X"10000095";
        ram_buffer(59747) := X"00000000";
        ram_buffer(59748) := X"8E220000";
        ram_buffer(59749) := X"00000000";
        ram_buffer(59750) := X"90420000";
        ram_buffer(59751) := X"00000000";
        ram_buffer(59752) := X"00409821";
        ram_buffer(59753) := X"2662FFD5";
        ram_buffer(59754) := X"2C43004E";
        ram_buffer(59755) := X"10600090";
        ram_buffer(59756) := X"00000000";
        ram_buffer(59757) := X"00021880";
        ram_buffer(59758) := X"3C02100D";
        ram_buffer(59759) := X"2442AF5C";
        ram_buffer(59760) := X"00621021";
        ram_buffer(59761) := X"8C420000";
        ram_buffer(59762) := X"00000000";
        ram_buffer(59763) := X"00400008";
        ram_buffer(59764) := X"00000000";
        ram_buffer(59765) := X"32020800";
        ram_buffer(59766) := X"10400066";
        ram_buffer(59767) := X"00000000";
        ram_buffer(59768) := X"8FC20020";
        ram_buffer(59769) := X"00000000";
        ram_buffer(59770) := X"14400004";
        ram_buffer(59771) := X"00000000";
        ram_buffer(59772) := X"24020008";
        ram_buffer(59773) := X"AFC20020";
        ram_buffer(59774) := X"36100200";
        ram_buffer(59775) := X"32020400";
        ram_buffer(59776) := X"10400005";
        ram_buffer(59777) := X"00000000";
        ram_buffer(59778) := X"2402FA7F";
        ram_buffer(59779) := X"02028024";
        ram_buffer(59780) := X"10000059";
        ram_buffer(59781) := X"00000000";
        ram_buffer(59782) := X"2402FC7F";
        ram_buffer(59783) := X"02028024";
        ram_buffer(59784) := X"8FC20034";
        ram_buffer(59785) := X"00000000";
        ram_buffer(59786) := X"10400006";
        ram_buffer(59787) := X"00000000";
        ram_buffer(59788) := X"8FC20034";
        ram_buffer(59789) := X"00000000";
        ram_buffer(59790) := X"2442FFFF";
        ram_buffer(59791) := X"AFC20034";
        ram_buffer(59792) := X"26520001";
        ram_buffer(59793) := X"8FC20038";
        ram_buffer(59794) := X"00000000";
        ram_buffer(59795) := X"24420001";
        ram_buffer(59796) := X"AFC20038";
        ram_buffer(59797) := X"1000004D";
        ram_buffer(59798) := X"00000000";
        ram_buffer(59799) := X"3C02100D";
        ram_buffer(59800) := X"8FC30020";
        ram_buffer(59801) := X"00000000";
        ram_buffer(59802) := X"00031840";
        ram_buffer(59803) := X"2442B094";
        ram_buffer(59804) := X"00621021";
        ram_buffer(59805) := X"84420000";
        ram_buffer(59806) := X"00000000";
        ram_buffer(59807) := X"AFC20020";
        ram_buffer(59808) := X"2402F47F";
        ram_buffer(59809) := X"02028024";
        ram_buffer(59810) := X"1000003B";
        ram_buffer(59811) := X"00000000";
        ram_buffer(59812) := X"3C02100D";
        ram_buffer(59813) := X"8FC30020";
        ram_buffer(59814) := X"00000000";
        ram_buffer(59815) := X"00031840";
        ram_buffer(59816) := X"2442B094";
        ram_buffer(59817) := X"00621021";
        ram_buffer(59818) := X"84420000";
        ram_buffer(59819) := X"00000000";
        ram_buffer(59820) := X"AFC20020";
        ram_buffer(59821) := X"8FC20020";
        ram_buffer(59822) := X"00000000";
        ram_buffer(59823) := X"28420009";
        ram_buffer(59824) := X"14400020";
        ram_buffer(59825) := X"00000000";
        ram_buffer(59826) := X"2402F47F";
        ram_buffer(59827) := X"02028024";
        ram_buffer(59828) := X"10000029";
        ram_buffer(59829) := X"00000000";
        ram_buffer(59830) := X"8FC20020";
        ram_buffer(59831) := X"00000000";
        ram_buffer(59832) := X"2842000B";
        ram_buffer(59833) := X"1440001A";
        ram_buffer(59834) := X"00000000";
        ram_buffer(59835) := X"2402F47F";
        ram_buffer(59836) := X"02028024";
        ram_buffer(59837) := X"10000020";
        ram_buffer(59838) := X"00000000";
        ram_buffer(59839) := X"32020080";
        ram_buffer(59840) := X"10400016";
        ram_buffer(59841) := X"00000000";
        ram_buffer(59842) := X"2402FF7F";
        ram_buffer(59843) := X"02028024";
        ram_buffer(59844) := X"10000019";
        ram_buffer(59845) := X"00000000";
        ram_buffer(59846) := X"32030600";
        ram_buffer(59847) := X"24020200";
        ram_buffer(59848) := X"14620011";
        ram_buffer(59849) := X"00000000";
        ram_buffer(59850) := X"24020010";
        ram_buffer(59851) := X"AFC20020";
        ram_buffer(59852) := X"2402FDFF";
        ram_buffer(59853) := X"02028024";
        ram_buffer(59854) := X"36100500";
        ram_buffer(59855) := X"1000000E";
        ram_buffer(59856) := X"00000000";
        ram_buffer(59857) := X"00000000";
        ram_buffer(59858) := X"10000029";
        ram_buffer(59859) := X"00000000";
        ram_buffer(59860) := X"00000000";
        ram_buffer(59861) := X"10000026";
        ram_buffer(59862) := X"00000000";
        ram_buffer(59863) := X"00000000";
        ram_buffer(59864) := X"10000023";
        ram_buffer(59865) := X"00000000";
        ram_buffer(59866) := X"00000000";
        ram_buffer(59867) := X"10000020";
        ram_buffer(59868) := X"00000000";
        ram_buffer(59869) := X"00000000";
        ram_buffer(59870) := X"02801021";
        ram_buffer(59871) := X"24540001";
        ram_buffer(59872) := X"00131E00";
        ram_buffer(59873) := X"00031E03";
        ram_buffer(59874) := X"A0430000";
        ram_buffer(59875) := X"8E220004";
        ram_buffer(59876) := X"00000000";
        ram_buffer(59877) := X"2442FFFF";
        ram_buffer(59878) := X"AE220004";
        ram_buffer(59879) := X"8E220004";
        ram_buffer(59880) := X"00000000";
        ram_buffer(59881) := X"18400007";
        ram_buffer(59882) := X"00000000";
        ram_buffer(59883) := X"8E220000";
        ram_buffer(59884) := X"00000000";
        ram_buffer(59885) := X"24420001";
        ram_buffer(59886) := X"AE220000";
        ram_buffer(59887) := X"10000007";
        ram_buffer(59888) := X"00000000";
        ram_buffer(59889) := X"02202821";
        ram_buffer(59890) := X"8FC401D8";
        ram_buffer(59891) := X"0C02E477";
        ram_buffer(59892) := X"00000000";
        ram_buffer(59893) := X"14400009";
        ram_buffer(59894) := X"00000000";
        ram_buffer(59895) := X"2652FFFF";
        ram_buffer(59896) := X"1640FF6B";
        ram_buffer(59897) := X"00000000";
        ram_buffer(59898) := X"10000005";
        ram_buffer(59899) := X"00000000";
        ram_buffer(59900) := X"00000000";
        ram_buffer(59901) := X"10000002";
        ram_buffer(59902) := X"00000000";
        ram_buffer(59903) := X"00000000";
        ram_buffer(59904) := X"32020100";
        ram_buffer(59905) := X"1040000F";
        ram_buffer(59906) := X"00000000";
        ram_buffer(59907) := X"27C20174";
        ram_buffer(59908) := X"0054102B";
        ram_buffer(59909) := X"10400008";
        ram_buffer(59910) := X"00000000";
        ram_buffer(59911) := X"2694FFFF";
        ram_buffer(59912) := X"82820000";
        ram_buffer(59913) := X"02203021";
        ram_buffer(59914) := X"00402821";
        ram_buffer(59915) := X"8FC401D8";
        ram_buffer(59916) := X"0C02E402";
        ram_buffer(59917) := X"00000000";
        ram_buffer(59918) := X"27C20174";
        ram_buffer(59919) := X"128200D5";
        ram_buffer(59920) := X"00000000";
        ram_buffer(59921) := X"32020010";
        ram_buffer(59922) := X"1440008B";
        ram_buffer(59923) := X"00000000";
        ram_buffer(59924) := X"A2800000";
        ram_buffer(59925) := X"27C30174";
        ram_buffer(59926) := X"8FC20028";
        ram_buffer(59927) := X"8FC70020";
        ram_buffer(59928) := X"00003021";
        ram_buffer(59929) := X"00602821";
        ram_buffer(59930) := X"8FC401D8";
        ram_buffer(59931) := X"0040F809";
        ram_buffer(59932) := X"00000000";
        ram_buffer(59933) := X"AFC20068";
        ram_buffer(59934) := X"32020020";
        ram_buffer(59935) := X"1040000E";
        ram_buffer(59936) := X"00000000";
        ram_buffer(59937) := X"8FC201E4";
        ram_buffer(59938) := X"00000000";
        ram_buffer(59939) := X"24430004";
        ram_buffer(59940) := X"AFC301E4";
        ram_buffer(59941) := X"8C420000";
        ram_buffer(59942) := X"00000000";
        ram_buffer(59943) := X"AFC2006C";
        ram_buffer(59944) := X"8FC30068";
        ram_buffer(59945) := X"8FC2006C";
        ram_buffer(59946) := X"00000000";
        ram_buffer(59947) := X"AC430000";
        ram_buffer(59948) := X"1000006D";
        ram_buffer(59949) := X"00000000";
        ram_buffer(59950) := X"32020008";
        ram_buffer(59951) := X"10400011";
        ram_buffer(59952) := X"00000000";
        ram_buffer(59953) := X"8FC201E4";
        ram_buffer(59954) := X"00000000";
        ram_buffer(59955) := X"24430004";
        ram_buffer(59956) := X"AFC301E4";
        ram_buffer(59957) := X"8C420000";
        ram_buffer(59958) := X"00000000";
        ram_buffer(59959) := X"AFC2004C";
        ram_buffer(59960) := X"8FC20068";
        ram_buffer(59961) := X"00000000";
        ram_buffer(59962) := X"00021E00";
        ram_buffer(59963) := X"00031E03";
        ram_buffer(59964) := X"8FC2004C";
        ram_buffer(59965) := X"00000000";
        ram_buffer(59966) := X"A0430000";
        ram_buffer(59967) := X"1000005A";
        ram_buffer(59968) := X"00000000";
        ram_buffer(59969) := X"32020004";
        ram_buffer(59970) := X"10400011";
        ram_buffer(59971) := X"00000000";
        ram_buffer(59972) := X"8FC201E4";
        ram_buffer(59973) := X"00000000";
        ram_buffer(59974) := X"24430004";
        ram_buffer(59975) := X"AFC301E4";
        ram_buffer(59976) := X"8C420000";
        ram_buffer(59977) := X"00000000";
        ram_buffer(59978) := X"AFC20050";
        ram_buffer(59979) := X"8FC20068";
        ram_buffer(59980) := X"00000000";
        ram_buffer(59981) := X"00021C00";
        ram_buffer(59982) := X"00031C03";
        ram_buffer(59983) := X"8FC20050";
        ram_buffer(59984) := X"00000000";
        ram_buffer(59985) := X"A4430000";
        ram_buffer(59986) := X"10000047";
        ram_buffer(59987) := X"00000000";
        ram_buffer(59988) := X"32020001";
        ram_buffer(59989) := X"1040000E";
        ram_buffer(59990) := X"00000000";
        ram_buffer(59991) := X"8FC201E4";
        ram_buffer(59992) := X"00000000";
        ram_buffer(59993) := X"24430004";
        ram_buffer(59994) := X"AFC301E4";
        ram_buffer(59995) := X"8C420000";
        ram_buffer(59996) := X"00000000";
        ram_buffer(59997) := X"AFC20054";
        ram_buffer(59998) := X"8FC30068";
        ram_buffer(59999) := X"8FC20054";
        ram_buffer(60000) := X"00000000";
        ram_buffer(60001) := X"AC430000";
        ram_buffer(60002) := X"10000037";
        ram_buffer(60003) := X"00000000";
        ram_buffer(60004) := X"32020002";
        ram_buffer(60005) := X"10400029";
        ram_buffer(60006) := X"00000000";
        ram_buffer(60007) := X"8FC30028";
        ram_buffer(60008) := X"3C02100B";
        ram_buffer(60009) := X"24426A64";
        ram_buffer(60010) := X"1462000C";
        ram_buffer(60011) := X"00000000";
        ram_buffer(60012) := X"27C20174";
        ram_buffer(60013) := X"8FC70020";
        ram_buffer(60014) := X"00003021";
        ram_buffer(60015) := X"00402821";
        ram_buffer(60016) := X"8FC401D8";
        ram_buffer(60017) := X"0C02DB85";
        ram_buffer(60018) := X"00000000";
        ram_buffer(60019) := X"AFC30044";
        ram_buffer(60020) := X"AFC20040";
        ram_buffer(60021) := X"1000000A";
        ram_buffer(60022) := X"00000000";
        ram_buffer(60023) := X"27C20174";
        ram_buffer(60024) := X"8FC70020";
        ram_buffer(60025) := X"00003021";
        ram_buffer(60026) := X"00402821";
        ram_buffer(60027) := X"8FC401D8";
        ram_buffer(60028) := X"0C02D961";
        ram_buffer(60029) := X"00000000";
        ram_buffer(60030) := X"AFC30044";
        ram_buffer(60031) := X"AFC20040";
        ram_buffer(60032) := X"8FC201E4";
        ram_buffer(60033) := X"00000000";
        ram_buffer(60034) := X"24430004";
        ram_buffer(60035) := X"AFC301E4";
        ram_buffer(60036) := X"8C420000";
        ram_buffer(60037) := X"00000000";
        ram_buffer(60038) := X"AFC20058";
        ram_buffer(60039) := X"8FC30044";
        ram_buffer(60040) := X"8FC20040";
        ram_buffer(60041) := X"8FC40058";
        ram_buffer(60042) := X"00000000";
        ram_buffer(60043) := X"AC830004";
        ram_buffer(60044) := X"AC820000";
        ram_buffer(60045) := X"1000000C";
        ram_buffer(60046) := X"00000000";
        ram_buffer(60047) := X"8FC201E4";
        ram_buffer(60048) := X"00000000";
        ram_buffer(60049) := X"24430004";
        ram_buffer(60050) := X"AFC301E4";
        ram_buffer(60051) := X"8C420000";
        ram_buffer(60052) := X"00000000";
        ram_buffer(60053) := X"AFC2005C";
        ram_buffer(60054) := X"8FC30068";
        ram_buffer(60055) := X"8FC2005C";
        ram_buffer(60056) := X"00000000";
        ram_buffer(60057) := X"AC430000";
        ram_buffer(60058) := X"8FC20018";
        ram_buffer(60059) := X"00000000";
        ram_buffer(60060) := X"24420001";
        ram_buffer(60061) := X"AFC20018";
        ram_buffer(60062) := X"02801821";
        ram_buffer(60063) := X"27C20174";
        ram_buffer(60064) := X"00621823";
        ram_buffer(60065) := X"8FC20038";
        ram_buffer(60066) := X"00000000";
        ram_buffer(60067) := X"00621021";
        ram_buffer(60068) := X"8FC3001C";
        ram_buffer(60069) := X"00000000";
        ram_buffer(60070) := X"00621021";
        ram_buffer(60071) := X"AFC2001C";
        ram_buffer(60072) := X"1000000B";
        ram_buffer(60073) := X"00000000";
        ram_buffer(60074) := X"00000000";
        ram_buffer(60075) := X"1000FA95";
        ram_buffer(60076) := X"00000000";
        ram_buffer(60077) := X"00000000";
        ram_buffer(60078) := X"1000FA92";
        ram_buffer(60079) := X"00000000";
        ram_buffer(60080) := X"00000000";
        ram_buffer(60081) := X"1000FA8F";
        ram_buffer(60082) := X"00000000";
        ram_buffer(60083) := X"00000000";
        ram_buffer(60084) := X"1000FA8C";
        ram_buffer(60085) := X"00000000";
        ram_buffer(60086) := X"00000000";
        ram_buffer(60087) := X"10000014";
        ram_buffer(60088) := X"00000000";
        ram_buffer(60089) := X"00000000";
        ram_buffer(60090) := X"10000011";
        ram_buffer(60091) := X"00000000";
        ram_buffer(60092) := X"00000000";
        ram_buffer(60093) := X"1000000E";
        ram_buffer(60094) := X"00000000";
        ram_buffer(60095) := X"00000000";
        ram_buffer(60096) := X"1000000B";
        ram_buffer(60097) := X"00000000";
        ram_buffer(60098) := X"00000000";
        ram_buffer(60099) := X"10000008";
        ram_buffer(60100) := X"00000000";
        ram_buffer(60101) := X"00000000";
        ram_buffer(60102) := X"10000005";
        ram_buffer(60103) := X"00000000";
        ram_buffer(60104) := X"00000000";
        ram_buffer(60105) := X"10000002";
        ram_buffer(60106) := X"00000000";
        ram_buffer(60107) := X"00000000";
        ram_buffer(60108) := X"8FC20018";
        ram_buffer(60109) := X"00000000";
        ram_buffer(60110) := X"1040000A";
        ram_buffer(60111) := X"00000000";
        ram_buffer(60112) := X"8622000C";
        ram_buffer(60113) := X"00000000";
        ram_buffer(60114) := X"3042FFFF";
        ram_buffer(60115) := X"30420040";
        ram_buffer(60116) := X"14400004";
        ram_buffer(60117) := X"00000000";
        ram_buffer(60118) := X"8FC20018";
        ram_buffer(60119) := X"1000000F";
        ram_buffer(60120) := X"00000000";
        ram_buffer(60121) := X"2402FFFF";
        ram_buffer(60122) := X"1000000C";
        ram_buffer(60123) := X"00000000";
        ram_buffer(60124) := X"00000000";
        ram_buffer(60125) := X"10000008";
        ram_buffer(60126) := X"00000000";
        ram_buffer(60127) := X"00000000";
        ram_buffer(60128) := X"10000005";
        ram_buffer(60129) := X"00000000";
        ram_buffer(60130) := X"00000000";
        ram_buffer(60131) := X"10000002";
        ram_buffer(60132) := X"00000000";
        ram_buffer(60133) := X"00000000";
        ram_buffer(60134) := X"8FC20018";
        ram_buffer(60135) := X"03C0E821";
        ram_buffer(60136) := X"8FBF01D4";
        ram_buffer(60137) := X"8FBE01D0";
        ram_buffer(60138) := X"8FB701CC";
        ram_buffer(60139) := X"8FB601C8";
        ram_buffer(60140) := X"8FB501C4";
        ram_buffer(60141) := X"8FB401C0";
        ram_buffer(60142) := X"8FB301BC";
        ram_buffer(60143) := X"8FB201B8";
        ram_buffer(60144) := X"8FB101B4";
        ram_buffer(60145) := X"8FB001B0";
        ram_buffer(60146) := X"27BD01D8";
        ram_buffer(60147) := X"03E00008";
        ram_buffer(60148) := X"00000000";
        ram_buffer(60149) := X"27BDFFD0";
        ram_buffer(60150) := X"AFBF002C";
        ram_buffer(60151) := X"AFBE0028";
        ram_buffer(60152) := X"AFB10024";
        ram_buffer(60153) := X"AFB00020";
        ram_buffer(60154) := X"03A0F021";
        ram_buffer(60155) := X"AFC40030";
        ram_buffer(60156) := X"AFC50034";
        ram_buffer(60157) := X"00C08021";
        ram_buffer(60158) := X"00008821";
        ram_buffer(60159) := X"8E020008";
        ram_buffer(60160) := X"00000000";
        ram_buffer(60161) := X"14400005";
        ram_buffer(60162) := X"00000000";
        ram_buffer(60163) := X"AE000004";
        ram_buffer(60164) := X"00001021";
        ram_buffer(60165) := X"10000051";
        ram_buffer(60166) := X"00000000";
        ram_buffer(60167) := X"8FC20034";
        ram_buffer(60168) := X"00000000";
        ram_buffer(60169) := X"8C420064";
        ram_buffer(60170) := X"00000000";
        ram_buffer(60171) := X"30422000";
        ram_buffer(60172) := X"10400041";
        ram_buffer(60173) := X"00000000";
        ram_buffer(60174) := X"8E020000";
        ram_buffer(60175) := X"00000000";
        ram_buffer(60176) := X"AFC20010";
        ram_buffer(60177) := X"10000036";
        ram_buffer(60178) := X"00000000";
        ram_buffer(60179) := X"8FC20010";
        ram_buffer(60180) := X"00000000";
        ram_buffer(60181) := X"8C420000";
        ram_buffer(60182) := X"00000000";
        ram_buffer(60183) := X"AFC20018";
        ram_buffer(60184) := X"8FC20010";
        ram_buffer(60185) := X"00000000";
        ram_buffer(60186) := X"8C420004";
        ram_buffer(60187) := X"00000000";
        ram_buffer(60188) := X"00021082";
        ram_buffer(60189) := X"AFC2001C";
        ram_buffer(60190) := X"AFC00014";
        ram_buffer(60191) := X"10000018";
        ram_buffer(60192) := X"00000000";
        ram_buffer(60193) := X"8FC20014";
        ram_buffer(60194) := X"00000000";
        ram_buffer(60195) := X"00021080";
        ram_buffer(60196) := X"8FC30018";
        ram_buffer(60197) := X"00000000";
        ram_buffer(60198) := X"00621021";
        ram_buffer(60199) := X"8C420000";
        ram_buffer(60200) := X"8FC60034";
        ram_buffer(60201) := X"00402821";
        ram_buffer(60202) := X"8FC40030";
        ram_buffer(60203) := X"0C02F386";
        ram_buffer(60204) := X"00000000";
        ram_buffer(60205) := X"00401821";
        ram_buffer(60206) := X"2402FFFF";
        ram_buffer(60207) := X"14620004";
        ram_buffer(60208) := X"00000000";
        ram_buffer(60209) := X"2411FFFF";
        ram_buffer(60210) := X"10000021";
        ram_buffer(60211) := X"00000000";
        ram_buffer(60212) := X"8FC20014";
        ram_buffer(60213) := X"00000000";
        ram_buffer(60214) := X"24420001";
        ram_buffer(60215) := X"AFC20014";
        ram_buffer(60216) := X"8FC30014";
        ram_buffer(60217) := X"8FC2001C";
        ram_buffer(60218) := X"00000000";
        ram_buffer(60219) := X"0062102A";
        ram_buffer(60220) := X"1440FFE4";
        ram_buffer(60221) := X"00000000";
        ram_buffer(60222) := X"8E030008";
        ram_buffer(60223) := X"8FC2001C";
        ram_buffer(60224) := X"00000000";
        ram_buffer(60225) := X"00021080";
        ram_buffer(60226) := X"00621023";
        ram_buffer(60227) := X"AE020008";
        ram_buffer(60228) := X"8FC20010";
        ram_buffer(60229) := X"00000000";
        ram_buffer(60230) := X"24420008";
        ram_buffer(60231) := X"AFC20010";
        ram_buffer(60232) := X"8E020008";
        ram_buffer(60233) := X"00000000";
        ram_buffer(60234) := X"1440FFC8";
        ram_buffer(60235) := X"00000000";
        ram_buffer(60236) := X"10000007";
        ram_buffer(60237) := X"00000000";
        ram_buffer(60238) := X"02003021";
        ram_buffer(60239) := X"8FC50034";
        ram_buffer(60240) := X"8FC40030";
        ram_buffer(60241) := X"0C02B89A";
        ram_buffer(60242) := X"00000000";
        ram_buffer(60243) := X"00408821";
        ram_buffer(60244) := X"AE000008";
        ram_buffer(60245) := X"AE000004";
        ram_buffer(60246) := X"02201021";
        ram_buffer(60247) := X"03C0E821";
        ram_buffer(60248) := X"8FBF002C";
        ram_buffer(60249) := X"8FBE0028";
        ram_buffer(60250) := X"8FB10024";
        ram_buffer(60251) := X"8FB00020";
        ram_buffer(60252) := X"27BD0030";
        ram_buffer(60253) := X"03E00008";
        ram_buffer(60254) := X"00000000";
        ram_buffer(60255) := X"27BDFB70";
        ram_buffer(60256) := X"AFBF048C";
        ram_buffer(60257) := X"AFBE0488";
        ram_buffer(60258) := X"AFB00484";
        ram_buffer(60259) := X"03A0F021";
        ram_buffer(60260) := X"AFC40490";
        ram_buffer(60261) := X"00A08021";
        ram_buffer(60262) := X"AFC60498";
        ram_buffer(60263) := X"AFC7049C";
        ram_buffer(60264) := X"8603000C";
        ram_buffer(60265) := X"2402FFFD";
        ram_buffer(60266) := X"00621024";
        ram_buffer(60267) := X"00021400";
        ram_buffer(60268) := X"00021403";
        ram_buffer(60269) := X"A7C20020";
        ram_buffer(60270) := X"8E020064";
        ram_buffer(60271) := X"00000000";
        ram_buffer(60272) := X"AFC20078";
        ram_buffer(60273) := X"8602000E";
        ram_buffer(60274) := X"00000000";
        ram_buffer(60275) := X"A7C20022";
        ram_buffer(60276) := X"8E02001C";
        ram_buffer(60277) := X"00000000";
        ram_buffer(60278) := X"AFC20030";
        ram_buffer(60279) := X"8E020024";
        ram_buffer(60280) := X"00000000";
        ram_buffer(60281) := X"AFC20038";
        ram_buffer(60282) := X"27C2007C";
        ram_buffer(60283) := X"AFC20014";
        ram_buffer(60284) := X"8FC20014";
        ram_buffer(60285) := X"00000000";
        ram_buffer(60286) := X"AFC20024";
        ram_buffer(60287) := X"24020400";
        ram_buffer(60288) := X"AFC2001C";
        ram_buffer(60289) := X"8FC2001C";
        ram_buffer(60290) := X"00000000";
        ram_buffer(60291) := X"AFC20028";
        ram_buffer(60292) := X"AFC0002C";
        ram_buffer(60293) := X"27C20014";
        ram_buffer(60294) := X"8FC7049C";
        ram_buffer(60295) := X"8FC60498";
        ram_buffer(60296) := X"00402821";
        ram_buffer(60297) := X"8FC40490";
        ram_buffer(60298) := X"0C02EBC4";
        ram_buffer(60299) := X"00000000";
        ram_buffer(60300) := X"AFC20010";
        ram_buffer(60301) := X"8FC20010";
        ram_buffer(60302) := X"00000000";
        ram_buffer(60303) := X"0440000A";
        ram_buffer(60304) := X"00000000";
        ram_buffer(60305) := X"27C20014";
        ram_buffer(60306) := X"00402821";
        ram_buffer(60307) := X"8FC40490";
        ram_buffer(60308) := X"0C026EE1";
        ram_buffer(60309) := X"00000000";
        ram_buffer(60310) := X"10400003";
        ram_buffer(60311) := X"00000000";
        ram_buffer(60312) := X"2402FFFF";
        ram_buffer(60313) := X"AFC20010";
        ram_buffer(60314) := X"87C20020";
        ram_buffer(60315) := X"00000000";
        ram_buffer(60316) := X"3042FFFF";
        ram_buffer(60317) := X"30420040";
        ram_buffer(60318) := X"10400007";
        ram_buffer(60319) := X"00000000";
        ram_buffer(60320) := X"8602000C";
        ram_buffer(60321) := X"00000000";
        ram_buffer(60322) := X"34420040";
        ram_buffer(60323) := X"00021400";
        ram_buffer(60324) := X"00021403";
        ram_buffer(60325) := X"A602000C";
        ram_buffer(60326) := X"8FC20010";
        ram_buffer(60327) := X"03C0E821";
        ram_buffer(60328) := X"8FBF048C";
        ram_buffer(60329) := X"8FBE0488";
        ram_buffer(60330) := X"8FB00484";
        ram_buffer(60331) := X"27BD0490";
        ram_buffer(60332) := X"03E00008";
        ram_buffer(60333) := X"00000000";
        ram_buffer(60334) := X"27BDFFE0";
        ram_buffer(60335) := X"AFBF001C";
        ram_buffer(60336) := X"AFBE0018";
        ram_buffer(60337) := X"03A0F021";
        ram_buffer(60338) := X"AFC40020";
        ram_buffer(60339) := X"AFC50024";
        ram_buffer(60340) := X"AFC60028";
        ram_buffer(60341) := X"8F828098";
        ram_buffer(60342) := X"8FC70028";
        ram_buffer(60343) := X"8FC60024";
        ram_buffer(60344) := X"8FC50020";
        ram_buffer(60345) := X"00402021";
        ram_buffer(60346) := X"0C02EBC4";
        ram_buffer(60347) := X"00000000";
        ram_buffer(60348) := X"AFC20010";
        ram_buffer(60349) := X"8FC20010";
        ram_buffer(60350) := X"03C0E821";
        ram_buffer(60351) := X"8FBF001C";
        ram_buffer(60352) := X"8FBE0018";
        ram_buffer(60353) := X"27BD0020";
        ram_buffer(60354) := X"03E00008";
        ram_buffer(60355) := X"00000000";
        ram_buffer(60356) := X"27BDFE70";
        ram_buffer(60357) := X"AFBF018C";
        ram_buffer(60358) := X"AFBE0188";
        ram_buffer(60359) := X"AFB70184";
        ram_buffer(60360) := X"AFB60180";
        ram_buffer(60361) := X"AFB5017C";
        ram_buffer(60362) := X"AFB40178";
        ram_buffer(60363) := X"AFB30174";
        ram_buffer(60364) := X"AFB20170";
        ram_buffer(60365) := X"AFB1016C";
        ram_buffer(60366) := X"AFB00168";
        ram_buffer(60367) := X"03A0F021";
        ram_buffer(60368) := X"AFC40190";
        ram_buffer(60369) := X"AFC50194";
        ram_buffer(60370) := X"AFC60198";
        ram_buffer(60371) := X"AFC7019C";
        ram_buffer(60372) := X"AFC0001C";
        ram_buffer(60373) := X"AFC00020";
        ram_buffer(60374) := X"AFC00024";
        ram_buffer(60375) := X"AFC00028";
        ram_buffer(60376) := X"AFC00048";
        ram_buffer(60377) := X"AFC0004C";
        ram_buffer(60378) := X"8FC20190";
        ram_buffer(60379) := X"00000000";
        ram_buffer(60380) := X"AFC20050";
        ram_buffer(60381) := X"8FC20050";
        ram_buffer(60382) := X"00000000";
        ram_buffer(60383) := X"1040000A";
        ram_buffer(60384) := X"00000000";
        ram_buffer(60385) := X"8FC20050";
        ram_buffer(60386) := X"00000000";
        ram_buffer(60387) := X"8C420038";
        ram_buffer(60388) := X"00000000";
        ram_buffer(60389) := X"14400004";
        ram_buffer(60390) := X"00000000";
        ram_buffer(60391) := X"8FC40050";
        ram_buffer(60392) := X"0C027069";
        ram_buffer(60393) := X"00000000";
        ram_buffer(60394) := X"8FC20194";
        ram_buffer(60395) := X"00000000";
        ram_buffer(60396) := X"8442000C";
        ram_buffer(60397) := X"00000000";
        ram_buffer(60398) := X"3042FFFF";
        ram_buffer(60399) := X"30422000";
        ram_buffer(60400) := X"14400013";
        ram_buffer(60401) := X"00000000";
        ram_buffer(60402) := X"8FC20194";
        ram_buffer(60403) := X"00000000";
        ram_buffer(60404) := X"8442000C";
        ram_buffer(60405) := X"00000000";
        ram_buffer(60406) := X"34422000";
        ram_buffer(60407) := X"00021C00";
        ram_buffer(60408) := X"00031C03";
        ram_buffer(60409) := X"8FC20194";
        ram_buffer(60410) := X"00000000";
        ram_buffer(60411) := X"A443000C";
        ram_buffer(60412) := X"8FC20194";
        ram_buffer(60413) := X"00000000";
        ram_buffer(60414) := X"8C430064";
        ram_buffer(60415) := X"2402DFFF";
        ram_buffer(60416) := X"00621824";
        ram_buffer(60417) := X"8FC20194";
        ram_buffer(60418) := X"00000000";
        ram_buffer(60419) := X"AC430064";
        ram_buffer(60420) := X"8FC20194";
        ram_buffer(60421) := X"00000000";
        ram_buffer(60422) := X"8442000C";
        ram_buffer(60423) := X"00000000";
        ram_buffer(60424) := X"3042FFFF";
        ram_buffer(60425) := X"30420008";
        ram_buffer(60426) := X"10400007";
        ram_buffer(60427) := X"00000000";
        ram_buffer(60428) := X"8FC20194";
        ram_buffer(60429) := X"00000000";
        ram_buffer(60430) := X"8C420010";
        ram_buffer(60431) := X"00000000";
        ram_buffer(60432) := X"1440000A";
        ram_buffer(60433) := X"00000000";
        ram_buffer(60434) := X"8FC50194";
        ram_buffer(60435) := X"8FC40190";
        ram_buffer(60436) := X"0C02ACF1";
        ram_buffer(60437) := X"00000000";
        ram_buffer(60438) := X"10400004";
        ram_buffer(60439) := X"00000000";
        ram_buffer(60440) := X"2402FFFF";
        ram_buffer(60441) := X"10000629";
        ram_buffer(60442) := X"00000000";
        ram_buffer(60443) := X"8FC20194";
        ram_buffer(60444) := X"00000000";
        ram_buffer(60445) := X"8442000C";
        ram_buffer(60446) := X"00000000";
        ram_buffer(60447) := X"3042FFFF";
        ram_buffer(60448) := X"3043001A";
        ram_buffer(60449) := X"2402000A";
        ram_buffer(60450) := X"1462000F";
        ram_buffer(60451) := X"00000000";
        ram_buffer(60452) := X"8FC20194";
        ram_buffer(60453) := X"00000000";
        ram_buffer(60454) := X"8442000E";
        ram_buffer(60455) := X"00000000";
        ram_buffer(60456) := X"04400009";
        ram_buffer(60457) := X"00000000";
        ram_buffer(60458) := X"8FC7019C";
        ram_buffer(60459) := X"8FC60198";
        ram_buffer(60460) := X"8FC50194";
        ram_buffer(60461) := X"8FC40190";
        ram_buffer(60462) := X"0C02EB5F";
        ram_buffer(60463) := X"00000000";
        ram_buffer(60464) := X"10000612";
        ram_buffer(60465) := X"00000000";
        ram_buffer(60466) := X"8FD50198";
        ram_buffer(60467) := X"27D1006C";
        ram_buffer(60468) := X"AFD10060";
        ram_buffer(60469) := X"AFC00068";
        ram_buffer(60470) := X"AFC00064";
        ram_buffer(60471) := X"AFC00010";
        ram_buffer(60472) := X"02A09821";
        ram_buffer(60473) := X"10000002";
        ram_buffer(60474) := X"00000000";
        ram_buffer(60475) := X"26B50001";
        ram_buffer(60476) := X"82A20000";
        ram_buffer(60477) := X"00000000";
        ram_buffer(60478) := X"10400005";
        ram_buffer(60479) := X"00000000";
        ram_buffer(60480) := X"82A30000";
        ram_buffer(60481) := X"24020025";
        ram_buffer(60482) := X"1462FFF8";
        ram_buffer(60483) := X"00000000";
        ram_buffer(60484) := X"02A01821";
        ram_buffer(60485) := X"02601021";
        ram_buffer(60486) := X"00628023";
        ram_buffer(60487) := X"1200001F";
        ram_buffer(60488) := X"00000000";
        ram_buffer(60489) := X"AE330000";
        ram_buffer(60490) := X"02001021";
        ram_buffer(60491) := X"AE220004";
        ram_buffer(60492) := X"8FC20068";
        ram_buffer(60493) := X"02001821";
        ram_buffer(60494) := X"00431021";
        ram_buffer(60495) := X"AFC20068";
        ram_buffer(60496) := X"26310008";
        ram_buffer(60497) := X"8FC20064";
        ram_buffer(60498) := X"00000000";
        ram_buffer(60499) := X"24420001";
        ram_buffer(60500) := X"AFC20064";
        ram_buffer(60501) := X"8FC20064";
        ram_buffer(60502) := X"00000000";
        ram_buffer(60503) := X"28420008";
        ram_buffer(60504) := X"1440000A";
        ram_buffer(60505) := X"00000000";
        ram_buffer(60506) := X"27C20060";
        ram_buffer(60507) := X"00403021";
        ram_buffer(60508) := X"8FC50194";
        ram_buffer(60509) := X"8FC40190";
        ram_buffer(60510) := X"0C02EAF5";
        ram_buffer(60511) := X"00000000";
        ram_buffer(60512) := X"144005A5";
        ram_buffer(60513) := X"00000000";
        ram_buffer(60514) := X"27D1006C";
        ram_buffer(60515) := X"8FC20010";
        ram_buffer(60516) := X"00000000";
        ram_buffer(60517) := X"00501021";
        ram_buffer(60518) := X"AFC20010";
        ram_buffer(60519) := X"82A20000";
        ram_buffer(60520) := X"00000000";
        ram_buffer(60521) := X"10400588";
        ram_buffer(60522) := X"00000000";
        ram_buffer(60523) := X"AFD50054";
        ram_buffer(60524) := X"26B50001";
        ram_buffer(60525) := X"00009021";
        ram_buffer(60526) := X"AFC0003C";
        ram_buffer(60527) := X"AFC00014";
        ram_buffer(60528) := X"2402FFFF";
        ram_buffer(60529) := X"AFC20018";
        ram_buffer(60530) := X"A3C0005C";
        ram_buffer(60531) := X"02A01021";
        ram_buffer(60532) := X"24550001";
        ram_buffer(60533) := X"80420000";
        ram_buffer(60534) := X"00000000";
        ram_buffer(60535) := X"0040A021";
        ram_buffer(60536) := X"2683FFE0";
        ram_buffer(60537) := X"2C62005B";
        ram_buffer(60538) := X"104003BF";
        ram_buffer(60539) := X"00000000";
        ram_buffer(60540) := X"00031880";
        ram_buffer(60541) := X"3C02100D";
        ram_buffer(60542) := X"2442B104";
        ram_buffer(60543) := X"00621021";
        ram_buffer(60544) := X"8C420000";
        ram_buffer(60545) := X"00000000";
        ram_buffer(60546) := X"00400008";
        ram_buffer(60547) := X"00000000";
        ram_buffer(60548) := X"8FC40190";
        ram_buffer(60549) := X"0C02BB25";
        ram_buffer(60550) := X"00000000";
        ram_buffer(60551) := X"8C420004";
        ram_buffer(60552) := X"00000000";
        ram_buffer(60553) := X"AFC2001C";
        ram_buffer(60554) := X"8FC4001C";
        ram_buffer(60555) := X"0C02851E";
        ram_buffer(60556) := X"00000000";
        ram_buffer(60557) := X"AFC20020";
        ram_buffer(60558) := X"8FC40190";
        ram_buffer(60559) := X"0C02BB25";
        ram_buffer(60560) := X"00000000";
        ram_buffer(60561) := X"8C420008";
        ram_buffer(60562) := X"00000000";
        ram_buffer(60563) := X"AFC20024";
        ram_buffer(60564) := X"8FC20020";
        ram_buffer(60565) := X"00000000";
        ram_buffer(60566) := X"1040FFDC";
        ram_buffer(60567) := X"00000000";
        ram_buffer(60568) := X"8FC20024";
        ram_buffer(60569) := X"00000000";
        ram_buffer(60570) := X"1040FFD8";
        ram_buffer(60571) := X"00000000";
        ram_buffer(60572) := X"8FC20024";
        ram_buffer(60573) := X"00000000";
        ram_buffer(60574) := X"80420000";
        ram_buffer(60575) := X"00000000";
        ram_buffer(60576) := X"1040FFD2";
        ram_buffer(60577) := X"00000000";
        ram_buffer(60578) := X"36520400";
        ram_buffer(60579) := X"1000FFCF";
        ram_buffer(60580) := X"00000000";
        ram_buffer(60581) := X"83C2005C";
        ram_buffer(60582) := X"00000000";
        ram_buffer(60583) := X"1440FFCB";
        ram_buffer(60584) := X"00000000";
        ram_buffer(60585) := X"24020020";
        ram_buffer(60586) := X"A3C2005C";
        ram_buffer(60587) := X"1000FFC7";
        ram_buffer(60588) := X"00000000";
        ram_buffer(60589) := X"36520001";
        ram_buffer(60590) := X"1000FFC4";
        ram_buffer(60591) := X"00000000";
        ram_buffer(60592) := X"8FC2019C";
        ram_buffer(60593) := X"00000000";
        ram_buffer(60594) := X"24430004";
        ram_buffer(60595) := X"AFC3019C";
        ram_buffer(60596) := X"8C420000";
        ram_buffer(60597) := X"00000000";
        ram_buffer(60598) := X"AFC20014";
        ram_buffer(60599) := X"8FC20014";
        ram_buffer(60600) := X"00000000";
        ram_buffer(60601) := X"04400003";
        ram_buffer(60602) := X"00000000";
        ram_buffer(60603) := X"1000FFB7";
        ram_buffer(60604) := X"00000000";
        ram_buffer(60605) := X"8FC20014";
        ram_buffer(60606) := X"00000000";
        ram_buffer(60607) := X"00021023";
        ram_buffer(60608) := X"AFC20014";
        ram_buffer(60609) := X"36520004";
        ram_buffer(60610) := X"1000FFB0";
        ram_buffer(60611) := X"00000000";
        ram_buffer(60612) := X"2402002B";
        ram_buffer(60613) := X"A3C2005C";
        ram_buffer(60614) := X"1000FFAC";
        ram_buffer(60615) := X"00000000";
        ram_buffer(60616) := X"02A01021";
        ram_buffer(60617) := X"24550001";
        ram_buffer(60618) := X"80420000";
        ram_buffer(60619) := X"00000000";
        ram_buffer(60620) := X"0040A021";
        ram_buffer(60621) := X"2402002A";
        ram_buffer(60622) := X"16820010";
        ram_buffer(60623) := X"00000000";
        ram_buffer(60624) := X"8FC2019C";
        ram_buffer(60625) := X"00000000";
        ram_buffer(60626) := X"24430004";
        ram_buffer(60627) := X"AFC3019C";
        ram_buffer(60628) := X"8C420000";
        ram_buffer(60629) := X"00000000";
        ram_buffer(60630) := X"AFC20018";
        ram_buffer(60631) := X"8FC20018";
        ram_buffer(60632) := X"00000000";
        ram_buffer(60633) := X"0441FF99";
        ram_buffer(60634) := X"00000000";
        ram_buffer(60635) := X"2402FFFF";
        ram_buffer(60636) := X"AFC20018";
        ram_buffer(60637) := X"1000FF95";
        ram_buffer(60638) := X"00000000";
        ram_buffer(60639) := X"00008021";
        ram_buffer(60640) := X"1000000D";
        ram_buffer(60641) := X"00000000";
        ram_buffer(60642) := X"02001821";
        ram_buffer(60643) := X"00031040";
        ram_buffer(60644) := X"00401821";
        ram_buffer(60645) := X"00031080";
        ram_buffer(60646) := X"00621821";
        ram_buffer(60647) := X"2682FFD0";
        ram_buffer(60648) := X"00628021";
        ram_buffer(60649) := X"02A01021";
        ram_buffer(60650) := X"24550001";
        ram_buffer(60651) := X"80420000";
        ram_buffer(60652) := X"00000000";
        ram_buffer(60653) := X"0040A021";
        ram_buffer(60654) := X"2682FFD0";
        ram_buffer(60655) := X"2C42000A";
        ram_buffer(60656) := X"1440FFF1";
        ram_buffer(60657) := X"00000000";
        ram_buffer(60658) := X"02001021";
        ram_buffer(60659) := X"04410002";
        ram_buffer(60660) := X"00000000";
        ram_buffer(60661) := X"2402FFFF";
        ram_buffer(60662) := X"AFC20018";
        ram_buffer(60663) := X"1000FF80";
        ram_buffer(60664) := X"00000000";
        ram_buffer(60665) := X"36520080";
        ram_buffer(60666) := X"1000FF78";
        ram_buffer(60667) := X"00000000";
        ram_buffer(60668) := X"00008021";
        ram_buffer(60669) := X"02001821";
        ram_buffer(60670) := X"00031040";
        ram_buffer(60671) := X"00401821";
        ram_buffer(60672) := X"00031080";
        ram_buffer(60673) := X"00621821";
        ram_buffer(60674) := X"2682FFD0";
        ram_buffer(60675) := X"00628021";
        ram_buffer(60676) := X"02A01021";
        ram_buffer(60677) := X"24550001";
        ram_buffer(60678) := X"80420000";
        ram_buffer(60679) := X"00000000";
        ram_buffer(60680) := X"0040A021";
        ram_buffer(60681) := X"2682FFD0";
        ram_buffer(60682) := X"2C42000A";
        ram_buffer(60683) := X"1440FFF1";
        ram_buffer(60684) := X"00000000";
        ram_buffer(60685) := X"AFD00014";
        ram_buffer(60686) := X"1000FF69";
        ram_buffer(60687) := X"00000000";
        ram_buffer(60688) := X"82A30000";
        ram_buffer(60689) := X"24020068";
        ram_buffer(60690) := X"14620005";
        ram_buffer(60691) := X"00000000";
        ram_buffer(60692) := X"26B50001";
        ram_buffer(60693) := X"36520200";
        ram_buffer(60694) := X"1000FF5C";
        ram_buffer(60695) := X"00000000";
        ram_buffer(60696) := X"36520040";
        ram_buffer(60697) := X"1000FF59";
        ram_buffer(60698) := X"00000000";
        ram_buffer(60699) := X"82A30000";
        ram_buffer(60700) := X"2402006C";
        ram_buffer(60701) := X"14620005";
        ram_buffer(60702) := X"00000000";
        ram_buffer(60703) := X"26B50001";
        ram_buffer(60704) := X"36520020";
        ram_buffer(60705) := X"1000FF51";
        ram_buffer(60706) := X"00000000";
        ram_buffer(60707) := X"36520010";
        ram_buffer(60708) := X"1000FF4E";
        ram_buffer(60709) := X"00000000";
        ram_buffer(60710) := X"36520020";
        ram_buffer(60711) := X"1000FF4B";
        ram_buffer(60712) := X"00000000";
        ram_buffer(60713) := X"36520020";
        ram_buffer(60714) := X"1000FF48";
        ram_buffer(60715) := X"00000000";
        ram_buffer(60716) := X"27D300AC";
        ram_buffer(60717) := X"8FC3019C";
        ram_buffer(60718) := X"00000000";
        ram_buffer(60719) := X"24620004";
        ram_buffer(60720) := X"AFC2019C";
        ram_buffer(60721) := X"8C620000";
        ram_buffer(60722) := X"00000000";
        ram_buffer(60723) := X"00021600";
        ram_buffer(60724) := X"00021603";
        ram_buffer(60725) := X"A2620000";
        ram_buffer(60726) := X"24020001";
        ram_buffer(60727) := X"AFC20044";
        ram_buffer(60728) := X"A3C0005C";
        ram_buffer(60729) := X"1000030A";
        ram_buffer(60730) := X"00000000";
        ram_buffer(60731) := X"36520010";
        ram_buffer(60732) := X"32420020";
        ram_buffer(60733) := X"1040000E";
        ram_buffer(60734) := X"00000000";
        ram_buffer(60735) := X"8FC2019C";
        ram_buffer(60736) := X"00000000";
        ram_buffer(60737) := X"24430007";
        ram_buffer(60738) := X"2402FFF8";
        ram_buffer(60739) := X"00621024";
        ram_buffer(60740) := X"24430008";
        ram_buffer(60741) := X"AFC3019C";
        ram_buffer(60742) := X"8C430004";
        ram_buffer(60743) := X"8C420000";
        ram_buffer(60744) := X"AFC3011C";
        ram_buffer(60745) := X"AFC20118";
        ram_buffer(60746) := X"10000038";
        ram_buffer(60747) := X"00000000";
        ram_buffer(60748) := X"32420010";
        ram_buffer(60749) := X"1040000C";
        ram_buffer(60750) := X"00000000";
        ram_buffer(60751) := X"8FC2019C";
        ram_buffer(60752) := X"00000000";
        ram_buffer(60753) := X"24430004";
        ram_buffer(60754) := X"AFC3019C";
        ram_buffer(60755) := X"8C420000";
        ram_buffer(60756) := X"00000000";
        ram_buffer(60757) := X"AFC2011C";
        ram_buffer(60758) := X"000217C3";
        ram_buffer(60759) := X"AFC20118";
        ram_buffer(60760) := X"1000002A";
        ram_buffer(60761) := X"00000000";
        ram_buffer(60762) := X"32420040";
        ram_buffer(60763) := X"1040000E";
        ram_buffer(60764) := X"00000000";
        ram_buffer(60765) := X"8FC2019C";
        ram_buffer(60766) := X"00000000";
        ram_buffer(60767) := X"24430004";
        ram_buffer(60768) := X"AFC3019C";
        ram_buffer(60769) := X"8C420000";
        ram_buffer(60770) := X"00000000";
        ram_buffer(60771) := X"00021400";
        ram_buffer(60772) := X"00021403";
        ram_buffer(60773) := X"AFC2011C";
        ram_buffer(60774) := X"000217C3";
        ram_buffer(60775) := X"AFC20118";
        ram_buffer(60776) := X"1000001A";
        ram_buffer(60777) := X"00000000";
        ram_buffer(60778) := X"32420200";
        ram_buffer(60779) := X"1040000E";
        ram_buffer(60780) := X"00000000";
        ram_buffer(60781) := X"8FC2019C";
        ram_buffer(60782) := X"00000000";
        ram_buffer(60783) := X"24430004";
        ram_buffer(60784) := X"AFC3019C";
        ram_buffer(60785) := X"8C420000";
        ram_buffer(60786) := X"00000000";
        ram_buffer(60787) := X"00021600";
        ram_buffer(60788) := X"00021603";
        ram_buffer(60789) := X"AFC2011C";
        ram_buffer(60790) := X"000217C3";
        ram_buffer(60791) := X"AFC20118";
        ram_buffer(60792) := X"1000000A";
        ram_buffer(60793) := X"00000000";
        ram_buffer(60794) := X"8FC2019C";
        ram_buffer(60795) := X"00000000";
        ram_buffer(60796) := X"24430004";
        ram_buffer(60797) := X"AFC3019C";
        ram_buffer(60798) := X"8C420000";
        ram_buffer(60799) := X"00000000";
        ram_buffer(60800) := X"AFC2011C";
        ram_buffer(60801) := X"000217C3";
        ram_buffer(60802) := X"AFC20118";
        ram_buffer(60803) := X"8FC3011C";
        ram_buffer(60804) := X"8FC20118";
        ram_buffer(60805) := X"AFC30034";
        ram_buffer(60806) := X"AFC20030";
        ram_buffer(60807) := X"8FC30034";
        ram_buffer(60808) := X"8FC20030";
        ram_buffer(60809) := X"00000000";
        ram_buffer(60810) := X"0441000E";
        ram_buffer(60811) := X"00000000";
        ram_buffer(60812) := X"00001821";
        ram_buffer(60813) := X"00001021";
        ram_buffer(60814) := X"8FC50034";
        ram_buffer(60815) := X"8FC40030";
        ram_buffer(60816) := X"00653823";
        ram_buffer(60817) := X"0067402B";
        ram_buffer(60818) := X"00443023";
        ram_buffer(60819) := X"00C81023";
        ram_buffer(60820) := X"00403021";
        ram_buffer(60821) := X"AFC70034";
        ram_buffer(60822) := X"AFC60030";
        ram_buffer(60823) := X"2402002D";
        ram_buffer(60824) := X"A3C2005C";
        ram_buffer(60825) := X"24020001";
        ram_buffer(60826) := X"A3C20038";
        ram_buffer(60827) := X"100001AB";
        ram_buffer(60828) := X"00000000";
        ram_buffer(60829) := X"32420020";
        ram_buffer(60830) := X"10400011";
        ram_buffer(60831) := X"00000000";
        ram_buffer(60832) := X"8FC2019C";
        ram_buffer(60833) := X"00000000";
        ram_buffer(60834) := X"24430004";
        ram_buffer(60835) := X"AFC3019C";
        ram_buffer(60836) := X"8C430000";
        ram_buffer(60837) := X"8FC20010";
        ram_buffer(60838) := X"00000000";
        ram_buffer(60839) := X"AFC20134";
        ram_buffer(60840) := X"000217C3";
        ram_buffer(60841) := X"AFC20130";
        ram_buffer(60842) := X"8FC50134";
        ram_buffer(60843) := X"8FC40130";
        ram_buffer(60844) := X"AC650004";
        ram_buffer(60845) := X"AC640000";
        ram_buffer(60846) := X"10000441";
        ram_buffer(60847) := X"00000000";
        ram_buffer(60848) := X"32420010";
        ram_buffer(60849) := X"1040000B";
        ram_buffer(60850) := X"00000000";
        ram_buffer(60851) := X"8FC2019C";
        ram_buffer(60852) := X"00000000";
        ram_buffer(60853) := X"24430004";
        ram_buffer(60854) := X"AFC3019C";
        ram_buffer(60855) := X"8C420000";
        ram_buffer(60856) := X"8FC30010";
        ram_buffer(60857) := X"00000000";
        ram_buffer(60858) := X"AC430000";
        ram_buffer(60859) := X"10000434";
        ram_buffer(60860) := X"00000000";
        ram_buffer(60861) := X"32420040";
        ram_buffer(60862) := X"1040000D";
        ram_buffer(60863) := X"00000000";
        ram_buffer(60864) := X"8FC2019C";
        ram_buffer(60865) := X"00000000";
        ram_buffer(60866) := X"24430004";
        ram_buffer(60867) := X"AFC3019C";
        ram_buffer(60868) := X"8C420000";
        ram_buffer(60869) := X"8FC30010";
        ram_buffer(60870) := X"00000000";
        ram_buffer(60871) := X"00031C00";
        ram_buffer(60872) := X"00031C03";
        ram_buffer(60873) := X"A4430000";
        ram_buffer(60874) := X"10000425";
        ram_buffer(60875) := X"00000000";
        ram_buffer(60876) := X"32420200";
        ram_buffer(60877) := X"1040000D";
        ram_buffer(60878) := X"00000000";
        ram_buffer(60879) := X"8FC2019C";
        ram_buffer(60880) := X"00000000";
        ram_buffer(60881) := X"24430004";
        ram_buffer(60882) := X"AFC3019C";
        ram_buffer(60883) := X"8C420000";
        ram_buffer(60884) := X"8FC30010";
        ram_buffer(60885) := X"00000000";
        ram_buffer(60886) := X"00031E00";
        ram_buffer(60887) := X"00031E03";
        ram_buffer(60888) := X"A0430000";
        ram_buffer(60889) := X"10000416";
        ram_buffer(60890) := X"00000000";
        ram_buffer(60891) := X"8FC2019C";
        ram_buffer(60892) := X"00000000";
        ram_buffer(60893) := X"24430004";
        ram_buffer(60894) := X"AFC3019C";
        ram_buffer(60895) := X"8C420000";
        ram_buffer(60896) := X"8FC30010";
        ram_buffer(60897) := X"00000000";
        ram_buffer(60898) := X"AC430000";
        ram_buffer(60899) := X"1000040C";
        ram_buffer(60900) := X"00000000";
        ram_buffer(60901) := X"36520010";
        ram_buffer(60902) := X"32420020";
        ram_buffer(60903) := X"1040000C";
        ram_buffer(60904) := X"00000000";
        ram_buffer(60905) := X"8FC2019C";
        ram_buffer(60906) := X"00000000";
        ram_buffer(60907) := X"24430007";
        ram_buffer(60908) := X"2402FFF8";
        ram_buffer(60909) := X"00621024";
        ram_buffer(60910) := X"24430008";
        ram_buffer(60911) := X"AFC3019C";
        ram_buffer(60912) := X"8C570004";
        ram_buffer(60913) := X"8C560000";
        ram_buffer(60914) := X"1000003C";
        ram_buffer(60915) := X"00000000";
        ram_buffer(60916) := X"32420010";
        ram_buffer(60917) := X"1040000B";
        ram_buffer(60918) := X"00000000";
        ram_buffer(60919) := X"8FC2019C";
        ram_buffer(60920) := X"00000000";
        ram_buffer(60921) := X"24430004";
        ram_buffer(60922) := X"AFC3019C";
        ram_buffer(60923) := X"8C420000";
        ram_buffer(60924) := X"00000000";
        ram_buffer(60925) := X"0040B821";
        ram_buffer(60926) := X"0000B021";
        ram_buffer(60927) := X"1000002F";
        ram_buffer(60928) := X"00000000";
        ram_buffer(60929) := X"32420040";
        ram_buffer(60930) := X"10400011";
        ram_buffer(60931) := X"00000000";
        ram_buffer(60932) := X"8FC2019C";
        ram_buffer(60933) := X"00000000";
        ram_buffer(60934) := X"24430004";
        ram_buffer(60935) := X"AFC3019C";
        ram_buffer(60936) := X"8C420000";
        ram_buffer(60937) := X"00000000";
        ram_buffer(60938) := X"AFC2013C";
        ram_buffer(60939) := X"AFC00138";
        ram_buffer(60940) := X"8FC3013C";
        ram_buffer(60941) := X"8FC20138";
        ram_buffer(60942) := X"00000000";
        ram_buffer(60943) := X"00402021";
        ram_buffer(60944) := X"30960000";
        ram_buffer(60945) := X"3077FFFF";
        ram_buffer(60946) := X"1000001C";
        ram_buffer(60947) := X"00000000";
        ram_buffer(60948) := X"32420200";
        ram_buffer(60949) := X"10400011";
        ram_buffer(60950) := X"00000000";
        ram_buffer(60951) := X"8FC2019C";
        ram_buffer(60952) := X"00000000";
        ram_buffer(60953) := X"24430004";
        ram_buffer(60954) := X"AFC3019C";
        ram_buffer(60955) := X"8C420000";
        ram_buffer(60956) := X"00000000";
        ram_buffer(60957) := X"AFC20144";
        ram_buffer(60958) := X"AFC00140";
        ram_buffer(60959) := X"8FC30144";
        ram_buffer(60960) := X"8FC20140";
        ram_buffer(60961) := X"00000000";
        ram_buffer(60962) := X"00402021";
        ram_buffer(60963) := X"30960000";
        ram_buffer(60964) := X"307700FF";
        ram_buffer(60965) := X"10000009";
        ram_buffer(60966) := X"00000000";
        ram_buffer(60967) := X"8FC2019C";
        ram_buffer(60968) := X"00000000";
        ram_buffer(60969) := X"24430004";
        ram_buffer(60970) := X"AFC3019C";
        ram_buffer(60971) := X"8C420000";
        ram_buffer(60972) := X"00000000";
        ram_buffer(60973) := X"0040B821";
        ram_buffer(60974) := X"0000B021";
        ram_buffer(60975) := X"AFD70034";
        ram_buffer(60976) := X"AFD60030";
        ram_buffer(60977) := X"A3C00038";
        ram_buffer(60978) := X"2402FBFF";
        ram_buffer(60979) := X"02429024";
        ram_buffer(60980) := X"10000111";
        ram_buffer(60981) := X"00000000";
        ram_buffer(60982) := X"8FC2019C";
        ram_buffer(60983) := X"00000000";
        ram_buffer(60984) := X"24430004";
        ram_buffer(60985) := X"AFC3019C";
        ram_buffer(60986) := X"8C420000";
        ram_buffer(60987) := X"00000000";
        ram_buffer(60988) := X"AFC20034";
        ram_buffer(60989) := X"AFC00030";
        ram_buffer(60990) := X"24020002";
        ram_buffer(60991) := X"A3C20038";
        ram_buffer(60992) := X"3C02100D";
        ram_buffer(60993) := X"2442B0B8";
        ram_buffer(60994) := X"AFC20048";
        ram_buffer(60995) := X"36520002";
        ram_buffer(60996) := X"24020030";
        ram_buffer(60997) := X"A3C20110";
        ram_buffer(60998) := X"24140078";
        ram_buffer(60999) := X"24020078";
        ram_buffer(61000) := X"A3C20111";
        ram_buffer(61001) := X"100000FC";
        ram_buffer(61002) := X"00000000";
        ram_buffer(61003) := X"8FC2019C";
        ram_buffer(61004) := X"00000000";
        ram_buffer(61005) := X"24430004";
        ram_buffer(61006) := X"AFC3019C";
        ram_buffer(61007) := X"8C530000";
        ram_buffer(61008) := X"A3C0005C";
        ram_buffer(61009) := X"1660000D";
        ram_buffer(61010) := X"00000000";
        ram_buffer(61011) := X"3C02100D";
        ram_buffer(61012) := X"2453B0CC";
        ram_buffer(61013) := X"8FC20018";
        ram_buffer(61014) := X"00000000";
        ram_buffer(61015) := X"00401821";
        ram_buffer(61016) := X"2C620007";
        ram_buffer(61017) := X"14400002";
        ram_buffer(61018) := X"00000000";
        ram_buffer(61019) := X"24030006";
        ram_buffer(61020) := X"AFC30044";
        ram_buffer(61021) := X"100001E6";
        ram_buffer(61022) := X"00000000";
        ram_buffer(61023) := X"8FC20018";
        ram_buffer(61024) := X"00000000";
        ram_buffer(61025) := X"04400018";
        ram_buffer(61026) := X"00000000";
        ram_buffer(61027) := X"8FC20018";
        ram_buffer(61028) := X"00000000";
        ram_buffer(61029) := X"00403021";
        ram_buffer(61030) := X"00002821";
        ram_buffer(61031) := X"02602021";
        ram_buffer(61032) := X"0C02BC51";
        ram_buffer(61033) := X"00000000";
        ram_buffer(61034) := X"AFC20058";
        ram_buffer(61035) := X"8FC20058";
        ram_buffer(61036) := X"00000000";
        ram_buffer(61037) := X"10400007";
        ram_buffer(61038) := X"00000000";
        ram_buffer(61039) := X"8FC30058";
        ram_buffer(61040) := X"02601021";
        ram_buffer(61041) := X"00621023";
        ram_buffer(61042) := X"AFC20044";
        ram_buffer(61043) := X"100001D0";
        ram_buffer(61044) := X"00000000";
        ram_buffer(61045) := X"8FC20018";
        ram_buffer(61046) := X"00000000";
        ram_buffer(61047) := X"AFC20044";
        ram_buffer(61048) := X"100001CB";
        ram_buffer(61049) := X"00000000";
        ram_buffer(61050) := X"02602021";
        ram_buffer(61051) := X"0C02851E";
        ram_buffer(61052) := X"00000000";
        ram_buffer(61053) := X"AFC20044";
        ram_buffer(61054) := X"100001C5";
        ram_buffer(61055) := X"00000000";
        ram_buffer(61056) := X"36520010";
        ram_buffer(61057) := X"32420020";
        ram_buffer(61058) := X"1040000E";
        ram_buffer(61059) := X"00000000";
        ram_buffer(61060) := X"8FC2019C";
        ram_buffer(61061) := X"00000000";
        ram_buffer(61062) := X"24430007";
        ram_buffer(61063) := X"2402FFF8";
        ram_buffer(61064) := X"00621024";
        ram_buffer(61065) := X"24430008";
        ram_buffer(61066) := X"AFC3019C";
        ram_buffer(61067) := X"8C430004";
        ram_buffer(61068) := X"8C420000";
        ram_buffer(61069) := X"AFC30124";
        ram_buffer(61070) := X"AFC20120";
        ram_buffer(61071) := X"10000040";
        ram_buffer(61072) := X"00000000";
        ram_buffer(61073) := X"32420010";
        ram_buffer(61074) := X"1040000B";
        ram_buffer(61075) := X"00000000";
        ram_buffer(61076) := X"8FC2019C";
        ram_buffer(61077) := X"00000000";
        ram_buffer(61078) := X"24430004";
        ram_buffer(61079) := X"AFC3019C";
        ram_buffer(61080) := X"8C420000";
        ram_buffer(61081) := X"00000000";
        ram_buffer(61082) := X"AFC20124";
        ram_buffer(61083) := X"AFC00120";
        ram_buffer(61084) := X"10000033";
        ram_buffer(61085) := X"00000000";
        ram_buffer(61086) := X"32420040";
        ram_buffer(61087) := X"10400013";
        ram_buffer(61088) := X"00000000";
        ram_buffer(61089) := X"8FC2019C";
        ram_buffer(61090) := X"00000000";
        ram_buffer(61091) := X"24430004";
        ram_buffer(61092) := X"AFC3019C";
        ram_buffer(61093) := X"8C420000";
        ram_buffer(61094) := X"00000000";
        ram_buffer(61095) := X"AFC2014C";
        ram_buffer(61096) := X"AFC00148";
        ram_buffer(61097) := X"8FC3014C";
        ram_buffer(61098) := X"8FC20148";
        ram_buffer(61099) := X"00000000";
        ram_buffer(61100) := X"00402021";
        ram_buffer(61101) := X"30840000";
        ram_buffer(61102) := X"AFC40120";
        ram_buffer(61103) := X"3062FFFF";
        ram_buffer(61104) := X"AFC20124";
        ram_buffer(61105) := X"1000001E";
        ram_buffer(61106) := X"00000000";
        ram_buffer(61107) := X"32420200";
        ram_buffer(61108) := X"10400013";
        ram_buffer(61109) := X"00000000";
        ram_buffer(61110) := X"8FC2019C";
        ram_buffer(61111) := X"00000000";
        ram_buffer(61112) := X"24430004";
        ram_buffer(61113) := X"AFC3019C";
        ram_buffer(61114) := X"8C420000";
        ram_buffer(61115) := X"00000000";
        ram_buffer(61116) := X"AFC20154";
        ram_buffer(61117) := X"AFC00150";
        ram_buffer(61118) := X"8FC30154";
        ram_buffer(61119) := X"8FC20150";
        ram_buffer(61120) := X"00000000";
        ram_buffer(61121) := X"00402021";
        ram_buffer(61122) := X"30840000";
        ram_buffer(61123) := X"AFC40120";
        ram_buffer(61124) := X"306200FF";
        ram_buffer(61125) := X"AFC20124";
        ram_buffer(61126) := X"10000009";
        ram_buffer(61127) := X"00000000";
        ram_buffer(61128) := X"8FC2019C";
        ram_buffer(61129) := X"00000000";
        ram_buffer(61130) := X"24430004";
        ram_buffer(61131) := X"AFC3019C";
        ram_buffer(61132) := X"8C420000";
        ram_buffer(61133) := X"00000000";
        ram_buffer(61134) := X"AFC20124";
        ram_buffer(61135) := X"AFC00120";
        ram_buffer(61136) := X"8FC30124";
        ram_buffer(61137) := X"8FC20120";
        ram_buffer(61138) := X"AFC30034";
        ram_buffer(61139) := X"AFC20030";
        ram_buffer(61140) := X"24020001";
        ram_buffer(61141) := X"A3C20038";
        ram_buffer(61142) := X"1000006F";
        ram_buffer(61143) := X"00000000";
        ram_buffer(61144) := X"3C02100D";
        ram_buffer(61145) := X"2442B0D4";
        ram_buffer(61146) := X"AFC20048";
        ram_buffer(61147) := X"10000004";
        ram_buffer(61148) := X"00000000";
        ram_buffer(61149) := X"3C02100D";
        ram_buffer(61150) := X"2442B0B8";
        ram_buffer(61151) := X"AFC20048";
        ram_buffer(61152) := X"32420020";
        ram_buffer(61153) := X"1040000E";
        ram_buffer(61154) := X"00000000";
        ram_buffer(61155) := X"8FC2019C";
        ram_buffer(61156) := X"00000000";
        ram_buffer(61157) := X"24430007";
        ram_buffer(61158) := X"2402FFF8";
        ram_buffer(61159) := X"00621024";
        ram_buffer(61160) := X"24430008";
        ram_buffer(61161) := X"AFC3019C";
        ram_buffer(61162) := X"8C430004";
        ram_buffer(61163) := X"8C420000";
        ram_buffer(61164) := X"AFC3012C";
        ram_buffer(61165) := X"AFC20128";
        ram_buffer(61166) := X"10000040";
        ram_buffer(61167) := X"00000000";
        ram_buffer(61168) := X"32420010";
        ram_buffer(61169) := X"1040000B";
        ram_buffer(61170) := X"00000000";
        ram_buffer(61171) := X"8FC3019C";
        ram_buffer(61172) := X"00000000";
        ram_buffer(61173) := X"24620004";
        ram_buffer(61174) := X"AFC2019C";
        ram_buffer(61175) := X"8C620000";
        ram_buffer(61176) := X"00000000";
        ram_buffer(61177) := X"AFC2012C";
        ram_buffer(61178) := X"AFC00128";
        ram_buffer(61179) := X"10000033";
        ram_buffer(61180) := X"00000000";
        ram_buffer(61181) := X"32420040";
        ram_buffer(61182) := X"10400013";
        ram_buffer(61183) := X"00000000";
        ram_buffer(61184) := X"8FC3019C";
        ram_buffer(61185) := X"00000000";
        ram_buffer(61186) := X"24620004";
        ram_buffer(61187) := X"AFC2019C";
        ram_buffer(61188) := X"8C620000";
        ram_buffer(61189) := X"00000000";
        ram_buffer(61190) := X"AFC2015C";
        ram_buffer(61191) := X"AFC00158";
        ram_buffer(61192) := X"8FC3015C";
        ram_buffer(61193) := X"8FC20158";
        ram_buffer(61194) := X"00000000";
        ram_buffer(61195) := X"00402021";
        ram_buffer(61196) := X"30840000";
        ram_buffer(61197) := X"AFC40128";
        ram_buffer(61198) := X"3062FFFF";
        ram_buffer(61199) := X"AFC2012C";
        ram_buffer(61200) := X"1000001E";
        ram_buffer(61201) := X"00000000";
        ram_buffer(61202) := X"32420200";
        ram_buffer(61203) := X"10400013";
        ram_buffer(61204) := X"00000000";
        ram_buffer(61205) := X"8FC3019C";
        ram_buffer(61206) := X"00000000";
        ram_buffer(61207) := X"24620004";
        ram_buffer(61208) := X"AFC2019C";
        ram_buffer(61209) := X"8C620000";
        ram_buffer(61210) := X"00000000";
        ram_buffer(61211) := X"AFC20164";
        ram_buffer(61212) := X"AFC00160";
        ram_buffer(61213) := X"8FC30164";
        ram_buffer(61214) := X"8FC20160";
        ram_buffer(61215) := X"00000000";
        ram_buffer(61216) := X"00402021";
        ram_buffer(61217) := X"30840000";
        ram_buffer(61218) := X"AFC40128";
        ram_buffer(61219) := X"306200FF";
        ram_buffer(61220) := X"AFC2012C";
        ram_buffer(61221) := X"10000009";
        ram_buffer(61222) := X"00000000";
        ram_buffer(61223) := X"8FC3019C";
        ram_buffer(61224) := X"00000000";
        ram_buffer(61225) := X"24620004";
        ram_buffer(61226) := X"AFC2019C";
        ram_buffer(61227) := X"8C620000";
        ram_buffer(61228) := X"00000000";
        ram_buffer(61229) := X"AFC2012C";
        ram_buffer(61230) := X"AFC00128";
        ram_buffer(61231) := X"8FC3012C";
        ram_buffer(61232) := X"8FC20128";
        ram_buffer(61233) := X"AFC30034";
        ram_buffer(61234) := X"AFC20030";
        ram_buffer(61235) := X"24020002";
        ram_buffer(61236) := X"A3C20038";
        ram_buffer(61237) := X"32420001";
        ram_buffer(61238) := X"1040000D";
        ram_buffer(61239) := X"00000000";
        ram_buffer(61240) := X"8FC20030";
        ram_buffer(61241) := X"8FC30034";
        ram_buffer(61242) := X"00000000";
        ram_buffer(61243) := X"00431025";
        ram_buffer(61244) := X"10400007";
        ram_buffer(61245) := X"00000000";
        ram_buffer(61246) := X"24020030";
        ram_buffer(61247) := X"A3C20110";
        ram_buffer(61248) := X"00141600";
        ram_buffer(61249) := X"00021603";
        ram_buffer(61250) := X"A3C20111";
        ram_buffer(61251) := X"36520002";
        ram_buffer(61252) := X"2402FBFF";
        ram_buffer(61253) := X"02429024";
        ram_buffer(61254) := X"A3C0005C";
        ram_buffer(61255) := X"8FC20018";
        ram_buffer(61256) := X"00000000";
        ram_buffer(61257) := X"AFC2003C";
        ram_buffer(61258) := X"8FC2003C";
        ram_buffer(61259) := X"00000000";
        ram_buffer(61260) := X"04400003";
        ram_buffer(61261) := X"00000000";
        ram_buffer(61262) := X"2402FF7F";
        ram_buffer(61263) := X"02429024";
        ram_buffer(61264) := X"27D300AC";
        ram_buffer(61265) := X"26730064";
        ram_buffer(61266) := X"8FC20030";
        ram_buffer(61267) := X"8FC30034";
        ram_buffer(61268) := X"00000000";
        ram_buffer(61269) := X"00431025";
        ram_buffer(61270) := X"14400005";
        ram_buffer(61271) := X"00000000";
        ram_buffer(61272) := X"8FC20018";
        ram_buffer(61273) := X"00000000";
        ram_buffer(61274) := X"104000CD";
        ram_buffer(61275) := X"00000000";
        ram_buffer(61276) := X"93C30038";
        ram_buffer(61277) := X"24020001";
        ram_buffer(61278) := X"1062002E";
        ram_buffer(61279) := X"00000000";
        ram_buffer(61280) := X"24020002";
        ram_buffer(61281) := X"1062009C";
        ram_buffer(61282) := X"00000000";
        ram_buffer(61283) := X"146000B8";
        ram_buffer(61284) := X"00000000";
        ram_buffer(61285) := X"2673FFFF";
        ram_buffer(61286) := X"93C20037";
        ram_buffer(61287) := X"00000000";
        ram_buffer(61288) := X"30420007";
        ram_buffer(61289) := X"304200FF";
        ram_buffer(61290) := X"24420030";
        ram_buffer(61291) := X"304200FF";
        ram_buffer(61292) := X"00021600";
        ram_buffer(61293) := X"00021603";
        ram_buffer(61294) := X"A2620000";
        ram_buffer(61295) := X"8FC20030";
        ram_buffer(61296) := X"00000000";
        ram_buffer(61297) := X"00021F40";
        ram_buffer(61298) := X"8FC20034";
        ram_buffer(61299) := X"00000000";
        ram_buffer(61300) := X"000210C2";
        ram_buffer(61301) := X"00431025";
        ram_buffer(61302) := X"AFC20034";
        ram_buffer(61303) := X"8FC20030";
        ram_buffer(61304) := X"00000000";
        ram_buffer(61305) := X"000210C2";
        ram_buffer(61306) := X"AFC20030";
        ram_buffer(61307) := X"8FC20030";
        ram_buffer(61308) := X"8FC30034";
        ram_buffer(61309) := X"00000000";
        ram_buffer(61310) := X"00431025";
        ram_buffer(61311) := X"1440FFE5";
        ram_buffer(61312) := X"00000000";
        ram_buffer(61313) := X"32420001";
        ram_buffer(61314) := X"104000A2";
        ram_buffer(61315) := X"00000000";
        ram_buffer(61316) := X"82630000";
        ram_buffer(61317) := X"24020030";
        ram_buffer(61318) := X"1062009E";
        ram_buffer(61319) := X"00000000";
        ram_buffer(61320) := X"2673FFFF";
        ram_buffer(61321) := X"24020030";
        ram_buffer(61322) := X"A2620000";
        ram_buffer(61323) := X"10000099";
        ram_buffer(61324) := X"00000000";
        ram_buffer(61325) := X"8FC20030";
        ram_buffer(61326) := X"00000000";
        ram_buffer(61327) := X"14400014";
        ram_buffer(61328) := X"00000000";
        ram_buffer(61329) := X"8FC20030";
        ram_buffer(61330) := X"00000000";
        ram_buffer(61331) := X"14400006";
        ram_buffer(61332) := X"00000000";
        ram_buffer(61333) := X"8FC20034";
        ram_buffer(61334) := X"00000000";
        ram_buffer(61335) := X"2C42000A";
        ram_buffer(61336) := X"1040000B";
        ram_buffer(61337) := X"00000000";
        ram_buffer(61338) := X"2673FFFF";
        ram_buffer(61339) := X"93C20037";
        ram_buffer(61340) := X"00000000";
        ram_buffer(61341) := X"24420030";
        ram_buffer(61342) := X"304200FF";
        ram_buffer(61343) := X"00021600";
        ram_buffer(61344) := X"00021603";
        ram_buffer(61345) := X"A2620000";
        ram_buffer(61346) := X"10000083";
        ram_buffer(61347) := X"00000000";
        ram_buffer(61348) := X"AFC00028";
        ram_buffer(61349) := X"2673FFFF";
        ram_buffer(61350) := X"8FC30034";
        ram_buffer(61351) := X"8FC20030";
        ram_buffer(61352) := X"2407000A";
        ram_buffer(61353) := X"00003021";
        ram_buffer(61354) := X"00602821";
        ram_buffer(61355) := X"00402021";
        ram_buffer(61356) := X"0C030BFE";
        ram_buffer(61357) := X"00000000";
        ram_buffer(61358) := X"306200FF";
        ram_buffer(61359) := X"24420030";
        ram_buffer(61360) := X"304200FF";
        ram_buffer(61361) := X"00021600";
        ram_buffer(61362) := X"00021603";
        ram_buffer(61363) := X"A2620000";
        ram_buffer(61364) := X"8FC20028";
        ram_buffer(61365) := X"00000000";
        ram_buffer(61366) := X"24420001";
        ram_buffer(61367) := X"AFC20028";
        ram_buffer(61368) := X"32420400";
        ram_buffer(61369) := X"10400032";
        ram_buffer(61370) := X"00000000";
        ram_buffer(61371) := X"8FC20024";
        ram_buffer(61372) := X"00000000";
        ram_buffer(61373) := X"80420000";
        ram_buffer(61374) := X"00000000";
        ram_buffer(61375) := X"00401821";
        ram_buffer(61376) := X"8FC20028";
        ram_buffer(61377) := X"00000000";
        ram_buffer(61378) := X"14620029";
        ram_buffer(61379) := X"00000000";
        ram_buffer(61380) := X"8FC20024";
        ram_buffer(61381) := X"00000000";
        ram_buffer(61382) := X"80430000";
        ram_buffer(61383) := X"2402007F";
        ram_buffer(61384) := X"10620023";
        ram_buffer(61385) := X"00000000";
        ram_buffer(61386) := X"8FC20030";
        ram_buffer(61387) := X"00000000";
        ram_buffer(61388) := X"1440000A";
        ram_buffer(61389) := X"00000000";
        ram_buffer(61390) := X"8FC20030";
        ram_buffer(61391) := X"00000000";
        ram_buffer(61392) := X"1440001B";
        ram_buffer(61393) := X"00000000";
        ram_buffer(61394) := X"8FC20034";
        ram_buffer(61395) := X"00000000";
        ram_buffer(61396) := X"2C42000A";
        ram_buffer(61397) := X"14400016";
        ram_buffer(61398) := X"00000000";
        ram_buffer(61399) := X"8FC20020";
        ram_buffer(61400) := X"00000000";
        ram_buffer(61401) := X"00021023";
        ram_buffer(61402) := X"02629821";
        ram_buffer(61403) := X"8FC60020";
        ram_buffer(61404) := X"8FC5001C";
        ram_buffer(61405) := X"02602021";
        ram_buffer(61406) := X"0C02CCBF";
        ram_buffer(61407) := X"00000000";
        ram_buffer(61408) := X"AFC00028";
        ram_buffer(61409) := X"8FC20024";
        ram_buffer(61410) := X"00000000";
        ram_buffer(61411) := X"24420001";
        ram_buffer(61412) := X"80420000";
        ram_buffer(61413) := X"00000000";
        ram_buffer(61414) := X"10400005";
        ram_buffer(61415) := X"00000000";
        ram_buffer(61416) := X"8FC20024";
        ram_buffer(61417) := X"00000000";
        ram_buffer(61418) := X"24420001";
        ram_buffer(61419) := X"AFC20024";
        ram_buffer(61420) := X"8FC30034";
        ram_buffer(61421) := X"8FC20030";
        ram_buffer(61422) := X"2407000A";
        ram_buffer(61423) := X"00003021";
        ram_buffer(61424) := X"00602821";
        ram_buffer(61425) := X"00402021";
        ram_buffer(61426) := X"0C030A67";
        ram_buffer(61427) := X"00000000";
        ram_buffer(61428) := X"AFC30034";
        ram_buffer(61429) := X"AFC20030";
        ram_buffer(61430) := X"8FC20030";
        ram_buffer(61431) := X"8FC30034";
        ram_buffer(61432) := X"00000000";
        ram_buffer(61433) := X"00431025";
        ram_buffer(61434) := X"1440FFAA";
        ram_buffer(61435) := X"00000000";
        ram_buffer(61436) := X"10000029";
        ram_buffer(61437) := X"00000000";
        ram_buffer(61438) := X"2673FFFF";
        ram_buffer(61439) := X"8FC20034";
        ram_buffer(61440) := X"00000000";
        ram_buffer(61441) := X"3043000F";
        ram_buffer(61442) := X"8FC20048";
        ram_buffer(61443) := X"00000000";
        ram_buffer(61444) := X"00431021";
        ram_buffer(61445) := X"80420000";
        ram_buffer(61446) := X"00000000";
        ram_buffer(61447) := X"A2620000";
        ram_buffer(61448) := X"8FC20030";
        ram_buffer(61449) := X"00000000";
        ram_buffer(61450) := X"00021F00";
        ram_buffer(61451) := X"8FC20034";
        ram_buffer(61452) := X"00000000";
        ram_buffer(61453) := X"00021102";
        ram_buffer(61454) := X"00431025";
        ram_buffer(61455) := X"AFC20034";
        ram_buffer(61456) := X"8FC20030";
        ram_buffer(61457) := X"00000000";
        ram_buffer(61458) := X"00021102";
        ram_buffer(61459) := X"AFC20030";
        ram_buffer(61460) := X"8FC20030";
        ram_buffer(61461) := X"8FC30034";
        ram_buffer(61462) := X"00000000";
        ram_buffer(61463) := X"00431025";
        ram_buffer(61464) := X"1440FFE5";
        ram_buffer(61465) := X"00000000";
        ram_buffer(61466) := X"1000000B";
        ram_buffer(61467) := X"00000000";
        ram_buffer(61468) := X"3C02100D";
        ram_buffer(61469) := X"2453B0E8";
        ram_buffer(61470) := X"02602021";
        ram_buffer(61471) := X"0C02851E";
        ram_buffer(61472) := X"00000000";
        ram_buffer(61473) := X"AFC20044";
        ram_buffer(61474) := X"00000000";
        ram_buffer(61475) := X"10000020";
        ram_buffer(61476) := X"00000000";
        ram_buffer(61477) := X"00000000";
        ram_buffer(61478) := X"1000000B";
        ram_buffer(61479) := X"00000000";
        ram_buffer(61480) := X"93C20038";
        ram_buffer(61481) := X"00000000";
        ram_buffer(61482) := X"14400007";
        ram_buffer(61483) := X"00000000";
        ram_buffer(61484) := X"32420001";
        ram_buffer(61485) := X"10400004";
        ram_buffer(61486) := X"00000000";
        ram_buffer(61487) := X"2673FFFF";
        ram_buffer(61488) := X"24020030";
        ram_buffer(61489) := X"A2620000";
        ram_buffer(61490) := X"27C200AC";
        ram_buffer(61491) := X"24420064";
        ram_buffer(61492) := X"00401821";
        ram_buffer(61493) := X"02601021";
        ram_buffer(61494) := X"00621023";
        ram_buffer(61495) := X"AFC20044";
        ram_buffer(61496) := X"1000000B";
        ram_buffer(61497) := X"00000000";
        ram_buffer(61498) := X"128001BA";
        ram_buffer(61499) := X"00000000";
        ram_buffer(61500) := X"27D300AC";
        ram_buffer(61501) := X"00141600";
        ram_buffer(61502) := X"00021603";
        ram_buffer(61503) := X"A2620000";
        ram_buffer(61504) := X"24020001";
        ram_buffer(61505) := X"AFC20044";
        ram_buffer(61506) := X"A3C0005C";
        ram_buffer(61507) := X"00000000";
        ram_buffer(61508) := X"8FC4003C";
        ram_buffer(61509) := X"8FC30044";
        ram_buffer(61510) := X"00000000";
        ram_buffer(61511) := X"0064102A";
        ram_buffer(61512) := X"10400002";
        ram_buffer(61513) := X"00000000";
        ram_buffer(61514) := X"00801821";
        ram_buffer(61515) := X"AFC30040";
        ram_buffer(61516) := X"83C2005C";
        ram_buffer(61517) := X"00000000";
        ram_buffer(61518) := X"10400005";
        ram_buffer(61519) := X"00000000";
        ram_buffer(61520) := X"8FC20040";
        ram_buffer(61521) := X"00000000";
        ram_buffer(61522) := X"24420001";
        ram_buffer(61523) := X"AFC20040";
        ram_buffer(61524) := X"32420002";
        ram_buffer(61525) := X"10400005";
        ram_buffer(61526) := X"00000000";
        ram_buffer(61527) := X"8FC20040";
        ram_buffer(61528) := X"00000000";
        ram_buffer(61529) := X"24420002";
        ram_buffer(61530) := X"AFC20040";
        ram_buffer(61531) := X"32420084";
        ram_buffer(61532) := X"14400045";
        ram_buffer(61533) := X"00000000";
        ram_buffer(61534) := X"8FC30014";
        ram_buffer(61535) := X"8FC20040";
        ram_buffer(61536) := X"00000000";
        ram_buffer(61537) := X"00628023";
        ram_buffer(61538) := X"1A00003F";
        ram_buffer(61539) := X"00000000";
        ram_buffer(61540) := X"1000001E";
        ram_buffer(61541) := X"00000000";
        ram_buffer(61542) := X"3C02100D";
        ram_buffer(61543) := X"2442B270";
        ram_buffer(61544) := X"AE220000";
        ram_buffer(61545) := X"24020010";
        ram_buffer(61546) := X"AE220004";
        ram_buffer(61547) := X"8FC20068";
        ram_buffer(61548) := X"00000000";
        ram_buffer(61549) := X"24420010";
        ram_buffer(61550) := X"AFC20068";
        ram_buffer(61551) := X"26310008";
        ram_buffer(61552) := X"8FC20064";
        ram_buffer(61553) := X"00000000";
        ram_buffer(61554) := X"24420001";
        ram_buffer(61555) := X"AFC20064";
        ram_buffer(61556) := X"8FC20064";
        ram_buffer(61557) := X"00000000";
        ram_buffer(61558) := X"28420008";
        ram_buffer(61559) := X"1440000A";
        ram_buffer(61560) := X"00000000";
        ram_buffer(61561) := X"27C20060";
        ram_buffer(61562) := X"00403021";
        ram_buffer(61563) := X"8FC50194";
        ram_buffer(61564) := X"8FC40190";
        ram_buffer(61565) := X"0C02EAF5";
        ram_buffer(61566) := X"00000000";
        ram_buffer(61567) := X"14400189";
        ram_buffer(61568) := X"00000000";
        ram_buffer(61569) := X"27D1006C";
        ram_buffer(61570) := X"2610FFF0";
        ram_buffer(61571) := X"2A020011";
        ram_buffer(61572) := X"1040FFE1";
        ram_buffer(61573) := X"00000000";
        ram_buffer(61574) := X"3C02100D";
        ram_buffer(61575) := X"2442B270";
        ram_buffer(61576) := X"AE220000";
        ram_buffer(61577) := X"02001021";
        ram_buffer(61578) := X"AE220004";
        ram_buffer(61579) := X"8FC30068";
        ram_buffer(61580) := X"02001021";
        ram_buffer(61581) := X"00621021";
        ram_buffer(61582) := X"AFC20068";
        ram_buffer(61583) := X"26310008";
        ram_buffer(61584) := X"8FC20064";
        ram_buffer(61585) := X"00000000";
        ram_buffer(61586) := X"24420001";
        ram_buffer(61587) := X"AFC20064";
        ram_buffer(61588) := X"8FC20064";
        ram_buffer(61589) := X"00000000";
        ram_buffer(61590) := X"28420008";
        ram_buffer(61591) := X"1440000A";
        ram_buffer(61592) := X"00000000";
        ram_buffer(61593) := X"27C20060";
        ram_buffer(61594) := X"00403021";
        ram_buffer(61595) := X"8FC50194";
        ram_buffer(61596) := X"8FC40190";
        ram_buffer(61597) := X"0C02EAF5";
        ram_buffer(61598) := X"00000000";
        ram_buffer(61599) := X"1440016C";
        ram_buffer(61600) := X"00000000";
        ram_buffer(61601) := X"27D1006C";
        ram_buffer(61602) := X"83C2005C";
        ram_buffer(61603) := X"00000000";
        ram_buffer(61604) := X"1040001C";
        ram_buffer(61605) := X"00000000";
        ram_buffer(61606) := X"27C2005C";
        ram_buffer(61607) := X"AE220000";
        ram_buffer(61608) := X"24020001";
        ram_buffer(61609) := X"AE220004";
        ram_buffer(61610) := X"8FC20068";
        ram_buffer(61611) := X"00000000";
        ram_buffer(61612) := X"24420001";
        ram_buffer(61613) := X"AFC20068";
        ram_buffer(61614) := X"26310008";
        ram_buffer(61615) := X"8FC20064";
        ram_buffer(61616) := X"00000000";
        ram_buffer(61617) := X"24420001";
        ram_buffer(61618) := X"AFC20064";
        ram_buffer(61619) := X"8FC20064";
        ram_buffer(61620) := X"00000000";
        ram_buffer(61621) := X"28420008";
        ram_buffer(61622) := X"1440000A";
        ram_buffer(61623) := X"00000000";
        ram_buffer(61624) := X"27C20060";
        ram_buffer(61625) := X"00403021";
        ram_buffer(61626) := X"8FC50194";
        ram_buffer(61627) := X"8FC40190";
        ram_buffer(61628) := X"0C02EAF5";
        ram_buffer(61629) := X"00000000";
        ram_buffer(61630) := X"14400150";
        ram_buffer(61631) := X"00000000";
        ram_buffer(61632) := X"27D1006C";
        ram_buffer(61633) := X"32420002";
        ram_buffer(61634) := X"1040001C";
        ram_buffer(61635) := X"00000000";
        ram_buffer(61636) := X"27C20110";
        ram_buffer(61637) := X"AE220000";
        ram_buffer(61638) := X"24020002";
        ram_buffer(61639) := X"AE220004";
        ram_buffer(61640) := X"8FC20068";
        ram_buffer(61641) := X"00000000";
        ram_buffer(61642) := X"24420002";
        ram_buffer(61643) := X"AFC20068";
        ram_buffer(61644) := X"26310008";
        ram_buffer(61645) := X"8FC20064";
        ram_buffer(61646) := X"00000000";
        ram_buffer(61647) := X"24420001";
        ram_buffer(61648) := X"AFC20064";
        ram_buffer(61649) := X"8FC20064";
        ram_buffer(61650) := X"00000000";
        ram_buffer(61651) := X"28420008";
        ram_buffer(61652) := X"1440000A";
        ram_buffer(61653) := X"00000000";
        ram_buffer(61654) := X"27C20060";
        ram_buffer(61655) := X"00403021";
        ram_buffer(61656) := X"8FC50194";
        ram_buffer(61657) := X"8FC40190";
        ram_buffer(61658) := X"0C02EAF5";
        ram_buffer(61659) := X"00000000";
        ram_buffer(61660) := X"14400135";
        ram_buffer(61661) := X"00000000";
        ram_buffer(61662) := X"27D1006C";
        ram_buffer(61663) := X"32430084";
        ram_buffer(61664) := X"24020080";
        ram_buffer(61665) := X"14620045";
        ram_buffer(61666) := X"00000000";
        ram_buffer(61667) := X"8FC30014";
        ram_buffer(61668) := X"8FC20040";
        ram_buffer(61669) := X"00000000";
        ram_buffer(61670) := X"00628023";
        ram_buffer(61671) := X"1A00003F";
        ram_buffer(61672) := X"00000000";
        ram_buffer(61673) := X"1000001E";
        ram_buffer(61674) := X"00000000";
        ram_buffer(61675) := X"3C02100D";
        ram_buffer(61676) := X"2442B280";
        ram_buffer(61677) := X"AE220000";
        ram_buffer(61678) := X"24020010";
        ram_buffer(61679) := X"AE220004";
        ram_buffer(61680) := X"8FC20068";
        ram_buffer(61681) := X"00000000";
        ram_buffer(61682) := X"24420010";
        ram_buffer(61683) := X"AFC20068";
        ram_buffer(61684) := X"26310008";
        ram_buffer(61685) := X"8FC20064";
        ram_buffer(61686) := X"00000000";
        ram_buffer(61687) := X"24420001";
        ram_buffer(61688) := X"AFC20064";
        ram_buffer(61689) := X"8FC20064";
        ram_buffer(61690) := X"00000000";
        ram_buffer(61691) := X"28420008";
        ram_buffer(61692) := X"1440000A";
        ram_buffer(61693) := X"00000000";
        ram_buffer(61694) := X"27C20060";
        ram_buffer(61695) := X"00403021";
        ram_buffer(61696) := X"8FC50194";
        ram_buffer(61697) := X"8FC40190";
        ram_buffer(61698) := X"0C02EAF5";
        ram_buffer(61699) := X"00000000";
        ram_buffer(61700) := X"14400110";
        ram_buffer(61701) := X"00000000";
        ram_buffer(61702) := X"27D1006C";
        ram_buffer(61703) := X"2610FFF0";
        ram_buffer(61704) := X"2A020011";
        ram_buffer(61705) := X"1040FFE1";
        ram_buffer(61706) := X"00000000";
        ram_buffer(61707) := X"3C02100D";
        ram_buffer(61708) := X"2442B280";
        ram_buffer(61709) := X"AE220000";
        ram_buffer(61710) := X"02001021";
        ram_buffer(61711) := X"AE220004";
        ram_buffer(61712) := X"8FC30068";
        ram_buffer(61713) := X"02001021";
        ram_buffer(61714) := X"00621021";
        ram_buffer(61715) := X"AFC20068";
        ram_buffer(61716) := X"26310008";
        ram_buffer(61717) := X"8FC20064";
        ram_buffer(61718) := X"00000000";
        ram_buffer(61719) := X"24420001";
        ram_buffer(61720) := X"AFC20064";
        ram_buffer(61721) := X"8FC20064";
        ram_buffer(61722) := X"00000000";
        ram_buffer(61723) := X"28420008";
        ram_buffer(61724) := X"1440000A";
        ram_buffer(61725) := X"00000000";
        ram_buffer(61726) := X"27C20060";
        ram_buffer(61727) := X"00403021";
        ram_buffer(61728) := X"8FC50194";
        ram_buffer(61729) := X"8FC40190";
        ram_buffer(61730) := X"0C02EAF5";
        ram_buffer(61731) := X"00000000";
        ram_buffer(61732) := X"144000F3";
        ram_buffer(61733) := X"00000000";
        ram_buffer(61734) := X"27D1006C";
        ram_buffer(61735) := X"8FC3003C";
        ram_buffer(61736) := X"8FC20044";
        ram_buffer(61737) := X"00000000";
        ram_buffer(61738) := X"00628023";
        ram_buffer(61739) := X"1A00003F";
        ram_buffer(61740) := X"00000000";
        ram_buffer(61741) := X"1000001E";
        ram_buffer(61742) := X"00000000";
        ram_buffer(61743) := X"3C02100D";
        ram_buffer(61744) := X"2442B280";
        ram_buffer(61745) := X"AE220000";
        ram_buffer(61746) := X"24020010";
        ram_buffer(61747) := X"AE220004";
        ram_buffer(61748) := X"8FC20068";
        ram_buffer(61749) := X"00000000";
        ram_buffer(61750) := X"24420010";
        ram_buffer(61751) := X"AFC20068";
        ram_buffer(61752) := X"26310008";
        ram_buffer(61753) := X"8FC20064";
        ram_buffer(61754) := X"00000000";
        ram_buffer(61755) := X"24420001";
        ram_buffer(61756) := X"AFC20064";
        ram_buffer(61757) := X"8FC20064";
        ram_buffer(61758) := X"00000000";
        ram_buffer(61759) := X"28420008";
        ram_buffer(61760) := X"1440000A";
        ram_buffer(61761) := X"00000000";
        ram_buffer(61762) := X"27C20060";
        ram_buffer(61763) := X"00403021";
        ram_buffer(61764) := X"8FC50194";
        ram_buffer(61765) := X"8FC40190";
        ram_buffer(61766) := X"0C02EAF5";
        ram_buffer(61767) := X"00000000";
        ram_buffer(61768) := X"144000D2";
        ram_buffer(61769) := X"00000000";
        ram_buffer(61770) := X"27D1006C";
        ram_buffer(61771) := X"2610FFF0";
        ram_buffer(61772) := X"2A020011";
        ram_buffer(61773) := X"1040FFE1";
        ram_buffer(61774) := X"00000000";
        ram_buffer(61775) := X"3C02100D";
        ram_buffer(61776) := X"2442B280";
        ram_buffer(61777) := X"AE220000";
        ram_buffer(61778) := X"02001021";
        ram_buffer(61779) := X"AE220004";
        ram_buffer(61780) := X"8FC30068";
        ram_buffer(61781) := X"02001021";
        ram_buffer(61782) := X"00621021";
        ram_buffer(61783) := X"AFC20068";
        ram_buffer(61784) := X"26310008";
        ram_buffer(61785) := X"8FC20064";
        ram_buffer(61786) := X"00000000";
        ram_buffer(61787) := X"24420001";
        ram_buffer(61788) := X"AFC20064";
        ram_buffer(61789) := X"8FC20064";
        ram_buffer(61790) := X"00000000";
        ram_buffer(61791) := X"28420008";
        ram_buffer(61792) := X"1440000A";
        ram_buffer(61793) := X"00000000";
        ram_buffer(61794) := X"27C20060";
        ram_buffer(61795) := X"00403021";
        ram_buffer(61796) := X"8FC50194";
        ram_buffer(61797) := X"8FC40190";
        ram_buffer(61798) := X"0C02EAF5";
        ram_buffer(61799) := X"00000000";
        ram_buffer(61800) := X"144000B5";
        ram_buffer(61801) := X"00000000";
        ram_buffer(61802) := X"27D1006C";
        ram_buffer(61803) := X"AE330000";
        ram_buffer(61804) := X"8FC20044";
        ram_buffer(61805) := X"00000000";
        ram_buffer(61806) := X"AE220004";
        ram_buffer(61807) := X"8FC30068";
        ram_buffer(61808) := X"8FC20044";
        ram_buffer(61809) := X"00000000";
        ram_buffer(61810) := X"00621021";
        ram_buffer(61811) := X"AFC20068";
        ram_buffer(61812) := X"26310008";
        ram_buffer(61813) := X"8FC20064";
        ram_buffer(61814) := X"00000000";
        ram_buffer(61815) := X"24420001";
        ram_buffer(61816) := X"AFC20064";
        ram_buffer(61817) := X"8FC20064";
        ram_buffer(61818) := X"00000000";
        ram_buffer(61819) := X"28420008";
        ram_buffer(61820) := X"1440000A";
        ram_buffer(61821) := X"00000000";
        ram_buffer(61822) := X"27C20060";
        ram_buffer(61823) := X"00403021";
        ram_buffer(61824) := X"8FC50194";
        ram_buffer(61825) := X"8FC40190";
        ram_buffer(61826) := X"0C02EAF5";
        ram_buffer(61827) := X"00000000";
        ram_buffer(61828) := X"1440009C";
        ram_buffer(61829) := X"00000000";
        ram_buffer(61830) := X"27D1006C";
        ram_buffer(61831) := X"32420004";
        ram_buffer(61832) := X"10400045";
        ram_buffer(61833) := X"00000000";
        ram_buffer(61834) := X"8FC30014";
        ram_buffer(61835) := X"8FC20040";
        ram_buffer(61836) := X"00000000";
        ram_buffer(61837) := X"00628023";
        ram_buffer(61838) := X"1A00003F";
        ram_buffer(61839) := X"00000000";
        ram_buffer(61840) := X"1000001E";
        ram_buffer(61841) := X"00000000";
        ram_buffer(61842) := X"3C02100D";
        ram_buffer(61843) := X"2442B270";
        ram_buffer(61844) := X"AE220000";
        ram_buffer(61845) := X"24020010";
        ram_buffer(61846) := X"AE220004";
        ram_buffer(61847) := X"8FC20068";
        ram_buffer(61848) := X"00000000";
        ram_buffer(61849) := X"24420010";
        ram_buffer(61850) := X"AFC20068";
        ram_buffer(61851) := X"26310008";
        ram_buffer(61852) := X"8FC20064";
        ram_buffer(61853) := X"00000000";
        ram_buffer(61854) := X"24420001";
        ram_buffer(61855) := X"AFC20064";
        ram_buffer(61856) := X"8FC20064";
        ram_buffer(61857) := X"00000000";
        ram_buffer(61858) := X"28420008";
        ram_buffer(61859) := X"1440000A";
        ram_buffer(61860) := X"00000000";
        ram_buffer(61861) := X"27C20060";
        ram_buffer(61862) := X"00403021";
        ram_buffer(61863) := X"8FC50194";
        ram_buffer(61864) := X"8FC40190";
        ram_buffer(61865) := X"0C02EAF5";
        ram_buffer(61866) := X"00000000";
        ram_buffer(61867) := X"14400078";
        ram_buffer(61868) := X"00000000";
        ram_buffer(61869) := X"27D1006C";
        ram_buffer(61870) := X"2610FFF0";
        ram_buffer(61871) := X"2A020011";
        ram_buffer(61872) := X"1040FFE1";
        ram_buffer(61873) := X"00000000";
        ram_buffer(61874) := X"3C02100D";
        ram_buffer(61875) := X"2442B270";
        ram_buffer(61876) := X"AE220000";
        ram_buffer(61877) := X"02001021";
        ram_buffer(61878) := X"AE220004";
        ram_buffer(61879) := X"8FC20068";
        ram_buffer(61880) := X"02001821";
        ram_buffer(61881) := X"00431021";
        ram_buffer(61882) := X"AFC20068";
        ram_buffer(61883) := X"26310008";
        ram_buffer(61884) := X"8FC20064";
        ram_buffer(61885) := X"00000000";
        ram_buffer(61886) := X"24420001";
        ram_buffer(61887) := X"AFC20064";
        ram_buffer(61888) := X"8FC20064";
        ram_buffer(61889) := X"00000000";
        ram_buffer(61890) := X"28420008";
        ram_buffer(61891) := X"1440000A";
        ram_buffer(61892) := X"00000000";
        ram_buffer(61893) := X"27C20060";
        ram_buffer(61894) := X"00403021";
        ram_buffer(61895) := X"8FC50194";
        ram_buffer(61896) := X"8FC40190";
        ram_buffer(61897) := X"0C02EAF5";
        ram_buffer(61898) := X"00000000";
        ram_buffer(61899) := X"1440005B";
        ram_buffer(61900) := X"00000000";
        ram_buffer(61901) := X"27D1006C";
        ram_buffer(61902) := X"8FC30014";
        ram_buffer(61903) := X"8FC20040";
        ram_buffer(61904) := X"00000000";
        ram_buffer(61905) := X"0043202A";
        ram_buffer(61906) := X"10800002";
        ram_buffer(61907) := X"00000000";
        ram_buffer(61908) := X"00601021";
        ram_buffer(61909) := X"8FC30010";
        ram_buffer(61910) := X"00000000";
        ram_buffer(61911) := X"00621021";
        ram_buffer(61912) := X"AFC20010";
        ram_buffer(61913) := X"8FC20068";
        ram_buffer(61914) := X"00000000";
        ram_buffer(61915) := X"10400009";
        ram_buffer(61916) := X"00000000";
        ram_buffer(61917) := X"27C20060";
        ram_buffer(61918) := X"00403021";
        ram_buffer(61919) := X"8FC50194";
        ram_buffer(61920) := X"8FC40190";
        ram_buffer(61921) := X"0C02EAF5";
        ram_buffer(61922) := X"00000000";
        ram_buffer(61923) := X"14400046";
        ram_buffer(61924) := X"00000000";
        ram_buffer(61925) := X"AFC00064";
        ram_buffer(61926) := X"27D1006C";
        ram_buffer(61927) := X"8FC2004C";
        ram_buffer(61928) := X"00000000";
        ram_buffer(61929) := X"1040FA4E";
        ram_buffer(61930) := X"00000000";
        ram_buffer(61931) := X"8FC5004C";
        ram_buffer(61932) := X"8FC40190";
        ram_buffer(61933) := X"0C027301";
        ram_buffer(61934) := X"00000000";
        ram_buffer(61935) := X"AFC0004C";
        ram_buffer(61936) := X"1000FA47";
        ram_buffer(61937) := X"00000000";
        ram_buffer(61938) := X"00000000";
        ram_buffer(61939) := X"10000002";
        ram_buffer(61940) := X"00000000";
        ram_buffer(61941) := X"00000000";
        ram_buffer(61942) := X"8FC20068";
        ram_buffer(61943) := X"00000000";
        ram_buffer(61944) := X"10400009";
        ram_buffer(61945) := X"00000000";
        ram_buffer(61946) := X"27C20060";
        ram_buffer(61947) := X"00403021";
        ram_buffer(61948) := X"8FC50194";
        ram_buffer(61949) := X"8FC40190";
        ram_buffer(61950) := X"0C02EAF5";
        ram_buffer(61951) := X"00000000";
        ram_buffer(61952) := X"1440002C";
        ram_buffer(61953) := X"00000000";
        ram_buffer(61954) := X"AFC00064";
        ram_buffer(61955) := X"27D1006C";
        ram_buffer(61956) := X"10000029";
        ram_buffer(61957) := X"00000000";
        ram_buffer(61958) := X"00000000";
        ram_buffer(61959) := X"10000026";
        ram_buffer(61960) := X"00000000";
        ram_buffer(61961) := X"00000000";
        ram_buffer(61962) := X"10000023";
        ram_buffer(61963) := X"00000000";
        ram_buffer(61964) := X"00000000";
        ram_buffer(61965) := X"10000020";
        ram_buffer(61966) := X"00000000";
        ram_buffer(61967) := X"00000000";
        ram_buffer(61968) := X"1000001D";
        ram_buffer(61969) := X"00000000";
        ram_buffer(61970) := X"00000000";
        ram_buffer(61971) := X"1000001A";
        ram_buffer(61972) := X"00000000";
        ram_buffer(61973) := X"00000000";
        ram_buffer(61974) := X"10000017";
        ram_buffer(61975) := X"00000000";
        ram_buffer(61976) := X"00000000";
        ram_buffer(61977) := X"10000014";
        ram_buffer(61978) := X"00000000";
        ram_buffer(61979) := X"00000000";
        ram_buffer(61980) := X"10000011";
        ram_buffer(61981) := X"00000000";
        ram_buffer(61982) := X"00000000";
        ram_buffer(61983) := X"1000000E";
        ram_buffer(61984) := X"00000000";
        ram_buffer(61985) := X"00000000";
        ram_buffer(61986) := X"1000000B";
        ram_buffer(61987) := X"00000000";
        ram_buffer(61988) := X"00000000";
        ram_buffer(61989) := X"10000008";
        ram_buffer(61990) := X"00000000";
        ram_buffer(61991) := X"00000000";
        ram_buffer(61992) := X"10000005";
        ram_buffer(61993) := X"00000000";
        ram_buffer(61994) := X"00000000";
        ram_buffer(61995) := X"10000002";
        ram_buffer(61996) := X"00000000";
        ram_buffer(61997) := X"00000000";
        ram_buffer(61998) := X"8FC2004C";
        ram_buffer(61999) := X"00000000";
        ram_buffer(62000) := X"10400005";
        ram_buffer(62001) := X"00000000";
        ram_buffer(62002) := X"8FC5004C";
        ram_buffer(62003) := X"8FC40190";
        ram_buffer(62004) := X"0C027301";
        ram_buffer(62005) := X"00000000";
        ram_buffer(62006) := X"8FC20194";
        ram_buffer(62007) := X"00000000";
        ram_buffer(62008) := X"8442000C";
        ram_buffer(62009) := X"00000000";
        ram_buffer(62010) := X"3042FFFF";
        ram_buffer(62011) := X"30420040";
        ram_buffer(62012) := X"14400004";
        ram_buffer(62013) := X"00000000";
        ram_buffer(62014) := X"8FC20010";
        ram_buffer(62015) := X"10000003";
        ram_buffer(62016) := X"00000000";
        ram_buffer(62017) := X"2402FFFF";
        ram_buffer(62018) := X"00000000";
        ram_buffer(62019) := X"03C0E821";
        ram_buffer(62020) := X"8FBF018C";
        ram_buffer(62021) := X"8FBE0188";
        ram_buffer(62022) := X"8FB70184";
        ram_buffer(62023) := X"8FB60180";
        ram_buffer(62024) := X"8FB5017C";
        ram_buffer(62025) := X"8FB40178";
        ram_buffer(62026) := X"8FB30174";
        ram_buffer(62027) := X"8FB20170";
        ram_buffer(62028) := X"8FB1016C";
        ram_buffer(62029) := X"8FB00168";
        ram_buffer(62030) := X"27BD0190";
        ram_buffer(62031) := X"03E00008";
        ram_buffer(62032) := X"00000000";
        ram_buffer(62033) := X"27BDFFD0";
        ram_buffer(62034) := X"AFBF002C";
        ram_buffer(62035) := X"AFBE0028";
        ram_buffer(62036) := X"03A0F021";
        ram_buffer(62037) := X"AFC40030";
        ram_buffer(62038) := X"AFC50034";
        ram_buffer(62039) := X"AFC60038";
        ram_buffer(62040) := X"8FC30034";
        ram_buffer(62041) := X"8FC20038";
        ram_buffer(62042) := X"00000000";
        ram_buffer(62043) := X"00620018";
        ram_buffer(62044) := X"00001012";
        ram_buffer(62045) := X"AFC20014";
        ram_buffer(62046) := X"8FC50014";
        ram_buffer(62047) := X"8FC40030";
        ram_buffer(62048) := X"0C027B8F";
        ram_buffer(62049) := X"00000000";
        ram_buffer(62050) := X"AFC20018";
        ram_buffer(62051) := X"8FC20018";
        ram_buffer(62052) := X"00000000";
        ram_buffer(62053) := X"14400004";
        ram_buffer(62054) := X"00000000";
        ram_buffer(62055) := X"00001021";
        ram_buffer(62056) := X"10000059";
        ram_buffer(62057) := X"00000000";
        ram_buffer(62058) := X"8FC20018";
        ram_buffer(62059) := X"00000000";
        ram_buffer(62060) := X"2442FFF8";
        ram_buffer(62061) := X"AFC2001C";
        ram_buffer(62062) := X"8FC2001C";
        ram_buffer(62063) := X"00000000";
        ram_buffer(62064) := X"8C430004";
        ram_buffer(62065) := X"2402FFFC";
        ram_buffer(62066) := X"00621024";
        ram_buffer(62067) := X"AFC20020";
        ram_buffer(62068) := X"8FC20020";
        ram_buffer(62069) := X"00000000";
        ram_buffer(62070) := X"2442FFFC";
        ram_buffer(62071) := X"AFC20024";
        ram_buffer(62072) := X"8FC20024";
        ram_buffer(62073) := X"00000000";
        ram_buffer(62074) := X"2C420025";
        ram_buffer(62075) := X"10400040";
        ram_buffer(62076) := X"00000000";
        ram_buffer(62077) := X"8FC20018";
        ram_buffer(62078) := X"00000000";
        ram_buffer(62079) := X"AFC20010";
        ram_buffer(62080) := X"8FC20024";
        ram_buffer(62081) := X"00000000";
        ram_buffer(62082) := X"2C420014";
        ram_buffer(62083) := X"14400029";
        ram_buffer(62084) := X"00000000";
        ram_buffer(62085) := X"8FC20010";
        ram_buffer(62086) := X"00000000";
        ram_buffer(62087) := X"24430004";
        ram_buffer(62088) := X"AFC30010";
        ram_buffer(62089) := X"AC400000";
        ram_buffer(62090) := X"8FC20010";
        ram_buffer(62091) := X"00000000";
        ram_buffer(62092) := X"24430004";
        ram_buffer(62093) := X"AFC30010";
        ram_buffer(62094) := X"AC400000";
        ram_buffer(62095) := X"8FC20024";
        ram_buffer(62096) := X"00000000";
        ram_buffer(62097) := X"2C42001C";
        ram_buffer(62098) := X"1440001A";
        ram_buffer(62099) := X"00000000";
        ram_buffer(62100) := X"8FC20010";
        ram_buffer(62101) := X"00000000";
        ram_buffer(62102) := X"24430004";
        ram_buffer(62103) := X"AFC30010";
        ram_buffer(62104) := X"AC400000";
        ram_buffer(62105) := X"8FC20010";
        ram_buffer(62106) := X"00000000";
        ram_buffer(62107) := X"24430004";
        ram_buffer(62108) := X"AFC30010";
        ram_buffer(62109) := X"AC400000";
        ram_buffer(62110) := X"8FC20024";
        ram_buffer(62111) := X"00000000";
        ram_buffer(62112) := X"2C420024";
        ram_buffer(62113) := X"1440000B";
        ram_buffer(62114) := X"00000000";
        ram_buffer(62115) := X"8FC20010";
        ram_buffer(62116) := X"00000000";
        ram_buffer(62117) := X"24430004";
        ram_buffer(62118) := X"AFC30010";
        ram_buffer(62119) := X"AC400000";
        ram_buffer(62120) := X"8FC20010";
        ram_buffer(62121) := X"00000000";
        ram_buffer(62122) := X"24430004";
        ram_buffer(62123) := X"AFC30010";
        ram_buffer(62124) := X"AC400000";
        ram_buffer(62125) := X"8FC20010";
        ram_buffer(62126) := X"00000000";
        ram_buffer(62127) := X"24430004";
        ram_buffer(62128) := X"AFC30010";
        ram_buffer(62129) := X"AC400000";
        ram_buffer(62130) := X"8FC20010";
        ram_buffer(62131) := X"00000000";
        ram_buffer(62132) := X"24430004";
        ram_buffer(62133) := X"AFC30010";
        ram_buffer(62134) := X"AC400000";
        ram_buffer(62135) := X"8FC20010";
        ram_buffer(62136) := X"00000000";
        ram_buffer(62137) := X"AC400000";
        ram_buffer(62138) := X"10000006";
        ram_buffer(62139) := X"00000000";
        ram_buffer(62140) := X"8FC60024";
        ram_buffer(62141) := X"00002821";
        ram_buffer(62142) := X"8FC40018";
        ram_buffer(62143) := X"0C02801D";
        ram_buffer(62144) := X"00000000";
        ram_buffer(62145) := X"8FC20018";
        ram_buffer(62146) := X"03C0E821";
        ram_buffer(62147) := X"8FBF002C";
        ram_buffer(62148) := X"8FBE0028";
        ram_buffer(62149) := X"27BD0030";
        ram_buffer(62150) := X"03E00008";
        ram_buffer(62151) := X"00000000";
        ram_buffer(62152) := X"27BDFFD8";
        ram_buffer(62153) := X"AFBF0024";
        ram_buffer(62154) := X"AFBE0020";
        ram_buffer(62155) := X"03A0F021";
        ram_buffer(62156) := X"AFC40028";
        ram_buffer(62157) := X"AFC5002C";
        ram_buffer(62158) := X"AFC60030";
        ram_buffer(62159) := X"0C02BB09";
        ram_buffer(62160) := X"00000000";
        ram_buffer(62161) := X"00401821";
        ram_buffer(62162) := X"24020001";
        ram_buffer(62163) := X"14620013";
        ram_buffer(62164) := X"00000000";
        ram_buffer(62165) := X"8FC2002C";
        ram_buffer(62166) := X"00000000";
        ram_buffer(62167) := X"1840000F";
        ram_buffer(62168) := X"00000000";
        ram_buffer(62169) := X"8FC2002C";
        ram_buffer(62170) := X"00000000";
        ram_buffer(62171) := X"28420100";
        ram_buffer(62172) := X"1040000A";
        ram_buffer(62173) := X"00000000";
        ram_buffer(62174) := X"8FC2002C";
        ram_buffer(62175) := X"00000000";
        ram_buffer(62176) := X"00021600";
        ram_buffer(62177) := X"00021603";
        ram_buffer(62178) := X"A3C20018";
        ram_buffer(62179) := X"24020001";
        ram_buffer(62180) := X"AFC20014";
        ram_buffer(62181) := X"1000001D";
        ram_buffer(62182) := X"00000000";
        ram_buffer(62183) := X"8FC20030";
        ram_buffer(62184) := X"00000000";
        ram_buffer(62185) := X"2443005C";
        ram_buffer(62186) := X"27C20018";
        ram_buffer(62187) := X"00603821";
        ram_buffer(62188) := X"8FC6002C";
        ram_buffer(62189) := X"00402821";
        ram_buffer(62190) := X"8FC40028";
        ram_buffer(62191) := X"0C02FA96";
        ram_buffer(62192) := X"00000000";
        ram_buffer(62193) := X"AFC20014";
        ram_buffer(62194) := X"8FC30014";
        ram_buffer(62195) := X"2402FFFF";
        ram_buffer(62196) := X"1462000E";
        ram_buffer(62197) := X"00000000";
        ram_buffer(62198) := X"8FC20030";
        ram_buffer(62199) := X"00000000";
        ram_buffer(62200) := X"8442000C";
        ram_buffer(62201) := X"00000000";
        ram_buffer(62202) := X"34420040";
        ram_buffer(62203) := X"00021C00";
        ram_buffer(62204) := X"00031C03";
        ram_buffer(62205) := X"8FC20030";
        ram_buffer(62206) := X"00000000";
        ram_buffer(62207) := X"A443000C";
        ram_buffer(62208) := X"2402FFFF";
        ram_buffer(62209) := X"1000007E";
        ram_buffer(62210) := X"00000000";
        ram_buffer(62211) := X"AFC00010";
        ram_buffer(62212) := X"10000074";
        ram_buffer(62213) := X"00000000";
        ram_buffer(62214) := X"8FC20030";
        ram_buffer(62215) := X"00000000";
        ram_buffer(62216) := X"8C420008";
        ram_buffer(62217) := X"00000000";
        ram_buffer(62218) := X"2443FFFF";
        ram_buffer(62219) := X"8FC20030";
        ram_buffer(62220) := X"00000000";
        ram_buffer(62221) := X"AC430008";
        ram_buffer(62222) := X"8FC20030";
        ram_buffer(62223) := X"00000000";
        ram_buffer(62224) := X"8C420008";
        ram_buffer(62225) := X"00000000";
        ram_buffer(62226) := X"04410046";
        ram_buffer(62227) := X"00000000";
        ram_buffer(62228) := X"8FC20030";
        ram_buffer(62229) := X"00000000";
        ram_buffer(62230) := X"8C430008";
        ram_buffer(62231) := X"8FC20030";
        ram_buffer(62232) := X"00000000";
        ram_buffer(62233) := X"8C420018";
        ram_buffer(62234) := X"00000000";
        ram_buffer(62235) := X"0062102A";
        ram_buffer(62236) := X"1440002C";
        ram_buffer(62237) := X"00000000";
        ram_buffer(62238) := X"8FC20030";
        ram_buffer(62239) := X"00000000";
        ram_buffer(62240) := X"8C420000";
        ram_buffer(62241) := X"8FC30010";
        ram_buffer(62242) := X"27C40010";
        ram_buffer(62243) := X"00831821";
        ram_buffer(62244) := X"80630008";
        ram_buffer(62245) := X"00000000";
        ram_buffer(62246) := X"306300FF";
        ram_buffer(62247) := X"A0430000";
        ram_buffer(62248) := X"8FC20030";
        ram_buffer(62249) := X"00000000";
        ram_buffer(62250) := X"8C420000";
        ram_buffer(62251) := X"00000000";
        ram_buffer(62252) := X"90430000";
        ram_buffer(62253) := X"2402000A";
        ram_buffer(62254) := X"10620010";
        ram_buffer(62255) := X"00000000";
        ram_buffer(62256) := X"8FC20030";
        ram_buffer(62257) := X"00000000";
        ram_buffer(62258) := X"8C420000";
        ram_buffer(62259) := X"00000000";
        ram_buffer(62260) := X"24440001";
        ram_buffer(62261) := X"8FC30030";
        ram_buffer(62262) := X"00000000";
        ram_buffer(62263) := X"AC640000";
        ram_buffer(62264) := X"90420000";
        ram_buffer(62265) := X"00000000";
        ram_buffer(62266) := X"24420001";
        ram_buffer(62267) := X"2C420001";
        ram_buffer(62268) := X"304200FF";
        ram_buffer(62269) := X"10000032";
        ram_buffer(62270) := X"00000000";
        ram_buffer(62271) := X"8FC60030";
        ram_buffer(62272) := X"2405000A";
        ram_buffer(62273) := X"8FC40028";
        ram_buffer(62274) := X"0C02FA03";
        ram_buffer(62275) := X"00000000";
        ram_buffer(62276) := X"24420001";
        ram_buffer(62277) := X"2C420001";
        ram_buffer(62278) := X"304200FF";
        ram_buffer(62279) := X"10000028";
        ram_buffer(62280) := X"00000000";
        ram_buffer(62281) := X"8FC20010";
        ram_buffer(62282) := X"27C30010";
        ram_buffer(62283) := X"00621021";
        ram_buffer(62284) := X"80420008";
        ram_buffer(62285) := X"00000000";
        ram_buffer(62286) := X"304200FF";
        ram_buffer(62287) := X"8FC60030";
        ram_buffer(62288) := X"00402821";
        ram_buffer(62289) := X"8FC40028";
        ram_buffer(62290) := X"0C02FA03";
        ram_buffer(62291) := X"00000000";
        ram_buffer(62292) := X"24420001";
        ram_buffer(62293) := X"2C420001";
        ram_buffer(62294) := X"304200FF";
        ram_buffer(62295) := X"10000018";
        ram_buffer(62296) := X"00000000";
        ram_buffer(62297) := X"8FC20030";
        ram_buffer(62298) := X"00000000";
        ram_buffer(62299) := X"8C420000";
        ram_buffer(62300) := X"8FC30010";
        ram_buffer(62301) := X"27C40010";
        ram_buffer(62302) := X"00831821";
        ram_buffer(62303) := X"80630008";
        ram_buffer(62304) := X"00000000";
        ram_buffer(62305) := X"306300FF";
        ram_buffer(62306) := X"A0430000";
        ram_buffer(62307) := X"8FC20030";
        ram_buffer(62308) := X"00000000";
        ram_buffer(62309) := X"8C420000";
        ram_buffer(62310) := X"00000000";
        ram_buffer(62311) := X"24440001";
        ram_buffer(62312) := X"8FC30030";
        ram_buffer(62313) := X"00000000";
        ram_buffer(62314) := X"AC640000";
        ram_buffer(62315) := X"90420000";
        ram_buffer(62316) := X"00000000";
        ram_buffer(62317) := X"24420001";
        ram_buffer(62318) := X"2C420001";
        ram_buffer(62319) := X"304200FF";
        ram_buffer(62320) := X"10400004";
        ram_buffer(62321) := X"00000000";
        ram_buffer(62322) := X"2402FFFF";
        ram_buffer(62323) := X"1000000C";
        ram_buffer(62324) := X"00000000";
        ram_buffer(62325) := X"8FC20010";
        ram_buffer(62326) := X"00000000";
        ram_buffer(62327) := X"24420001";
        ram_buffer(62328) := X"AFC20010";
        ram_buffer(62329) := X"8FC30010";
        ram_buffer(62330) := X"8FC20014";
        ram_buffer(62331) := X"00000000";
        ram_buffer(62332) := X"0062102B";
        ram_buffer(62333) := X"1440FF88";
        ram_buffer(62334) := X"00000000";
        ram_buffer(62335) := X"8FC2002C";
        ram_buffer(62336) := X"03C0E821";
        ram_buffer(62337) := X"8FBF0024";
        ram_buffer(62338) := X"8FBE0020";
        ram_buffer(62339) := X"27BD0028";
        ram_buffer(62340) := X"03E00008";
        ram_buffer(62341) := X"00000000";
        ram_buffer(62342) := X"27BDFFE0";
        ram_buffer(62343) := X"AFBF001C";
        ram_buffer(62344) := X"AFBE0018";
        ram_buffer(62345) := X"03A0F021";
        ram_buffer(62346) := X"AFC40020";
        ram_buffer(62347) := X"AFC50024";
        ram_buffer(62348) := X"AFC60028";
        ram_buffer(62349) := X"8FC20028";
        ram_buffer(62350) := X"00000000";
        ram_buffer(62351) := X"8442000C";
        ram_buffer(62352) := X"00000000";
        ram_buffer(62353) := X"3042FFFF";
        ram_buffer(62354) := X"30422000";
        ram_buffer(62355) := X"14400013";
        ram_buffer(62356) := X"00000000";
        ram_buffer(62357) := X"8FC20028";
        ram_buffer(62358) := X"00000000";
        ram_buffer(62359) := X"8442000C";
        ram_buffer(62360) := X"00000000";
        ram_buffer(62361) := X"34422000";
        ram_buffer(62362) := X"00021C00";
        ram_buffer(62363) := X"00031C03";
        ram_buffer(62364) := X"8FC20028";
        ram_buffer(62365) := X"00000000";
        ram_buffer(62366) := X"A443000C";
        ram_buffer(62367) := X"8FC20028";
        ram_buffer(62368) := X"00000000";
        ram_buffer(62369) := X"8C420064";
        ram_buffer(62370) := X"00000000";
        ram_buffer(62371) := X"34432000";
        ram_buffer(62372) := X"8FC20028";
        ram_buffer(62373) := X"00000000";
        ram_buffer(62374) := X"AC430064";
        ram_buffer(62375) := X"8FC60028";
        ram_buffer(62376) := X"8FC50024";
        ram_buffer(62377) := X"8FC40020";
        ram_buffer(62378) := X"0C02F2C8";
        ram_buffer(62379) := X"00000000";
        ram_buffer(62380) := X"AFC20010";
        ram_buffer(62381) := X"8FC20010";
        ram_buffer(62382) := X"03C0E821";
        ram_buffer(62383) := X"8FBF001C";
        ram_buffer(62384) := X"8FBE0018";
        ram_buffer(62385) := X"27BD0020";
        ram_buffer(62386) := X"03E00008";
        ram_buffer(62387) := X"00000000";
        ram_buffer(62388) := X"27BDFFE0";
        ram_buffer(62389) := X"AFBF001C";
        ram_buffer(62390) := X"AFBE0018";
        ram_buffer(62391) := X"03A0F021";
        ram_buffer(62392) := X"AFC40020";
        ram_buffer(62393) := X"AFC50024";
        ram_buffer(62394) := X"8F828098";
        ram_buffer(62395) := X"00000000";
        ram_buffer(62396) := X"AFC20010";
        ram_buffer(62397) := X"8FC20010";
        ram_buffer(62398) := X"00000000";
        ram_buffer(62399) := X"AFC20014";
        ram_buffer(62400) := X"8FC20014";
        ram_buffer(62401) := X"00000000";
        ram_buffer(62402) := X"1040000A";
        ram_buffer(62403) := X"00000000";
        ram_buffer(62404) := X"8FC20014";
        ram_buffer(62405) := X"00000000";
        ram_buffer(62406) := X"8C420038";
        ram_buffer(62407) := X"00000000";
        ram_buffer(62408) := X"14400004";
        ram_buffer(62409) := X"00000000";
        ram_buffer(62410) := X"8FC40014";
        ram_buffer(62411) := X"0C027069";
        ram_buffer(62412) := X"00000000";
        ram_buffer(62413) := X"8FC60024";
        ram_buffer(62414) := X"8FC50020";
        ram_buffer(62415) := X"8FC40010";
        ram_buffer(62416) := X"0C02F386";
        ram_buffer(62417) := X"00000000";
        ram_buffer(62418) := X"03C0E821";
        ram_buffer(62419) := X"8FBF001C";
        ram_buffer(62420) := X"8FBE0018";
        ram_buffer(62421) := X"27BD0020";
        ram_buffer(62422) := X"03E00008";
        ram_buffer(62423) := X"00000000";
        ram_buffer(62424) := X"27BDFFE0";
        ram_buffer(62425) := X"AFBE001C";
        ram_buffer(62426) := X"03A0F021";
        ram_buffer(62427) := X"AFC40020";
        ram_buffer(62428) := X"AFC50024";
        ram_buffer(62429) := X"8FC20020";
        ram_buffer(62430) := X"00000000";
        ram_buffer(62431) := X"24420014";
        ram_buffer(62432) := X"AFC20004";
        ram_buffer(62433) := X"8FC20004";
        ram_buffer(62434) := X"00000000";
        ram_buffer(62435) := X"AFC20000";
        ram_buffer(62436) := X"8FC20024";
        ram_buffer(62437) := X"00000000";
        ram_buffer(62438) := X"00021143";
        ram_buffer(62439) := X"AFC2000C";
        ram_buffer(62440) := X"8FC20020";
        ram_buffer(62441) := X"00000000";
        ram_buffer(62442) := X"8C430010";
        ram_buffer(62443) := X"8FC2000C";
        ram_buffer(62444) := X"00000000";
        ram_buffer(62445) := X"0043102A";
        ram_buffer(62446) := X"10400067";
        ram_buffer(62447) := X"00000000";
        ram_buffer(62448) := X"8FC20020";
        ram_buffer(62449) := X"00000000";
        ram_buffer(62450) := X"8C420010";
        ram_buffer(62451) := X"00000000";
        ram_buffer(62452) := X"00021080";
        ram_buffer(62453) := X"8FC30000";
        ram_buffer(62454) := X"00000000";
        ram_buffer(62455) := X"00621021";
        ram_buffer(62456) := X"AFC20010";
        ram_buffer(62457) := X"8FC2000C";
        ram_buffer(62458) := X"00000000";
        ram_buffer(62459) := X"00021080";
        ram_buffer(62460) := X"8FC30000";
        ram_buffer(62461) := X"00000000";
        ram_buffer(62462) := X"00621021";
        ram_buffer(62463) := X"AFC20000";
        ram_buffer(62464) := X"8FC20024";
        ram_buffer(62465) := X"00000000";
        ram_buffer(62466) := X"3042001F";
        ram_buffer(62467) := X"AFC20024";
        ram_buffer(62468) := X"8FC20024";
        ram_buffer(62469) := X"00000000";
        ram_buffer(62470) := X"10400049";
        ram_buffer(62471) := X"00000000";
        ram_buffer(62472) := X"24030020";
        ram_buffer(62473) := X"8FC20024";
        ram_buffer(62474) := X"00000000";
        ram_buffer(62475) := X"00621023";
        ram_buffer(62476) := X"AFC2000C";
        ram_buffer(62477) := X"8FC20000";
        ram_buffer(62478) := X"00000000";
        ram_buffer(62479) := X"24430004";
        ram_buffer(62480) := X"AFC30000";
        ram_buffer(62481) := X"8C430000";
        ram_buffer(62482) := X"8FC20024";
        ram_buffer(62483) := X"00000000";
        ram_buffer(62484) := X"00431006";
        ram_buffer(62485) := X"AFC20008";
        ram_buffer(62486) := X"10000018";
        ram_buffer(62487) := X"00000000";
        ram_buffer(62488) := X"8FC20004";
        ram_buffer(62489) := X"00000000";
        ram_buffer(62490) := X"24430004";
        ram_buffer(62491) := X"AFC30004";
        ram_buffer(62492) := X"8FC30000";
        ram_buffer(62493) := X"00000000";
        ram_buffer(62494) := X"8C640000";
        ram_buffer(62495) := X"8FC3000C";
        ram_buffer(62496) := X"00000000";
        ram_buffer(62497) := X"00642004";
        ram_buffer(62498) := X"8FC30008";
        ram_buffer(62499) := X"00000000";
        ram_buffer(62500) := X"00831825";
        ram_buffer(62501) := X"AC430000";
        ram_buffer(62502) := X"8FC20000";
        ram_buffer(62503) := X"00000000";
        ram_buffer(62504) := X"24430004";
        ram_buffer(62505) := X"AFC30000";
        ram_buffer(62506) := X"8C430000";
        ram_buffer(62507) := X"8FC20024";
        ram_buffer(62508) := X"00000000";
        ram_buffer(62509) := X"00431006";
        ram_buffer(62510) := X"AFC20008";
        ram_buffer(62511) := X"8FC30000";
        ram_buffer(62512) := X"8FC20010";
        ram_buffer(62513) := X"00000000";
        ram_buffer(62514) := X"0062102B";
        ram_buffer(62515) := X"1440FFE4";
        ram_buffer(62516) := X"00000000";
        ram_buffer(62517) := X"8FC20004";
        ram_buffer(62518) := X"8FC30008";
        ram_buffer(62519) := X"00000000";
        ram_buffer(62520) := X"AC430000";
        ram_buffer(62521) := X"8FC20004";
        ram_buffer(62522) := X"00000000";
        ram_buffer(62523) := X"8C420000";
        ram_buffer(62524) := X"00000000";
        ram_buffer(62525) := X"10400018";
        ram_buffer(62526) := X"00000000";
        ram_buffer(62527) := X"8FC20004";
        ram_buffer(62528) := X"00000000";
        ram_buffer(62529) := X"24420004";
        ram_buffer(62530) := X"AFC20004";
        ram_buffer(62531) := X"10000012";
        ram_buffer(62532) := X"00000000";
        ram_buffer(62533) := X"8FC20004";
        ram_buffer(62534) := X"00000000";
        ram_buffer(62535) := X"24430004";
        ram_buffer(62536) := X"AFC30004";
        ram_buffer(62537) := X"8FC30000";
        ram_buffer(62538) := X"00000000";
        ram_buffer(62539) := X"24640004";
        ram_buffer(62540) := X"AFC40000";
        ram_buffer(62541) := X"8C630000";
        ram_buffer(62542) := X"00000000";
        ram_buffer(62543) := X"AC430000";
        ram_buffer(62544) := X"8FC30000";
        ram_buffer(62545) := X"8FC20010";
        ram_buffer(62546) := X"00000000";
        ram_buffer(62547) := X"0062102B";
        ram_buffer(62548) := X"1440FFF0";
        ram_buffer(62549) := X"00000000";
        ram_buffer(62550) := X"8FC20004";
        ram_buffer(62551) := X"8FC30020";
        ram_buffer(62552) := X"00000000";
        ram_buffer(62553) := X"24630014";
        ram_buffer(62554) := X"00431023";
        ram_buffer(62555) := X"00021083";
        ram_buffer(62556) := X"00401821";
        ram_buffer(62557) := X"8FC20020";
        ram_buffer(62558) := X"00000000";
        ram_buffer(62559) := X"AC430010";
        ram_buffer(62560) := X"8FC20020";
        ram_buffer(62561) := X"00000000";
        ram_buffer(62562) := X"8C420010";
        ram_buffer(62563) := X"00000000";
        ram_buffer(62564) := X"14400004";
        ram_buffer(62565) := X"00000000";
        ram_buffer(62566) := X"8FC20020";
        ram_buffer(62567) := X"00000000";
        ram_buffer(62568) := X"AC400014";
        ram_buffer(62569) := X"00000000";
        ram_buffer(62570) := X"03C0E821";
        ram_buffer(62571) := X"8FBE001C";
        ram_buffer(62572) := X"27BD0020";
        ram_buffer(62573) := X"03E00008";
        ram_buffer(62574) := X"00000000";
        ram_buffer(62575) := X"27BDFFD8";
        ram_buffer(62576) := X"AFBF0024";
        ram_buffer(62577) := X"AFBE0020";
        ram_buffer(62578) := X"03A0F021";
        ram_buffer(62579) := X"AFC40028";
        ram_buffer(62580) := X"AFC5002C";
        ram_buffer(62581) := X"8FC2002C";
        ram_buffer(62582) := X"00000000";
        ram_buffer(62583) := X"24420014";
        ram_buffer(62584) := X"AFC20010";
        ram_buffer(62585) := X"8FC2002C";
        ram_buffer(62586) := X"00000000";
        ram_buffer(62587) := X"8C420010";
        ram_buffer(62588) := X"00000000";
        ram_buffer(62589) := X"00021080";
        ram_buffer(62590) := X"8FC30010";
        ram_buffer(62591) := X"00000000";
        ram_buffer(62592) := X"00621021";
        ram_buffer(62593) := X"AFC20014";
        ram_buffer(62594) := X"8FC20010";
        ram_buffer(62595) := X"00000000";
        ram_buffer(62596) := X"8C430000";
        ram_buffer(62597) := X"2402FFFF";
        ram_buffer(62598) := X"1062000C";
        ram_buffer(62599) := X"00000000";
        ram_buffer(62600) := X"8FC20010";
        ram_buffer(62601) := X"00000000";
        ram_buffer(62602) := X"8C420000";
        ram_buffer(62603) := X"00000000";
        ram_buffer(62604) := X"24430001";
        ram_buffer(62605) := X"8FC20010";
        ram_buffer(62606) := X"00000000";
        ram_buffer(62607) := X"AC430000";
        ram_buffer(62608) := X"8FC2002C";
        ram_buffer(62609) := X"10000047";
        ram_buffer(62610) := X"00000000";
        ram_buffer(62611) := X"8FC20010";
        ram_buffer(62612) := X"00000000";
        ram_buffer(62613) := X"24430004";
        ram_buffer(62614) := X"AFC30010";
        ram_buffer(62615) := X"AC400000";
        ram_buffer(62616) := X"8FC30010";
        ram_buffer(62617) := X"8FC20014";
        ram_buffer(62618) := X"00000000";
        ram_buffer(62619) := X"0062102B";
        ram_buffer(62620) := X"1440FFE5";
        ram_buffer(62621) := X"00000000";
        ram_buffer(62622) := X"8FC2002C";
        ram_buffer(62623) := X"00000000";
        ram_buffer(62624) := X"8C430010";
        ram_buffer(62625) := X"8FC2002C";
        ram_buffer(62626) := X"00000000";
        ram_buffer(62627) := X"8C420008";
        ram_buffer(62628) := X"00000000";
        ram_buffer(62629) := X"0062102A";
        ram_buffer(62630) := X"14400023";
        ram_buffer(62631) := X"00000000";
        ram_buffer(62632) := X"8FC2002C";
        ram_buffer(62633) := X"00000000";
        ram_buffer(62634) := X"8C420004";
        ram_buffer(62635) := X"00000000";
        ram_buffer(62636) := X"24420001";
        ram_buffer(62637) := X"00402821";
        ram_buffer(62638) := X"8FC40028";
        ram_buffer(62639) := X"0C02BDA8";
        ram_buffer(62640) := X"00000000";
        ram_buffer(62641) := X"AFC20018";
        ram_buffer(62642) := X"8FC20018";
        ram_buffer(62643) := X"00000000";
        ram_buffer(62644) := X"2443000C";
        ram_buffer(62645) := X"8FC2002C";
        ram_buffer(62646) := X"00000000";
        ram_buffer(62647) := X"2444000C";
        ram_buffer(62648) := X"8FC2002C";
        ram_buffer(62649) := X"00000000";
        ram_buffer(62650) := X"8C420010";
        ram_buffer(62651) := X"00000000";
        ram_buffer(62652) := X"24420002";
        ram_buffer(62653) := X"00021080";
        ram_buffer(62654) := X"00403021";
        ram_buffer(62655) := X"00802821";
        ram_buffer(62656) := X"00602021";
        ram_buffer(62657) := X"0C027F93";
        ram_buffer(62658) := X"00000000";
        ram_buffer(62659) := X"8FC5002C";
        ram_buffer(62660) := X"8FC40028";
        ram_buffer(62661) := X"0C02BE10";
        ram_buffer(62662) := X"00000000";
        ram_buffer(62663) := X"8FC20018";
        ram_buffer(62664) := X"00000000";
        ram_buffer(62665) := X"AFC2002C";
        ram_buffer(62666) := X"8FC2002C";
        ram_buffer(62667) := X"00000000";
        ram_buffer(62668) := X"8C420010";
        ram_buffer(62669) := X"00000000";
        ram_buffer(62670) := X"24440001";
        ram_buffer(62671) := X"8FC3002C";
        ram_buffer(62672) := X"00000000";
        ram_buffer(62673) := X"AC640010";
        ram_buffer(62674) := X"8FC3002C";
        ram_buffer(62675) := X"24420004";
        ram_buffer(62676) := X"00021080";
        ram_buffer(62677) := X"00621021";
        ram_buffer(62678) := X"24030001";
        ram_buffer(62679) := X"AC430004";
        ram_buffer(62680) := X"8FC2002C";
        ram_buffer(62681) := X"03C0E821";
        ram_buffer(62682) := X"8FBF0024";
        ram_buffer(62683) := X"8FBE0020";
        ram_buffer(62684) := X"27BD0028";
        ram_buffer(62685) := X"03E00008";
        ram_buffer(62686) := X"00000000";
        ram_buffer(62687) := X"27BDFF88";
        ram_buffer(62688) := X"AFBF0074";
        ram_buffer(62689) := X"AFBE0070";
        ram_buffer(62690) := X"AFB0006C";
        ram_buffer(62691) := X"03A0F021";
        ram_buffer(62692) := X"AFC40078";
        ram_buffer(62693) := X"AFC5007C";
        ram_buffer(62694) := X"AFC60080";
        ram_buffer(62695) := X"AFC70084";
        ram_buffer(62696) := X"8FC40078";
        ram_buffer(62697) := X"0C02BB25";
        ram_buffer(62698) := X"00000000";
        ram_buffer(62699) := X"8C420000";
        ram_buffer(62700) := X"00000000";
        ram_buffer(62701) := X"AFC20058";
        ram_buffer(62702) := X"8FC40058";
        ram_buffer(62703) := X"0C02851E";
        ram_buffer(62704) := X"00000000";
        ram_buffer(62705) := X"AFC2005C";
        ram_buffer(62706) := X"8FC2005C";
        ram_buffer(62707) := X"00000000";
        ram_buffer(62708) := X"2442FFFF";
        ram_buffer(62709) := X"8FC30058";
        ram_buffer(62710) := X"00000000";
        ram_buffer(62711) := X"00621021";
        ram_buffer(62712) := X"90420000";
        ram_buffer(62713) := X"00000000";
        ram_buffer(62714) := X"A3C20060";
        ram_buffer(62715) := X"AFC00028";
        ram_buffer(62716) := X"8FC2007C";
        ram_buffer(62717) := X"00000000";
        ram_buffer(62718) := X"8C420000";
        ram_buffer(62719) := X"00000000";
        ram_buffer(62720) := X"24420002";
        ram_buffer(62721) := X"AFC20018";
        ram_buffer(62722) := X"10000005";
        ram_buffer(62723) := X"00000000";
        ram_buffer(62724) := X"8FC20028";
        ram_buffer(62725) := X"00000000";
        ram_buffer(62726) := X"24420001";
        ram_buffer(62727) := X"AFC20028";
        ram_buffer(62728) := X"8FC20028";
        ram_buffer(62729) := X"8FC30018";
        ram_buffer(62730) := X"00000000";
        ram_buffer(62731) := X"00621021";
        ram_buffer(62732) := X"90430000";
        ram_buffer(62733) := X"24020030";
        ram_buffer(62734) := X"1062FFF5";
        ram_buffer(62735) := X"00000000";
        ram_buffer(62736) := X"8FC20028";
        ram_buffer(62737) := X"8FC30018";
        ram_buffer(62738) := X"00000000";
        ram_buffer(62739) := X"00621021";
        ram_buffer(62740) := X"AFC20018";
        ram_buffer(62741) := X"8FC20018";
        ram_buffer(62742) := X"00000000";
        ram_buffer(62743) := X"AFC2001C";
        ram_buffer(62744) := X"AFC00014";
        ram_buffer(62745) := X"AFC00040";
        ram_buffer(62746) := X"AFC00050";
        ram_buffer(62747) := X"8FC2001C";
        ram_buffer(62748) := X"00000000";
        ram_buffer(62749) := X"90420000";
        ram_buffer(62750) := X"00000000";
        ram_buffer(62751) := X"00401821";
        ram_buffer(62752) := X"3C02100D";
        ram_buffer(62753) := X"2442B290";
        ram_buffer(62754) := X"00621021";
        ram_buffer(62755) := X"90420000";
        ram_buffer(62756) := X"00000000";
        ram_buffer(62757) := X"14400042";
        ram_buffer(62758) := X"00000000";
        ram_buffer(62759) := X"24020001";
        ram_buffer(62760) := X"AFC20040";
        ram_buffer(62761) := X"8FC6005C";
        ram_buffer(62762) := X"8FC50058";
        ram_buffer(62763) := X"8FC4001C";
        ram_buffer(62764) := X"0C028525";
        ram_buffer(62765) := X"00000000";
        ram_buffer(62766) := X"14400077";
        ram_buffer(62767) := X"00000000";
        ram_buffer(62768) := X"8FC3001C";
        ram_buffer(62769) := X"8FC2005C";
        ram_buffer(62770) := X"00000000";
        ram_buffer(62771) := X"00621021";
        ram_buffer(62772) := X"AFC2001C";
        ram_buffer(62773) := X"8FC2001C";
        ram_buffer(62774) := X"00000000";
        ram_buffer(62775) := X"AFC20014";
        ram_buffer(62776) := X"8FC2001C";
        ram_buffer(62777) := X"00000000";
        ram_buffer(62778) := X"90420000";
        ram_buffer(62779) := X"00000000";
        ram_buffer(62780) := X"00401821";
        ram_buffer(62781) := X"3C02100D";
        ram_buffer(62782) := X"2442B290";
        ram_buffer(62783) := X"00621021";
        ram_buffer(62784) := X"90420000";
        ram_buffer(62785) := X"00000000";
        ram_buffer(62786) := X"10400066";
        ram_buffer(62787) := X"00000000";
        ram_buffer(62788) := X"10000005";
        ram_buffer(62789) := X"00000000";
        ram_buffer(62790) := X"8FC2001C";
        ram_buffer(62791) := X"00000000";
        ram_buffer(62792) := X"24420001";
        ram_buffer(62793) := X"AFC2001C";
        ram_buffer(62794) := X"8FC2001C";
        ram_buffer(62795) := X"00000000";
        ram_buffer(62796) := X"90430000";
        ram_buffer(62797) := X"24020030";
        ram_buffer(62798) := X"1062FFF7";
        ram_buffer(62799) := X"00000000";
        ram_buffer(62800) := X"8FC2001C";
        ram_buffer(62801) := X"00000000";
        ram_buffer(62802) := X"90420000";
        ram_buffer(62803) := X"00000000";
        ram_buffer(62804) := X"00401821";
        ram_buffer(62805) := X"3C02100D";
        ram_buffer(62806) := X"2442B290";
        ram_buffer(62807) := X"00621021";
        ram_buffer(62808) := X"90420000";
        ram_buffer(62809) := X"00000000";
        ram_buffer(62810) := X"10400002";
        ram_buffer(62811) := X"00000000";
        ram_buffer(62812) := X"AFC00040";
        ram_buffer(62813) := X"24020001";
        ram_buffer(62814) := X"AFC20028";
        ram_buffer(62815) := X"8FC2001C";
        ram_buffer(62816) := X"00000000";
        ram_buffer(62817) := X"AFC20018";
        ram_buffer(62818) := X"10000005";
        ram_buffer(62819) := X"00000000";
        ram_buffer(62820) := X"8FC2001C";
        ram_buffer(62821) := X"00000000";
        ram_buffer(62822) := X"24420001";
        ram_buffer(62823) := X"AFC2001C";
        ram_buffer(62824) := X"8FC2001C";
        ram_buffer(62825) := X"00000000";
        ram_buffer(62826) := X"90420000";
        ram_buffer(62827) := X"00000000";
        ram_buffer(62828) := X"00401821";
        ram_buffer(62829) := X"3C02100D";
        ram_buffer(62830) := X"2442B290";
        ram_buffer(62831) := X"00621021";
        ram_buffer(62832) := X"90420000";
        ram_buffer(62833) := X"00000000";
        ram_buffer(62834) := X"1440FFF1";
        ram_buffer(62835) := X"00000000";
        ram_buffer(62836) := X"8FC6005C";
        ram_buffer(62837) := X"8FC50058";
        ram_buffer(62838) := X"8FC4001C";
        ram_buffer(62839) := X"0C028525";
        ram_buffer(62840) := X"00000000";
        ram_buffer(62841) := X"1440001F";
        ram_buffer(62842) := X"00000000";
        ram_buffer(62843) := X"8FC20014";
        ram_buffer(62844) := X"00000000";
        ram_buffer(62845) := X"1440001B";
        ram_buffer(62846) := X"00000000";
        ram_buffer(62847) := X"8FC3001C";
        ram_buffer(62848) := X"8FC2005C";
        ram_buffer(62849) := X"00000000";
        ram_buffer(62850) := X"00621021";
        ram_buffer(62851) := X"AFC2001C";
        ram_buffer(62852) := X"8FC2001C";
        ram_buffer(62853) := X"00000000";
        ram_buffer(62854) := X"AFC20014";
        ram_buffer(62855) := X"10000005";
        ram_buffer(62856) := X"00000000";
        ram_buffer(62857) := X"8FC2001C";
        ram_buffer(62858) := X"00000000";
        ram_buffer(62859) := X"24420001";
        ram_buffer(62860) := X"AFC2001C";
        ram_buffer(62861) := X"8FC2001C";
        ram_buffer(62862) := X"00000000";
        ram_buffer(62863) := X"90420000";
        ram_buffer(62864) := X"00000000";
        ram_buffer(62865) := X"00401821";
        ram_buffer(62866) := X"3C02100D";
        ram_buffer(62867) := X"2442B290";
        ram_buffer(62868) := X"00621021";
        ram_buffer(62869) := X"90420000";
        ram_buffer(62870) := X"00000000";
        ram_buffer(62871) := X"1440FFF1";
        ram_buffer(62872) := X"00000000";
        ram_buffer(62873) := X"8FC20014";
        ram_buffer(62874) := X"00000000";
        ram_buffer(62875) := X"1040000E";
        ram_buffer(62876) := X"00000000";
        ram_buffer(62877) := X"8FC3001C";
        ram_buffer(62878) := X"8FC20014";
        ram_buffer(62879) := X"00000000";
        ram_buffer(62880) := X"00621023";
        ram_buffer(62881) := X"00021080";
        ram_buffer(62882) := X"00021023";
        ram_buffer(62883) := X"AFC20050";
        ram_buffer(62884) := X"10000005";
        ram_buffer(62885) := X"00000000";
        ram_buffer(62886) := X"00000000";
        ram_buffer(62887) := X"10000002";
        ram_buffer(62888) := X"00000000";
        ram_buffer(62889) := X"00000000";
        ram_buffer(62890) := X"8FC2001C";
        ram_buffer(62891) := X"00000000";
        ram_buffer(62892) := X"AFC20020";
        ram_buffer(62893) := X"8FC2001C";
        ram_buffer(62894) := X"00000000";
        ram_buffer(62895) := X"90420000";
        ram_buffer(62896) := X"24030050";
        ram_buffer(62897) := X"10430004";
        ram_buffer(62898) := X"00000000";
        ram_buffer(62899) := X"24030070";
        ram_buffer(62900) := X"14430063";
        ram_buffer(62901) := X"00000000";
        ram_buffer(62902) := X"AFC00024";
        ram_buffer(62903) := X"8FC2001C";
        ram_buffer(62904) := X"00000000";
        ram_buffer(62905) := X"24420001";
        ram_buffer(62906) := X"AFC2001C";
        ram_buffer(62907) := X"8FC2001C";
        ram_buffer(62908) := X"00000000";
        ram_buffer(62909) := X"90420000";
        ram_buffer(62910) := X"2403002B";
        ram_buffer(62911) := X"10430006";
        ram_buffer(62912) := X"00000000";
        ram_buffer(62913) := X"2403002D";
        ram_buffer(62914) := X"14430007";
        ram_buffer(62915) := X"00000000";
        ram_buffer(62916) := X"24020001";
        ram_buffer(62917) := X"AFC20024";
        ram_buffer(62918) := X"8FC2001C";
        ram_buffer(62919) := X"00000000";
        ram_buffer(62920) := X"24420001";
        ram_buffer(62921) := X"AFC2001C";
        ram_buffer(62922) := X"8FC2001C";
        ram_buffer(62923) := X"00000000";
        ram_buffer(62924) := X"90420000";
        ram_buffer(62925) := X"00000000";
        ram_buffer(62926) := X"00401821";
        ram_buffer(62927) := X"3C02100D";
        ram_buffer(62928) := X"2442B290";
        ram_buffer(62929) := X"00621021";
        ram_buffer(62930) := X"90420000";
        ram_buffer(62931) := X"00000000";
        ram_buffer(62932) := X"AFC20034";
        ram_buffer(62933) := X"8FC20034";
        ram_buffer(62934) := X"00000000";
        ram_buffer(62935) := X"10400006";
        ram_buffer(62936) := X"00000000";
        ram_buffer(62937) := X"8FC20034";
        ram_buffer(62938) := X"00000000";
        ram_buffer(62939) := X"2842001A";
        ram_buffer(62940) := X"14400006";
        ram_buffer(62941) := X"00000000";
        ram_buffer(62942) := X"8FC20020";
        ram_buffer(62943) := X"00000000";
        ram_buffer(62944) := X"AFC2001C";
        ram_buffer(62945) := X"10000036";
        ram_buffer(62946) := X"00000000";
        ram_buffer(62947) := X"8FC20034";
        ram_buffer(62948) := X"00000000";
        ram_buffer(62949) := X"2442FFF0";
        ram_buffer(62950) := X"AFC20054";
        ram_buffer(62951) := X"1000000B";
        ram_buffer(62952) := X"00000000";
        ram_buffer(62953) := X"8FC20054";
        ram_buffer(62954) := X"00000000";
        ram_buffer(62955) := X"00021040";
        ram_buffer(62956) := X"00021880";
        ram_buffer(62957) := X"00431821";
        ram_buffer(62958) := X"8FC20034";
        ram_buffer(62959) := X"00000000";
        ram_buffer(62960) := X"00621021";
        ram_buffer(62961) := X"2442FFF0";
        ram_buffer(62962) := X"AFC20054";
        ram_buffer(62963) := X"8FC2001C";
        ram_buffer(62964) := X"00000000";
        ram_buffer(62965) := X"24420001";
        ram_buffer(62966) := X"AFC2001C";
        ram_buffer(62967) := X"8FC2001C";
        ram_buffer(62968) := X"00000000";
        ram_buffer(62969) := X"90420000";
        ram_buffer(62970) := X"00000000";
        ram_buffer(62971) := X"00401821";
        ram_buffer(62972) := X"3C02100D";
        ram_buffer(62973) := X"2442B290";
        ram_buffer(62974) := X"00621021";
        ram_buffer(62975) := X"90420000";
        ram_buffer(62976) := X"00000000";
        ram_buffer(62977) := X"AFC20034";
        ram_buffer(62978) := X"8FC20034";
        ram_buffer(62979) := X"00000000";
        ram_buffer(62980) := X"10400006";
        ram_buffer(62981) := X"00000000";
        ram_buffer(62982) := X"8FC20034";
        ram_buffer(62983) := X"00000000";
        ram_buffer(62984) := X"2842001A";
        ram_buffer(62985) := X"1440FFDF";
        ram_buffer(62986) := X"00000000";
        ram_buffer(62987) := X"8FC20024";
        ram_buffer(62988) := X"00000000";
        ram_buffer(62989) := X"10400005";
        ram_buffer(62990) := X"00000000";
        ram_buffer(62991) := X"8FC20054";
        ram_buffer(62992) := X"00000000";
        ram_buffer(62993) := X"00021023";
        ram_buffer(62994) := X"AFC20054";
        ram_buffer(62995) := X"8FC30050";
        ram_buffer(62996) := X"8FC20054";
        ram_buffer(62997) := X"00000000";
        ram_buffer(62998) := X"00621021";
        ram_buffer(62999) := X"AFC20050";
        ram_buffer(63000) := X"8FC2007C";
        ram_buffer(63001) := X"8FC3001C";
        ram_buffer(63002) := X"00000000";
        ram_buffer(63003) := X"AC430000";
        ram_buffer(63004) := X"8FC20040";
        ram_buffer(63005) := X"00000000";
        ram_buffer(63006) := X"1040000B";
        ram_buffer(63007) := X"00000000";
        ram_buffer(63008) := X"8FC20028";
        ram_buffer(63009) := X"00000000";
        ram_buffer(63010) := X"10400004";
        ram_buffer(63011) := X"00000000";
        ram_buffer(63012) := X"00001021";
        ram_buffer(63013) := X"10000266";
        ram_buffer(63014) := X"00000000";
        ram_buffer(63015) := X"24020006";
        ram_buffer(63016) := X"10000263";
        ram_buffer(63017) := X"00000000";
        ram_buffer(63018) := X"8FC30020";
        ram_buffer(63019) := X"8FC20018";
        ram_buffer(63020) := X"00000000";
        ram_buffer(63021) := X"00621023";
        ram_buffer(63022) := X"2442FFFF";
        ram_buffer(63023) := X"AFC20034";
        ram_buffer(63024) := X"AFC00030";
        ram_buffer(63025) := X"10000009";
        ram_buffer(63026) := X"00000000";
        ram_buffer(63027) := X"8FC20030";
        ram_buffer(63028) := X"00000000";
        ram_buffer(63029) := X"24420001";
        ram_buffer(63030) := X"AFC20030";
        ram_buffer(63031) := X"8FC20034";
        ram_buffer(63032) := X"00000000";
        ram_buffer(63033) := X"00021043";
        ram_buffer(63034) := X"AFC20034";
        ram_buffer(63035) := X"8FC20034";
        ram_buffer(63036) := X"00000000";
        ram_buffer(63037) := X"28420008";
        ram_buffer(63038) := X"1040FFF4";
        ram_buffer(63039) := X"00000000";
        ram_buffer(63040) := X"8FC50030";
        ram_buffer(63041) := X"8FC40078";
        ram_buffer(63042) := X"0C02BDA8";
        ram_buffer(63043) := X"00000000";
        ram_buffer(63044) := X"AFC20010";
        ram_buffer(63045) := X"8FC20010";
        ram_buffer(63046) := X"00000000";
        ram_buffer(63047) := X"24420014";
        ram_buffer(63048) := X"AFC2004C";
        ram_buffer(63049) := X"AFC00034";
        ram_buffer(63050) := X"AFC00044";
        ram_buffer(63051) := X"10000054";
        ram_buffer(63052) := X"00000000";
        ram_buffer(63053) := X"8FC20020";
        ram_buffer(63054) := X"00000000";
        ram_buffer(63055) := X"2442FFFF";
        ram_buffer(63056) := X"AFC20020";
        ram_buffer(63057) := X"8FC20020";
        ram_buffer(63058) := X"00000000";
        ram_buffer(63059) := X"90420000";
        ram_buffer(63060) := X"93C30060";
        ram_buffer(63061) := X"00000000";
        ram_buffer(63062) := X"14620025";
        ram_buffer(63063) := X"00000000";
        ram_buffer(63064) := X"24030001";
        ram_buffer(63065) := X"8FC2005C";
        ram_buffer(63066) := X"00000000";
        ram_buffer(63067) := X"00621023";
        ram_buffer(63068) := X"8FC30020";
        ram_buffer(63069) := X"00000000";
        ram_buffer(63070) := X"00621821";
        ram_buffer(63071) := X"8FC20018";
        ram_buffer(63072) := X"00000000";
        ram_buffer(63073) := X"0062102B";
        ram_buffer(63074) := X"14400019";
        ram_buffer(63075) := X"00000000";
        ram_buffer(63076) := X"24030001";
        ram_buffer(63077) := X"8FC2005C";
        ram_buffer(63078) := X"00000000";
        ram_buffer(63079) := X"00621023";
        ram_buffer(63080) := X"8FC30020";
        ram_buffer(63081) := X"00000000";
        ram_buffer(63082) := X"00621021";
        ram_buffer(63083) := X"8FC6005C";
        ram_buffer(63084) := X"8FC50058";
        ram_buffer(63085) := X"00402021";
        ram_buffer(63086) := X"0C028525";
        ram_buffer(63087) := X"00000000";
        ram_buffer(63088) := X"1440000B";
        ram_buffer(63089) := X"00000000";
        ram_buffer(63090) := X"24030001";
        ram_buffer(63091) := X"8FC2005C";
        ram_buffer(63092) := X"00000000";
        ram_buffer(63093) := X"00621023";
        ram_buffer(63094) := X"8FC30020";
        ram_buffer(63095) := X"00000000";
        ram_buffer(63096) := X"00621021";
        ram_buffer(63097) := X"AFC20020";
        ram_buffer(63098) := X"10000025";
        ram_buffer(63099) := X"00000000";
        ram_buffer(63100) := X"8FC30034";
        ram_buffer(63101) := X"24020020";
        ram_buffer(63102) := X"1462000A";
        ram_buffer(63103) := X"00000000";
        ram_buffer(63104) := X"8FC2004C";
        ram_buffer(63105) := X"00000000";
        ram_buffer(63106) := X"24430004";
        ram_buffer(63107) := X"AFC3004C";
        ram_buffer(63108) := X"8FC30044";
        ram_buffer(63109) := X"00000000";
        ram_buffer(63110) := X"AC430000";
        ram_buffer(63111) := X"AFC00044";
        ram_buffer(63112) := X"AFC00034";
        ram_buffer(63113) := X"8FC20020";
        ram_buffer(63114) := X"00000000";
        ram_buffer(63115) := X"90420000";
        ram_buffer(63116) := X"00000000";
        ram_buffer(63117) := X"00401821";
        ram_buffer(63118) := X"3C02100D";
        ram_buffer(63119) := X"2442B290";
        ram_buffer(63120) := X"00621021";
        ram_buffer(63121) := X"90420000";
        ram_buffer(63122) := X"00000000";
        ram_buffer(63123) := X"3043000F";
        ram_buffer(63124) := X"8FC20034";
        ram_buffer(63125) := X"00000000";
        ram_buffer(63126) := X"00431004";
        ram_buffer(63127) := X"00401821";
        ram_buffer(63128) := X"8FC20044";
        ram_buffer(63129) := X"00000000";
        ram_buffer(63130) := X"00431025";
        ram_buffer(63131) := X"AFC20044";
        ram_buffer(63132) := X"8FC20034";
        ram_buffer(63133) := X"00000000";
        ram_buffer(63134) := X"24420004";
        ram_buffer(63135) := X"AFC20034";
        ram_buffer(63136) := X"8FC30020";
        ram_buffer(63137) := X"8FC20018";
        ram_buffer(63138) := X"00000000";
        ram_buffer(63139) := X"0043102B";
        ram_buffer(63140) := X"1440FFA8";
        ram_buffer(63141) := X"00000000";
        ram_buffer(63142) := X"8FC2004C";
        ram_buffer(63143) := X"00000000";
        ram_buffer(63144) := X"24430004";
        ram_buffer(63145) := X"AFC3004C";
        ram_buffer(63146) := X"8FC30044";
        ram_buffer(63147) := X"00000000";
        ram_buffer(63148) := X"AC430000";
        ram_buffer(63149) := X"8FC2004C";
        ram_buffer(63150) := X"8FC30010";
        ram_buffer(63151) := X"00000000";
        ram_buffer(63152) := X"24630014";
        ram_buffer(63153) := X"00431023";
        ram_buffer(63154) := X"00021083";
        ram_buffer(63155) := X"AFC20034";
        ram_buffer(63156) := X"8FC20010";
        ram_buffer(63157) := X"8FC30034";
        ram_buffer(63158) := X"00000000";
        ram_buffer(63159) := X"AC430010";
        ram_buffer(63160) := X"8FC20034";
        ram_buffer(63161) := X"00000000";
        ram_buffer(63162) := X"00028140";
        ram_buffer(63163) := X"8FC40044";
        ram_buffer(63164) := X"0C02BF41";
        ram_buffer(63165) := X"00000000";
        ram_buffer(63166) := X"02021023";
        ram_buffer(63167) := X"AFC20034";
        ram_buffer(63168) := X"8FC20080";
        ram_buffer(63169) := X"00000000";
        ram_buffer(63170) := X"8C420000";
        ram_buffer(63171) := X"00000000";
        ram_buffer(63172) := X"AFC20038";
        ram_buffer(63173) := X"AFC00048";
        ram_buffer(63174) := X"8FC20010";
        ram_buffer(63175) := X"00000000";
        ram_buffer(63176) := X"24420014";
        ram_buffer(63177) := X"AFC2004C";
        ram_buffer(63178) := X"8FC30034";
        ram_buffer(63179) := X"8FC20038";
        ram_buffer(63180) := X"00000000";
        ram_buffer(63181) := X"0043102A";
        ram_buffer(63182) := X"1040003F";
        ram_buffer(63183) := X"00000000";
        ram_buffer(63184) := X"8FC30034";
        ram_buffer(63185) := X"8FC20038";
        ram_buffer(63186) := X"00000000";
        ram_buffer(63187) := X"00621023";
        ram_buffer(63188) := X"AFC20034";
        ram_buffer(63189) := X"8FC50034";
        ram_buffer(63190) := X"8FC40010";
        ram_buffer(63191) := X"0C02C617";
        ram_buffer(63192) := X"00000000";
        ram_buffer(63193) := X"10400029";
        ram_buffer(63194) := X"00000000";
        ram_buffer(63195) := X"24020001";
        ram_buffer(63196) := X"AFC20048";
        ram_buffer(63197) := X"8FC20034";
        ram_buffer(63198) := X"00000000";
        ram_buffer(63199) := X"2442FFFF";
        ram_buffer(63200) := X"AFC20030";
        ram_buffer(63201) := X"8FC20030";
        ram_buffer(63202) := X"00000000";
        ram_buffer(63203) := X"00021143";
        ram_buffer(63204) := X"00021080";
        ram_buffer(63205) := X"8FC3004C";
        ram_buffer(63206) := X"00000000";
        ram_buffer(63207) := X"00621021";
        ram_buffer(63208) := X"8C420000";
        ram_buffer(63209) := X"8FC30030";
        ram_buffer(63210) := X"00000000";
        ram_buffer(63211) := X"3063001F";
        ram_buffer(63212) := X"24040001";
        ram_buffer(63213) := X"00641804";
        ram_buffer(63214) := X"00431024";
        ram_buffer(63215) := X"10400013";
        ram_buffer(63216) := X"00000000";
        ram_buffer(63217) := X"24020002";
        ram_buffer(63218) := X"AFC20048";
        ram_buffer(63219) := X"8FC20030";
        ram_buffer(63220) := X"00000000";
        ram_buffer(63221) := X"28420002";
        ram_buffer(63222) := X"1440000C";
        ram_buffer(63223) := X"00000000";
        ram_buffer(63224) := X"8FC20030";
        ram_buffer(63225) := X"00000000";
        ram_buffer(63226) := X"2442FFFF";
        ram_buffer(63227) := X"00402821";
        ram_buffer(63228) := X"8FC40010";
        ram_buffer(63229) := X"0C02C617";
        ram_buffer(63230) := X"00000000";
        ram_buffer(63231) := X"10400003";
        ram_buffer(63232) := X"00000000";
        ram_buffer(63233) := X"24020003";
        ram_buffer(63234) := X"AFC20048";
        ram_buffer(63235) := X"8FC50034";
        ram_buffer(63236) := X"8FC40010";
        ram_buffer(63237) := X"0C02F3D8";
        ram_buffer(63238) := X"00000000";
        ram_buffer(63239) := X"8FC30050";
        ram_buffer(63240) := X"8FC20034";
        ram_buffer(63241) := X"00000000";
        ram_buffer(63242) := X"00621021";
        ram_buffer(63243) := X"AFC20050";
        ram_buffer(63244) := X"1000001B";
        ram_buffer(63245) := X"00000000";
        ram_buffer(63246) := X"8FC30034";
        ram_buffer(63247) := X"8FC20038";
        ram_buffer(63248) := X"00000000";
        ram_buffer(63249) := X"0062102A";
        ram_buffer(63250) := X"10400015";
        ram_buffer(63251) := X"00000000";
        ram_buffer(63252) := X"8FC30038";
        ram_buffer(63253) := X"8FC20034";
        ram_buffer(63254) := X"00000000";
        ram_buffer(63255) := X"00621023";
        ram_buffer(63256) := X"AFC20034";
        ram_buffer(63257) := X"8FC60034";
        ram_buffer(63258) := X"8FC50010";
        ram_buffer(63259) := X"8FC40078";
        ram_buffer(63260) := X"0C02C1BB";
        ram_buffer(63261) := X"00000000";
        ram_buffer(63262) := X"AFC20010";
        ram_buffer(63263) := X"8FC30050";
        ram_buffer(63264) := X"8FC20034";
        ram_buffer(63265) := X"00000000";
        ram_buffer(63266) := X"00621023";
        ram_buffer(63267) := X"AFC20050";
        ram_buffer(63268) := X"8FC20010";
        ram_buffer(63269) := X"00000000";
        ram_buffer(63270) := X"24420014";
        ram_buffer(63271) := X"AFC2004C";
        ram_buffer(63272) := X"8FC20080";
        ram_buffer(63273) := X"00000000";
        ram_buffer(63274) := X"8C430008";
        ram_buffer(63275) := X"8FC20050";
        ram_buffer(63276) := X"00000000";
        ram_buffer(63277) := X"0062102A";
        ram_buffer(63278) := X"1040000E";
        ram_buffer(63279) := X"00000000";
        ram_buffer(63280) := X"10000002";
        ram_buffer(63281) := X"00000000";
        ram_buffer(63282) := X"00000000";
        ram_buffer(63283) := X"8FC50010";
        ram_buffer(63284) := X"8FC40078";
        ram_buffer(63285) := X"0C02BE10";
        ram_buffer(63286) := X"00000000";
        ram_buffer(63287) := X"8FC20088";
        ram_buffer(63288) := X"00000000";
        ram_buffer(63289) := X"AC400000";
        ram_buffer(63290) := X"240200A3";
        ram_buffer(63291) := X"10000150";
        ram_buffer(63292) := X"00000000";
        ram_buffer(63293) := X"24020001";
        ram_buffer(63294) := X"AFC2002C";
        ram_buffer(63295) := X"8FC20080";
        ram_buffer(63296) := X"00000000";
        ram_buffer(63297) := X"8C430004";
        ram_buffer(63298) := X"8FC20050";
        ram_buffer(63299) := X"00000000";
        ram_buffer(63300) := X"0043102A";
        ram_buffer(63301) := X"10400093";
        ram_buffer(63302) := X"00000000";
        ram_buffer(63303) := X"24020002";
        ram_buffer(63304) := X"AFC2002C";
        ram_buffer(63305) := X"8FC20080";
        ram_buffer(63306) := X"00000000";
        ram_buffer(63307) := X"8C430004";
        ram_buffer(63308) := X"8FC20050";
        ram_buffer(63309) := X"00000000";
        ram_buffer(63310) := X"00621023";
        ram_buffer(63311) := X"AFC20034";
        ram_buffer(63312) := X"8FC30034";
        ram_buffer(63313) := X"8FC20038";
        ram_buffer(63314) := X"00000000";
        ram_buffer(63315) := X"0062102A";
        ram_buffer(63316) := X"1440004D";
        ram_buffer(63317) := X"00000000";
        ram_buffer(63318) := X"8FC20080";
        ram_buffer(63319) := X"00000000";
        ram_buffer(63320) := X"8C42000C";
        ram_buffer(63321) := X"24030002";
        ram_buffer(63322) := X"1043001C";
        ram_buffer(63323) := X"00000000";
        ram_buffer(63324) := X"24030003";
        ram_buffer(63325) := X"1043001F";
        ram_buffer(63326) := X"00000000";
        ram_buffer(63327) := X"24030001";
        ram_buffer(63328) := X"14430037";
        ram_buffer(63329) := X"00000000";
        ram_buffer(63330) := X"8FC30034";
        ram_buffer(63331) := X"8FC20038";
        ram_buffer(63332) := X"00000000";
        ram_buffer(63333) := X"1462002E";
        ram_buffer(63334) := X"00000000";
        ram_buffer(63335) := X"8FC20034";
        ram_buffer(63336) := X"00000000";
        ram_buffer(63337) := X"28420002";
        ram_buffer(63338) := X"14400016";
        ram_buffer(63339) := X"00000000";
        ram_buffer(63340) := X"8FC20034";
        ram_buffer(63341) := X"00000000";
        ram_buffer(63342) := X"2442FFFF";
        ram_buffer(63343) := X"00402821";
        ram_buffer(63344) := X"8FC40010";
        ram_buffer(63345) := X"0C02C617";
        ram_buffer(63346) := X"00000000";
        ram_buffer(63347) := X"1440000D";
        ram_buffer(63348) := X"00000000";
        ram_buffer(63349) := X"1000001E";
        ram_buffer(63350) := X"00000000";
        ram_buffer(63351) := X"8FC2008C";
        ram_buffer(63352) := X"00000000";
        ram_buffer(63353) := X"1440001D";
        ram_buffer(63354) := X"00000000";
        ram_buffer(63355) := X"10000005";
        ram_buffer(63356) := X"00000000";
        ram_buffer(63357) := X"8FC2008C";
        ram_buffer(63358) := X"00000000";
        ram_buffer(63359) := X"10400018";
        ram_buffer(63360) := X"00000000";
        ram_buffer(63361) := X"8FC20080";
        ram_buffer(63362) := X"00000000";
        ram_buffer(63363) := X"8C430004";
        ram_buffer(63364) := X"8FC20084";
        ram_buffer(63365) := X"00000000";
        ram_buffer(63366) := X"AC430000";
        ram_buffer(63367) := X"8FC20010";
        ram_buffer(63368) := X"24030001";
        ram_buffer(63369) := X"AC430010";
        ram_buffer(63370) := X"8FC2004C";
        ram_buffer(63371) := X"24030001";
        ram_buffer(63372) := X"AC430000";
        ram_buffer(63373) := X"8FC20088";
        ram_buffer(63374) := X"8FC30010";
        ram_buffer(63375) := X"00000000";
        ram_buffer(63376) := X"AC430000";
        ram_buffer(63377) := X"24020062";
        ram_buffer(63378) := X"100000F9";
        ram_buffer(63379) := X"00000000";
        ram_buffer(63380) := X"00000000";
        ram_buffer(63381) := X"10000002";
        ram_buffer(63382) := X"00000000";
        ram_buffer(63383) := X"00000000";
        ram_buffer(63384) := X"8FC50010";
        ram_buffer(63385) := X"8FC40078";
        ram_buffer(63386) := X"0C02BE10";
        ram_buffer(63387) := X"00000000";
        ram_buffer(63388) := X"8FC20088";
        ram_buffer(63389) := X"00000000";
        ram_buffer(63390) := X"AC400000";
        ram_buffer(63391) := X"24020050";
        ram_buffer(63392) := X"100000EB";
        ram_buffer(63393) := X"00000000";
        ram_buffer(63394) := X"8FC20034";
        ram_buffer(63395) := X"00000000";
        ram_buffer(63396) := X"2442FFFF";
        ram_buffer(63397) := X"AFC20030";
        ram_buffer(63398) := X"8FC20048";
        ram_buffer(63399) := X"00000000";
        ram_buffer(63400) := X"10400005";
        ram_buffer(63401) := X"00000000";
        ram_buffer(63402) := X"24020001";
        ram_buffer(63403) := X"AFC20048";
        ram_buffer(63404) := X"1000000A";
        ram_buffer(63405) := X"00000000";
        ram_buffer(63406) := X"8FC20030";
        ram_buffer(63407) := X"00000000";
        ram_buffer(63408) := X"18400006";
        ram_buffer(63409) := X"00000000";
        ram_buffer(63410) := X"8FC50030";
        ram_buffer(63411) := X"8FC40010";
        ram_buffer(63412) := X"0C02C617";
        ram_buffer(63413) := X"00000000";
        ram_buffer(63414) := X"AFC20048";
        ram_buffer(63415) := X"8FC20030";
        ram_buffer(63416) := X"00000000";
        ram_buffer(63417) := X"00021143";
        ram_buffer(63418) := X"00021080";
        ram_buffer(63419) := X"8FC3004C";
        ram_buffer(63420) := X"00000000";
        ram_buffer(63421) := X"00621021";
        ram_buffer(63422) := X"8C420000";
        ram_buffer(63423) := X"8FC30030";
        ram_buffer(63424) := X"00000000";
        ram_buffer(63425) := X"3063001F";
        ram_buffer(63426) := X"24040001";
        ram_buffer(63427) := X"00641804";
        ram_buffer(63428) := X"00431024";
        ram_buffer(63429) := X"10400005";
        ram_buffer(63430) := X"00000000";
        ram_buffer(63431) := X"8FC20048";
        ram_buffer(63432) := X"00000000";
        ram_buffer(63433) := X"34420002";
        ram_buffer(63434) := X"AFC20048";
        ram_buffer(63435) := X"8FC30038";
        ram_buffer(63436) := X"8FC20034";
        ram_buffer(63437) := X"00000000";
        ram_buffer(63438) := X"00621023";
        ram_buffer(63439) := X"AFC20038";
        ram_buffer(63440) := X"8FC50034";
        ram_buffer(63441) := X"8FC40010";
        ram_buffer(63442) := X"0C02F3D8";
        ram_buffer(63443) := X"00000000";
        ram_buffer(63444) := X"8FC20080";
        ram_buffer(63445) := X"00000000";
        ram_buffer(63446) := X"8C420004";
        ram_buffer(63447) := X"00000000";
        ram_buffer(63448) := X"AFC20050";
        ram_buffer(63449) := X"8FC20048";
        ram_buffer(63450) := X"00000000";
        ram_buffer(63451) := X"104000A7";
        ram_buffer(63452) := X"00000000";
        ram_buffer(63453) := X"AFC0003C";
        ram_buffer(63454) := X"8FC20080";
        ram_buffer(63455) := X"00000000";
        ram_buffer(63456) := X"8C42000C";
        ram_buffer(63457) := X"24030001";
        ram_buffer(63458) := X"1043000C";
        ram_buffer(63459) := X"00000000";
        ram_buffer(63460) := X"28430002";
        ram_buffer(63461) := X"14600027";
        ram_buffer(63462) := X"00000000";
        ram_buffer(63463) := X"24030002";
        ram_buffer(63464) := X"10430018";
        ram_buffer(63465) := X"00000000";
        ram_buffer(63466) := X"24030003";
        ram_buffer(63467) := X"1043001C";
        ram_buffer(63468) := X"00000000";
        ram_buffer(63469) := X"10000023";
        ram_buffer(63470) := X"00000000";
        ram_buffer(63471) := X"8FC20048";
        ram_buffer(63472) := X"00000000";
        ram_buffer(63473) := X"30420002";
        ram_buffer(63474) := X"1040001D";
        ram_buffer(63475) := X"00000000";
        ram_buffer(63476) := X"8FC2004C";
        ram_buffer(63477) := X"00000000";
        ram_buffer(63478) := X"8C430000";
        ram_buffer(63479) := X"8FC20048";
        ram_buffer(63480) := X"00000000";
        ram_buffer(63481) := X"00621025";
        ram_buffer(63482) := X"30420001";
        ram_buffer(63483) := X"10400014";
        ram_buffer(63484) := X"00000000";
        ram_buffer(63485) := X"24020001";
        ram_buffer(63486) := X"AFC2003C";
        ram_buffer(63487) := X"10000010";
        ram_buffer(63488) := X"00000000";
        ram_buffer(63489) := X"24030001";
        ram_buffer(63490) := X"8FC2008C";
        ram_buffer(63491) := X"00000000";
        ram_buffer(63492) := X"00621023";
        ram_buffer(63493) := X"AFC2003C";
        ram_buffer(63494) := X"1000000A";
        ram_buffer(63495) := X"00000000";
        ram_buffer(63496) := X"8FC2008C";
        ram_buffer(63497) := X"00000000";
        ram_buffer(63498) := X"AFC2003C";
        ram_buffer(63499) := X"10000005";
        ram_buffer(63500) := X"00000000";
        ram_buffer(63501) := X"00000000";
        ram_buffer(63502) := X"10000002";
        ram_buffer(63503) := X"00000000";
        ram_buffer(63504) := X"00000000";
        ram_buffer(63505) := X"8FC2003C";
        ram_buffer(63506) := X"00000000";
        ram_buffer(63507) := X"1040006B";
        ram_buffer(63508) := X"00000000";
        ram_buffer(63509) := X"8FC20010";
        ram_buffer(63510) := X"00000000";
        ram_buffer(63511) := X"8C420010";
        ram_buffer(63512) := X"00000000";
        ram_buffer(63513) := X"AFC20030";
        ram_buffer(63514) := X"8FC50010";
        ram_buffer(63515) := X"8FC40078";
        ram_buffer(63516) := X"0C02F46F";
        ram_buffer(63517) := X"00000000";
        ram_buffer(63518) := X"AFC20010";
        ram_buffer(63519) := X"8FC20010";
        ram_buffer(63520) := X"00000000";
        ram_buffer(63521) := X"24420014";
        ram_buffer(63522) := X"AFC2004C";
        ram_buffer(63523) := X"8FC3002C";
        ram_buffer(63524) := X"24020002";
        ram_buffer(63525) := X"1462001E";
        ram_buffer(63526) := X"00000000";
        ram_buffer(63527) := X"8FC20080";
        ram_buffer(63528) := X"00000000";
        ram_buffer(63529) := X"8C420000";
        ram_buffer(63530) := X"00000000";
        ram_buffer(63531) := X"2443FFFF";
        ram_buffer(63532) := X"8FC20038";
        ram_buffer(63533) := X"00000000";
        ram_buffer(63534) := X"1462004A";
        ram_buffer(63535) := X"00000000";
        ram_buffer(63536) := X"8FC20038";
        ram_buffer(63537) := X"00000000";
        ram_buffer(63538) := X"00021143";
        ram_buffer(63539) := X"00021080";
        ram_buffer(63540) := X"8FC3004C";
        ram_buffer(63541) := X"00000000";
        ram_buffer(63542) := X"00621021";
        ram_buffer(63543) := X"8C420000";
        ram_buffer(63544) := X"8FC30038";
        ram_buffer(63545) := X"00000000";
        ram_buffer(63546) := X"3063001F";
        ram_buffer(63547) := X"24040001";
        ram_buffer(63548) := X"00641804";
        ram_buffer(63549) := X"00431024";
        ram_buffer(63550) := X"1040003A";
        ram_buffer(63551) := X"00000000";
        ram_buffer(63552) := X"24020001";
        ram_buffer(63553) := X"AFC2002C";
        ram_buffer(63554) := X"10000036";
        ram_buffer(63555) := X"00000000";
        ram_buffer(63556) := X"8FC20010";
        ram_buffer(63557) := X"00000000";
        ram_buffer(63558) := X"8C430010";
        ram_buffer(63559) := X"8FC20030";
        ram_buffer(63560) := X"00000000";
        ram_buffer(63561) := X"0043102A";
        ram_buffer(63562) := X"1440001E";
        ram_buffer(63563) := X"00000000";
        ram_buffer(63564) := X"8FC20038";
        ram_buffer(63565) := X"00000000";
        ram_buffer(63566) := X"3042001F";
        ram_buffer(63567) := X"AFC20034";
        ram_buffer(63568) := X"8FC20034";
        ram_buffer(63569) := X"00000000";
        ram_buffer(63570) := X"10400026";
        ram_buffer(63571) := X"00000000";
        ram_buffer(63572) := X"8FC30030";
        ram_buffer(63573) := X"3C023FFF";
        ram_buffer(63574) := X"3442FFFF";
        ram_buffer(63575) := X"00621021";
        ram_buffer(63576) := X"00021080";
        ram_buffer(63577) := X"8FC3004C";
        ram_buffer(63578) := X"00000000";
        ram_buffer(63579) := X"00621021";
        ram_buffer(63580) := X"8C420000";
        ram_buffer(63581) := X"00000000";
        ram_buffer(63582) := X"00402021";
        ram_buffer(63583) := X"0C02BF41";
        ram_buffer(63584) := X"00000000";
        ram_buffer(63585) := X"00402021";
        ram_buffer(63586) := X"24030020";
        ram_buffer(63587) := X"8FC20034";
        ram_buffer(63588) := X"00000000";
        ram_buffer(63589) := X"00621023";
        ram_buffer(63590) := X"0082102A";
        ram_buffer(63591) := X"10400011";
        ram_buffer(63592) := X"00000000";
        ram_buffer(63593) := X"24050001";
        ram_buffer(63594) := X"8FC40010";
        ram_buffer(63595) := X"0C02F3D8";
        ram_buffer(63596) := X"00000000";
        ram_buffer(63597) := X"8FC20050";
        ram_buffer(63598) := X"00000000";
        ram_buffer(63599) := X"24420001";
        ram_buffer(63600) := X"AFC20050";
        ram_buffer(63601) := X"8FC20080";
        ram_buffer(63602) := X"00000000";
        ram_buffer(63603) := X"8C420008";
        ram_buffer(63604) := X"8FC30050";
        ram_buffer(63605) := X"00000000";
        ram_buffer(63606) := X"0043102A";
        ram_buffer(63607) := X"1440FEBA";
        ram_buffer(63608) := X"00000000";
        ram_buffer(63609) := X"8FC2002C";
        ram_buffer(63610) := X"00000000";
        ram_buffer(63611) := X"34420020";
        ram_buffer(63612) := X"AFC2002C";
        ram_buffer(63613) := X"10000005";
        ram_buffer(63614) := X"00000000";
        ram_buffer(63615) := X"8FC2002C";
        ram_buffer(63616) := X"00000000";
        ram_buffer(63617) := X"34420010";
        ram_buffer(63618) := X"AFC2002C";
        ram_buffer(63619) := X"8FC20088";
        ram_buffer(63620) := X"8FC30010";
        ram_buffer(63621) := X"00000000";
        ram_buffer(63622) := X"AC430000";
        ram_buffer(63623) := X"8FC20084";
        ram_buffer(63624) := X"8FC30050";
        ram_buffer(63625) := X"00000000";
        ram_buffer(63626) := X"AC430000";
        ram_buffer(63627) := X"8FC2002C";
        ram_buffer(63628) := X"03C0E821";
        ram_buffer(63629) := X"8FBF0074";
        ram_buffer(63630) := X"8FBE0070";
        ram_buffer(63631) := X"8FB0006C";
        ram_buffer(63632) := X"27BD0078";
        ram_buffer(63633) := X"03E00008";
        ram_buffer(63634) := X"00000000";
        ram_buffer(63635) := X"27BDFFF0";
        ram_buffer(63636) := X"AFBE000C";
        ram_buffer(63637) := X"03A0F021";
        ram_buffer(63638) := X"AFC40010";
        ram_buffer(63639) := X"AFC50014";
        ram_buffer(63640) := X"AFC60018";
        ram_buffer(63641) := X"24030008";
        ram_buffer(63642) := X"8FC20018";
        ram_buffer(63643) := X"00000000";
        ram_buffer(63644) := X"00621023";
        ram_buffer(63645) := X"AFC20018";
        ram_buffer(63646) := X"8FC20018";
        ram_buffer(63647) := X"00000000";
        ram_buffer(63648) := X"00021080";
        ram_buffer(63649) := X"AFC20018";
        ram_buffer(63650) := X"24030020";
        ram_buffer(63651) := X"8FC20018";
        ram_buffer(63652) := X"00000000";
        ram_buffer(63653) := X"00621023";
        ram_buffer(63654) := X"AFC20000";
        ram_buffer(63655) := X"8FC20010";
        ram_buffer(63656) := X"00000000";
        ram_buffer(63657) := X"8C430000";
        ram_buffer(63658) := X"8FC20010";
        ram_buffer(63659) := X"00000000";
        ram_buffer(63660) := X"24420004";
        ram_buffer(63661) := X"8C440000";
        ram_buffer(63662) := X"8FC20000";
        ram_buffer(63663) := X"00000000";
        ram_buffer(63664) := X"00441004";
        ram_buffer(63665) := X"00621825";
        ram_buffer(63666) := X"8FC20010";
        ram_buffer(63667) := X"00000000";
        ram_buffer(63668) := X"AC430000";
        ram_buffer(63669) := X"8FC20010";
        ram_buffer(63670) := X"00000000";
        ram_buffer(63671) := X"24420004";
        ram_buffer(63672) := X"8FC30010";
        ram_buffer(63673) := X"00000000";
        ram_buffer(63674) := X"24630004";
        ram_buffer(63675) := X"8C640000";
        ram_buffer(63676) := X"8FC30018";
        ram_buffer(63677) := X"00000000";
        ram_buffer(63678) := X"00641806";
        ram_buffer(63679) := X"AC430000";
        ram_buffer(63680) := X"8FC20010";
        ram_buffer(63681) := X"00000000";
        ram_buffer(63682) := X"24420004";
        ram_buffer(63683) := X"AFC20010";
        ram_buffer(63684) := X"8FC30010";
        ram_buffer(63685) := X"8FC20014";
        ram_buffer(63686) := X"00000000";
        ram_buffer(63687) := X"0062102B";
        ram_buffer(63688) := X"1440FFDE";
        ram_buffer(63689) := X"00000000";
        ram_buffer(63690) := X"00000000";
        ram_buffer(63691) := X"03C0E821";
        ram_buffer(63692) := X"8FBE000C";
        ram_buffer(63693) := X"27BD0010";
        ram_buffer(63694) := X"03E00008";
        ram_buffer(63695) := X"00000000";
        ram_buffer(63696) := X"27BDFFC0";
        ram_buffer(63697) := X"AFBF003C";
        ram_buffer(63698) := X"AFBE0038";
        ram_buffer(63699) := X"03A0F021";
        ram_buffer(63700) := X"AFC40040";
        ram_buffer(63701) := X"AFC50044";
        ram_buffer(63702) := X"AFC60048";
        ram_buffer(63703) := X"8FC20044";
        ram_buffer(63704) := X"00000000";
        ram_buffer(63705) := X"8C420000";
        ram_buffer(63706) := X"00000000";
        ram_buffer(63707) := X"AFC20028";
        ram_buffer(63708) := X"8FC20028";
        ram_buffer(63709) := X"00000000";
        ram_buffer(63710) := X"00021143";
        ram_buffer(63711) := X"00021080";
        ram_buffer(63712) := X"8FC30048";
        ram_buffer(63713) := X"00000000";
        ram_buffer(63714) := X"00621021";
        ram_buffer(63715) := X"AFC20010";
        ram_buffer(63716) := X"8FC20028";
        ram_buffer(63717) := X"00000000";
        ram_buffer(63718) := X"3042001F";
        ram_buffer(63719) := X"10400005";
        ram_buffer(63720) := X"00000000";
        ram_buffer(63721) := X"8FC20010";
        ram_buffer(63722) := X"00000000";
        ram_buffer(63723) := X"24420004";
        ram_buffer(63724) := X"AFC20010";
        ram_buffer(63725) := X"8FC20010";
        ram_buffer(63726) := X"00000000";
        ram_buffer(63727) := X"2442FFFC";
        ram_buffer(63728) := X"AFC20010";
        ram_buffer(63729) := X"8FC20010";
        ram_buffer(63730) := X"00000000";
        ram_buffer(63731) := X"AC400000";
        ram_buffer(63732) := X"8FC20010";
        ram_buffer(63733) := X"00000000";
        ram_buffer(63734) := X"AFC2002C";
        ram_buffer(63735) := X"8FC2002C";
        ram_buffer(63736) := X"00000000";
        ram_buffer(63737) := X"AFC20014";
        ram_buffer(63738) := X"AFC00024";
        ram_buffer(63739) := X"8FC20024";
        ram_buffer(63740) := X"00000000";
        ram_buffer(63741) := X"AFC20020";
        ram_buffer(63742) := X"8FC20020";
        ram_buffer(63743) := X"00000000";
        ram_buffer(63744) := X"AFC2001C";
        ram_buffer(63745) := X"8FC20040";
        ram_buffer(63746) := X"00000000";
        ram_buffer(63747) := X"8C420000";
        ram_buffer(63748) := X"00000000";
        ram_buffer(63749) := X"AFC20018";
        ram_buffer(63750) := X"1000007B";
        ram_buffer(63751) := X"00000000";
        ram_buffer(63752) := X"3C02100D";
        ram_buffer(63753) := X"2443B290";
        ram_buffer(63754) := X"8FC20030";
        ram_buffer(63755) := X"00000000";
        ram_buffer(63756) := X"00621021";
        ram_buffer(63757) := X"90420000";
        ram_buffer(63758) := X"00000000";
        ram_buffer(63759) := X"AFC20034";
        ram_buffer(63760) := X"8FC20034";
        ram_buffer(63761) := X"00000000";
        ram_buffer(63762) := X"14400045";
        ram_buffer(63763) := X"00000000";
        ram_buffer(63764) := X"8FC20030";
        ram_buffer(63765) := X"00000000";
        ram_buffer(63766) := X"2C420021";
        ram_buffer(63767) := X"10400031";
        ram_buffer(63768) := X"00000000";
        ram_buffer(63769) := X"8FC30020";
        ram_buffer(63770) := X"8FC2001C";
        ram_buffer(63771) := X"00000000";
        ram_buffer(63772) := X"0062102A";
        ram_buffer(63773) := X"10400064";
        ram_buffer(63774) := X"00000000";
        ram_buffer(63775) := X"8FC30010";
        ram_buffer(63776) := X"8FC20014";
        ram_buffer(63777) := X"00000000";
        ram_buffer(63778) := X"0062102B";
        ram_buffer(63779) := X"1040000B";
        ram_buffer(63780) := X"00000000";
        ram_buffer(63781) := X"8FC20024";
        ram_buffer(63782) := X"00000000";
        ram_buffer(63783) := X"28420008";
        ram_buffer(63784) := X"10400006";
        ram_buffer(63785) := X"00000000";
        ram_buffer(63786) := X"8FC60024";
        ram_buffer(63787) := X"8FC50014";
        ram_buffer(63788) := X"8FC40010";
        ram_buffer(63789) := X"0C02F893";
        ram_buffer(63790) := X"00000000";
        ram_buffer(63791) := X"8FC30010";
        ram_buffer(63792) := X"8FC20048";
        ram_buffer(63793) := X"00000000";
        ram_buffer(63794) := X"0043102B";
        ram_buffer(63795) := X"14400005";
        ram_buffer(63796) := X"00000000";
        ram_buffer(63797) := X"24020008";
        ram_buffer(63798) := X"AFC20024";
        ram_buffer(63799) := X"1000004A";
        ram_buffer(63800) := X"00000000";
        ram_buffer(63801) := X"8FC2001C";
        ram_buffer(63802) := X"00000000";
        ram_buffer(63803) := X"AFC20020";
        ram_buffer(63804) := X"8FC20010";
        ram_buffer(63805) := X"00000000";
        ram_buffer(63806) := X"2442FFFC";
        ram_buffer(63807) := X"AFC20010";
        ram_buffer(63808) := X"8FC20010";
        ram_buffer(63809) := X"00000000";
        ram_buffer(63810) := X"AC400000";
        ram_buffer(63811) := X"8FC20010";
        ram_buffer(63812) := X"00000000";
        ram_buffer(63813) := X"AFC20014";
        ram_buffer(63814) := X"AFC00024";
        ram_buffer(63815) := X"1000003A";
        ram_buffer(63816) := X"00000000";
        ram_buffer(63817) := X"8FC30030";
        ram_buffer(63818) := X"24020029";
        ram_buffer(63819) := X"14620009";
        ram_buffer(63820) := X"00000000";
        ram_buffer(63821) := X"8FC20018";
        ram_buffer(63822) := X"00000000";
        ram_buffer(63823) := X"24430001";
        ram_buffer(63824) := X"8FC20040";
        ram_buffer(63825) := X"00000000";
        ram_buffer(63826) := X"AC430000";
        ram_buffer(63827) := X"1000003B";
        ram_buffer(63828) := X"00000000";
        ram_buffer(63829) := X"24020004";
        ram_buffer(63830) := X"100000A6";
        ram_buffer(63831) := X"00000000";
        ram_buffer(63832) := X"8FC2001C";
        ram_buffer(63833) := X"00000000";
        ram_buffer(63834) := X"24420001";
        ram_buffer(63835) := X"AFC2001C";
        ram_buffer(63836) := X"8FC20024";
        ram_buffer(63837) := X"00000000";
        ram_buffer(63838) := X"24420001";
        ram_buffer(63839) := X"AFC20024";
        ram_buffer(63840) := X"8FC20024";
        ram_buffer(63841) := X"00000000";
        ram_buffer(63842) := X"28420009";
        ram_buffer(63843) := X"14400012";
        ram_buffer(63844) := X"00000000";
        ram_buffer(63845) := X"8FC30010";
        ram_buffer(63846) := X"8FC20048";
        ram_buffer(63847) := X"00000000";
        ram_buffer(63848) := X"0043102B";
        ram_buffer(63849) := X"14400003";
        ram_buffer(63850) := X"00000000";
        ram_buffer(63851) := X"10000016";
        ram_buffer(63852) := X"00000000";
        ram_buffer(63853) := X"24020001";
        ram_buffer(63854) := X"AFC20024";
        ram_buffer(63855) := X"8FC20010";
        ram_buffer(63856) := X"00000000";
        ram_buffer(63857) := X"2442FFFC";
        ram_buffer(63858) := X"AFC20010";
        ram_buffer(63859) := X"8FC20010";
        ram_buffer(63860) := X"00000000";
        ram_buffer(63861) := X"AC400000";
        ram_buffer(63862) := X"8FC20010";
        ram_buffer(63863) := X"00000000";
        ram_buffer(63864) := X"8C420000";
        ram_buffer(63865) := X"00000000";
        ram_buffer(63866) := X"00021900";
        ram_buffer(63867) := X"8FC20034";
        ram_buffer(63868) := X"00000000";
        ram_buffer(63869) := X"3042000F";
        ram_buffer(63870) := X"00621825";
        ram_buffer(63871) := X"8FC20010";
        ram_buffer(63872) := X"00000000";
        ram_buffer(63873) := X"AC430000";
        ram_buffer(63874) := X"8FC20018";
        ram_buffer(63875) := X"00000000";
        ram_buffer(63876) := X"24420001";
        ram_buffer(63877) := X"AFC20018";
        ram_buffer(63878) := X"8FC20018";
        ram_buffer(63879) := X"00000000";
        ram_buffer(63880) := X"90420000";
        ram_buffer(63881) := X"00000000";
        ram_buffer(63882) := X"AFC20030";
        ram_buffer(63883) := X"8FC20030";
        ram_buffer(63884) := X"00000000";
        ram_buffer(63885) := X"1440FF7A";
        ram_buffer(63886) := X"00000000";
        ram_buffer(63887) := X"8FC2001C";
        ram_buffer(63888) := X"00000000";
        ram_buffer(63889) := X"14400004";
        ram_buffer(63890) := X"00000000";
        ram_buffer(63891) := X"24020004";
        ram_buffer(63892) := X"10000068";
        ram_buffer(63893) := X"00000000";
        ram_buffer(63894) := X"8FC30010";
        ram_buffer(63895) := X"8FC20014";
        ram_buffer(63896) := X"00000000";
        ram_buffer(63897) := X"0062102B";
        ram_buffer(63898) := X"1040000B";
        ram_buffer(63899) := X"00000000";
        ram_buffer(63900) := X"8FC20024";
        ram_buffer(63901) := X"00000000";
        ram_buffer(63902) := X"28420008";
        ram_buffer(63903) := X"10400006";
        ram_buffer(63904) := X"00000000";
        ram_buffer(63905) := X"8FC60024";
        ram_buffer(63906) := X"8FC50014";
        ram_buffer(63907) := X"8FC40010";
        ram_buffer(63908) := X"0C02F893";
        ram_buffer(63909) := X"00000000";
        ram_buffer(63910) := X"8FC30010";
        ram_buffer(63911) := X"8FC20048";
        ram_buffer(63912) := X"00000000";
        ram_buffer(63913) := X"0043102B";
        ram_buffer(63914) := X"10400022";
        ram_buffer(63915) := X"00000000";
        ram_buffer(63916) := X"8FC20048";
        ram_buffer(63917) := X"00000000";
        ram_buffer(63918) := X"AFC20014";
        ram_buffer(63919) := X"8FC20014";
        ram_buffer(63920) := X"00000000";
        ram_buffer(63921) := X"24430004";
        ram_buffer(63922) := X"AFC30014";
        ram_buffer(63923) := X"8FC30010";
        ram_buffer(63924) := X"00000000";
        ram_buffer(63925) := X"24640004";
        ram_buffer(63926) := X"AFC40010";
        ram_buffer(63927) := X"8C630000";
        ram_buffer(63928) := X"00000000";
        ram_buffer(63929) := X"AC430000";
        ram_buffer(63930) := X"8FC30010";
        ram_buffer(63931) := X"8FC2002C";
        ram_buffer(63932) := X"00000000";
        ram_buffer(63933) := X"0043102B";
        ram_buffer(63934) := X"1040FFF0";
        ram_buffer(63935) := X"00000000";
        ram_buffer(63936) := X"8FC20014";
        ram_buffer(63937) := X"00000000";
        ram_buffer(63938) := X"24430004";
        ram_buffer(63939) := X"AFC30014";
        ram_buffer(63940) := X"AC400000";
        ram_buffer(63941) := X"8FC30014";
        ram_buffer(63942) := X"8FC2002C";
        ram_buffer(63943) := X"00000000";
        ram_buffer(63944) := X"0043102B";
        ram_buffer(63945) := X"1040FFF6";
        ram_buffer(63946) := X"00000000";
        ram_buffer(63947) := X"10000016";
        ram_buffer(63948) := X"00000000";
        ram_buffer(63949) := X"8FC20028";
        ram_buffer(63950) := X"00000000";
        ram_buffer(63951) := X"3042001F";
        ram_buffer(63952) := X"AFC20024";
        ram_buffer(63953) := X"8FC20024";
        ram_buffer(63954) := X"00000000";
        ram_buffer(63955) := X"1040000E";
        ram_buffer(63956) := X"00000000";
        ram_buffer(63957) := X"8FC2002C";
        ram_buffer(63958) := X"00000000";
        ram_buffer(63959) := X"8C430000";
        ram_buffer(63960) := X"24040020";
        ram_buffer(63961) := X"8FC20024";
        ram_buffer(63962) := X"00000000";
        ram_buffer(63963) := X"00821023";
        ram_buffer(63964) := X"2404FFFF";
        ram_buffer(63965) := X"00441006";
        ram_buffer(63966) := X"00621824";
        ram_buffer(63967) := X"8FC2002C";
        ram_buffer(63968) := X"00000000";
        ram_buffer(63969) := X"AC430000";
        ram_buffer(63970) := X"8FC2002C";
        ram_buffer(63971) := X"00000000";
        ram_buffer(63972) := X"AFC20014";
        ram_buffer(63973) := X"8FC20014";
        ram_buffer(63974) := X"00000000";
        ram_buffer(63975) := X"8C420000";
        ram_buffer(63976) := X"00000000";
        ram_buffer(63977) := X"14400011";
        ram_buffer(63978) := X"00000000";
        ram_buffer(63979) := X"8FC30014";
        ram_buffer(63980) := X"8FC20048";
        ram_buffer(63981) := X"00000000";
        ram_buffer(63982) := X"14620006";
        ram_buffer(63983) := X"00000000";
        ram_buffer(63984) := X"8FC20014";
        ram_buffer(63985) := X"24030001";
        ram_buffer(63986) := X"AC430000";
        ram_buffer(63987) := X"10000008";
        ram_buffer(63988) := X"00000000";
        ram_buffer(63989) := X"8FC20014";
        ram_buffer(63990) := X"00000000";
        ram_buffer(63991) := X"2442FFFC";
        ram_buffer(63992) := X"AFC20014";
        ram_buffer(63993) := X"1000FFEB";
        ram_buffer(63994) := X"00000000";
        ram_buffer(63995) := X"00000000";
        ram_buffer(63996) := X"24020005";
        ram_buffer(63997) := X"03C0E821";
        ram_buffer(63998) := X"8FBF003C";
        ram_buffer(63999) := X"8FBE0038";
        ram_buffer(64000) := X"27BD0040";
        ram_buffer(64001) := X"03E00008";
        ram_buffer(64002) := X"00000000";
        ram_buffer(64003) := X"27BDFFD0";
        ram_buffer(64004) := X"AFBF002C";
        ram_buffer(64005) := X"AFBE0028";
        ram_buffer(64006) := X"AFB20024";
        ram_buffer(64007) := X"AFB10020";
        ram_buffer(64008) := X"AFB0001C";
        ram_buffer(64009) := X"03A0F021";
        ram_buffer(64010) := X"AFC40030";
        ram_buffer(64011) := X"00A09021";
        ram_buffer(64012) := X"00C08021";
        ram_buffer(64013) := X"8FC20030";
        ram_buffer(64014) := X"00000000";
        ram_buffer(64015) := X"AFC20010";
        ram_buffer(64016) := X"8FC20010";
        ram_buffer(64017) := X"00000000";
        ram_buffer(64018) := X"1040000A";
        ram_buffer(64019) := X"00000000";
        ram_buffer(64020) := X"8FC20010";
        ram_buffer(64021) := X"00000000";
        ram_buffer(64022) := X"8C420038";
        ram_buffer(64023) := X"00000000";
        ram_buffer(64024) := X"14400004";
        ram_buffer(64025) := X"00000000";
        ram_buffer(64026) := X"8FC40010";
        ram_buffer(64027) := X"0C027069";
        ram_buffer(64028) := X"00000000";
        ram_buffer(64029) := X"8E020018";
        ram_buffer(64030) := X"00000000";
        ram_buffer(64031) := X"AE020008";
        ram_buffer(64032) := X"8602000C";
        ram_buffer(64033) := X"00000000";
        ram_buffer(64034) := X"3042FFFF";
        ram_buffer(64035) := X"30420008";
        ram_buffer(64036) := X"10400005";
        ram_buffer(64037) := X"00000000";
        ram_buffer(64038) := X"8E020010";
        ram_buffer(64039) := X"00000000";
        ram_buffer(64040) := X"1440000A";
        ram_buffer(64041) := X"00000000";
        ram_buffer(64042) := X"02002821";
        ram_buffer(64043) := X"8FC40030";
        ram_buffer(64044) := X"0C02ACF1";
        ram_buffer(64045) := X"00000000";
        ram_buffer(64046) := X"10400004";
        ram_buffer(64047) := X"00000000";
        ram_buffer(64048) := X"2402FFFF";
        ram_buffer(64049) := X"10000049";
        ram_buffer(64050) := X"00000000";
        ram_buffer(64051) := X"325200FF";
        ram_buffer(64052) := X"8602000C";
        ram_buffer(64053) := X"00000000";
        ram_buffer(64054) := X"3042FFFF";
        ram_buffer(64055) := X"30422000";
        ram_buffer(64056) := X"1440000B";
        ram_buffer(64057) := X"00000000";
        ram_buffer(64058) := X"8602000C";
        ram_buffer(64059) := X"00000000";
        ram_buffer(64060) := X"34422000";
        ram_buffer(64061) := X"00021400";
        ram_buffer(64062) := X"00021403";
        ram_buffer(64063) := X"A602000C";
        ram_buffer(64064) := X"8E030064";
        ram_buffer(64065) := X"2402DFFF";
        ram_buffer(64066) := X"00621024";
        ram_buffer(64067) := X"AE020064";
        ram_buffer(64068) := X"8E020000";
        ram_buffer(64069) := X"00000000";
        ram_buffer(64070) := X"00401821";
        ram_buffer(64071) := X"8E020010";
        ram_buffer(64072) := X"00000000";
        ram_buffer(64073) := X"00628823";
        ram_buffer(64074) := X"8E020014";
        ram_buffer(64075) := X"00000000";
        ram_buffer(64076) := X"0222102A";
        ram_buffer(64077) := X"1440000B";
        ram_buffer(64078) := X"00000000";
        ram_buffer(64079) := X"02002821";
        ram_buffer(64080) := X"8FC40030";
        ram_buffer(64081) := X"0C026EE1";
        ram_buffer(64082) := X"00000000";
        ram_buffer(64083) := X"10400004";
        ram_buffer(64084) := X"00000000";
        ram_buffer(64085) := X"2402FFFF";
        ram_buffer(64086) := X"10000024";
        ram_buffer(64087) := X"00000000";
        ram_buffer(64088) := X"00008821";
        ram_buffer(64089) := X"8E020008";
        ram_buffer(64090) := X"00000000";
        ram_buffer(64091) := X"2442FFFF";
        ram_buffer(64092) := X"AE020008";
        ram_buffer(64093) := X"8E020000";
        ram_buffer(64094) := X"00000000";
        ram_buffer(64095) := X"24430001";
        ram_buffer(64096) := X"AE030000";
        ram_buffer(64097) := X"324300FF";
        ram_buffer(64098) := X"A0430000";
        ram_buffer(64099) := X"26310001";
        ram_buffer(64100) := X"8E020014";
        ram_buffer(64101) := X"00000000";
        ram_buffer(64102) := X"1222000A";
        ram_buffer(64103) := X"00000000";
        ram_buffer(64104) := X"8602000C";
        ram_buffer(64105) := X"00000000";
        ram_buffer(64106) := X"3042FFFF";
        ram_buffer(64107) := X"30420001";
        ram_buffer(64108) := X"1040000D";
        ram_buffer(64109) := X"00000000";
        ram_buffer(64110) := X"2402000A";
        ram_buffer(64111) := X"1642000A";
        ram_buffer(64112) := X"00000000";
        ram_buffer(64113) := X"02002821";
        ram_buffer(64114) := X"8FC40030";
        ram_buffer(64115) := X"0C026EE1";
        ram_buffer(64116) := X"00000000";
        ram_buffer(64117) := X"10400004";
        ram_buffer(64118) := X"00000000";
        ram_buffer(64119) := X"2402FFFF";
        ram_buffer(64120) := X"10000002";
        ram_buffer(64121) := X"00000000";
        ram_buffer(64122) := X"02401021";
        ram_buffer(64123) := X"03C0E821";
        ram_buffer(64124) := X"8FBF002C";
        ram_buffer(64125) := X"8FBE0028";
        ram_buffer(64126) := X"8FB20024";
        ram_buffer(64127) := X"8FB10020";
        ram_buffer(64128) := X"8FB0001C";
        ram_buffer(64129) := X"27BD0030";
        ram_buffer(64130) := X"03E00008";
        ram_buffer(64131) := X"00000000";
        ram_buffer(64132) := X"27BDFFE8";
        ram_buffer(64133) := X"AFBF0014";
        ram_buffer(64134) := X"AFBE0010";
        ram_buffer(64135) := X"03A0F021";
        ram_buffer(64136) := X"00801821";
        ram_buffer(64137) := X"00A02021";
        ram_buffer(64138) := X"8F828098";
        ram_buffer(64139) := X"00803021";
        ram_buffer(64140) := X"00602821";
        ram_buffer(64141) := X"00402021";
        ram_buffer(64142) := X"0C02FA03";
        ram_buffer(64143) := X"00000000";
        ram_buffer(64144) := X"03C0E821";
        ram_buffer(64145) := X"8FBF0014";
        ram_buffer(64146) := X"8FBE0010";
        ram_buffer(64147) := X"27BD0018";
        ram_buffer(64148) := X"03E00008";
        ram_buffer(64149) := X"00000000";
        ram_buffer(64150) := X"27BDFFC8";
        ram_buffer(64151) := X"AFBF0034";
        ram_buffer(64152) := X"AFBE0030";
        ram_buffer(64153) := X"AFB0002C";
        ram_buffer(64154) := X"03A0F021";
        ram_buffer(64155) := X"AFC40038";
        ram_buffer(64156) := X"AFC5003C";
        ram_buffer(64157) := X"AFC60040";
        ram_buffer(64158) := X"AFC70044";
        ram_buffer(64159) := X"AFC00018";
        ram_buffer(64160) := X"8FC2003C";
        ram_buffer(64161) := X"00000000";
        ram_buffer(64162) := X"14400012";
        ram_buffer(64163) := X"00000000";
        ram_buffer(64164) := X"8F908198";
        ram_buffer(64165) := X"0C02BAFF";
        ram_buffer(64166) := X"00000000";
        ram_buffer(64167) := X"00402021";
        ram_buffer(64168) := X"27C3001C";
        ram_buffer(64169) := X"8FC20044";
        ram_buffer(64170) := X"00000000";
        ram_buffer(64171) := X"AFA20010";
        ram_buffer(64172) := X"00803821";
        ram_buffer(64173) := X"00003021";
        ram_buffer(64174) := X"00602821";
        ram_buffer(64175) := X"8FC40038";
        ram_buffer(64176) := X"0200F809";
        ram_buffer(64177) := X"00000000";
        ram_buffer(64178) := X"AFC20018";
        ram_buffer(64179) := X"1000000F";
        ram_buffer(64180) := X"00000000";
        ram_buffer(64181) := X"8F908198";
        ram_buffer(64182) := X"0C02BAFF";
        ram_buffer(64183) := X"00000000";
        ram_buffer(64184) := X"00401821";
        ram_buffer(64185) := X"8FC20044";
        ram_buffer(64186) := X"00000000";
        ram_buffer(64187) := X"AFA20010";
        ram_buffer(64188) := X"00603821";
        ram_buffer(64189) := X"8FC60040";
        ram_buffer(64190) := X"8FC5003C";
        ram_buffer(64191) := X"8FC40038";
        ram_buffer(64192) := X"0200F809";
        ram_buffer(64193) := X"00000000";
        ram_buffer(64194) := X"AFC20018";
        ram_buffer(64195) := X"8FC30018";
        ram_buffer(64196) := X"2402FFFF";
        ram_buffer(64197) := X"1462000A";
        ram_buffer(64198) := X"00000000";
        ram_buffer(64199) := X"8FC20044";
        ram_buffer(64200) := X"00000000";
        ram_buffer(64201) := X"AC400000";
        ram_buffer(64202) := X"8FC20038";
        ram_buffer(64203) := X"2403008A";
        ram_buffer(64204) := X"AC430000";
        ram_buffer(64205) := X"2402FFFF";
        ram_buffer(64206) := X"10000002";
        ram_buffer(64207) := X"00000000";
        ram_buffer(64208) := X"8FC20018";
        ram_buffer(64209) := X"03C0E821";
        ram_buffer(64210) := X"8FBF0034";
        ram_buffer(64211) := X"8FBE0030";
        ram_buffer(64212) := X"8FB0002C";
        ram_buffer(64213) := X"27BD0038";
        ram_buffer(64214) := X"03E00008";
        ram_buffer(64215) := X"00000000";
        ram_buffer(64216) := X"27BDFFC0";
        ram_buffer(64217) := X"AFBF003C";
        ram_buffer(64218) := X"AFBE0038";
        ram_buffer(64219) := X"AFB00034";
        ram_buffer(64220) := X"03A0F021";
        ram_buffer(64221) := X"AFC40040";
        ram_buffer(64222) := X"AFC50044";
        ram_buffer(64223) := X"AFC60048";
        ram_buffer(64224) := X"AFC00018";
        ram_buffer(64225) := X"8F828098";
        ram_buffer(64226) := X"00000000";
        ram_buffer(64227) := X"AFC2001C";
        ram_buffer(64228) := X"8FC20040";
        ram_buffer(64229) := X"00000000";
        ram_buffer(64230) := X"14400012";
        ram_buffer(64231) := X"00000000";
        ram_buffer(64232) := X"8F908198";
        ram_buffer(64233) := X"0C02BAFF";
        ram_buffer(64234) := X"00000000";
        ram_buffer(64235) := X"00402021";
        ram_buffer(64236) := X"27C30020";
        ram_buffer(64237) := X"8FC20048";
        ram_buffer(64238) := X"00000000";
        ram_buffer(64239) := X"AFA20010";
        ram_buffer(64240) := X"00803821";
        ram_buffer(64241) := X"00003021";
        ram_buffer(64242) := X"00602821";
        ram_buffer(64243) := X"8FC4001C";
        ram_buffer(64244) := X"0200F809";
        ram_buffer(64245) := X"00000000";
        ram_buffer(64246) := X"AFC20018";
        ram_buffer(64247) := X"1000000F";
        ram_buffer(64248) := X"00000000";
        ram_buffer(64249) := X"8F908198";
        ram_buffer(64250) := X"0C02BAFF";
        ram_buffer(64251) := X"00000000";
        ram_buffer(64252) := X"00401821";
        ram_buffer(64253) := X"8FC20048";
        ram_buffer(64254) := X"00000000";
        ram_buffer(64255) := X"AFA20010";
        ram_buffer(64256) := X"00603821";
        ram_buffer(64257) := X"8FC60044";
        ram_buffer(64258) := X"8FC50040";
        ram_buffer(64259) := X"8FC4001C";
        ram_buffer(64260) := X"0200F809";
        ram_buffer(64261) := X"00000000";
        ram_buffer(64262) := X"AFC20018";
        ram_buffer(64263) := X"8FC30018";
        ram_buffer(64264) := X"2402FFFF";
        ram_buffer(64265) := X"1462000A";
        ram_buffer(64266) := X"00000000";
        ram_buffer(64267) := X"8FC20048";
        ram_buffer(64268) := X"00000000";
        ram_buffer(64269) := X"AC400000";
        ram_buffer(64270) := X"8FC2001C";
        ram_buffer(64271) := X"2403008A";
        ram_buffer(64272) := X"AC430000";
        ram_buffer(64273) := X"2402FFFF";
        ram_buffer(64274) := X"10000002";
        ram_buffer(64275) := X"00000000";
        ram_buffer(64276) := X"8FC20018";
        ram_buffer(64277) := X"03C0E821";
        ram_buffer(64278) := X"8FBF003C";
        ram_buffer(64279) := X"8FBE0038";
        ram_buffer(64280) := X"8FB00034";
        ram_buffer(64281) := X"27BD0040";
        ram_buffer(64282) := X"03E00008";
        ram_buffer(64283) := X"00000000";
        ram_buffer(64284) := X"27BDFFD8";
        ram_buffer(64285) := X"AFBF0024";
        ram_buffer(64286) := X"AFBE0020";
        ram_buffer(64287) := X"AFB0001C";
        ram_buffer(64288) := X"03A0F021";
        ram_buffer(64289) := X"AFC40028";
        ram_buffer(64290) := X"AFC5002C";
        ram_buffer(64291) := X"AFC60030";
        ram_buffer(64292) := X"AFC70034";
        ram_buffer(64293) := X"8F908198";
        ram_buffer(64294) := X"0C02BAFF";
        ram_buffer(64295) := X"00000000";
        ram_buffer(64296) := X"00401821";
        ram_buffer(64297) := X"8FC20034";
        ram_buffer(64298) := X"00000000";
        ram_buffer(64299) := X"AFA20010";
        ram_buffer(64300) := X"00603821";
        ram_buffer(64301) := X"8FC60030";
        ram_buffer(64302) := X"8FC5002C";
        ram_buffer(64303) := X"8FC40028";
        ram_buffer(64304) := X"0200F809";
        ram_buffer(64305) := X"00000000";
        ram_buffer(64306) := X"03C0E821";
        ram_buffer(64307) := X"8FBF0024";
        ram_buffer(64308) := X"8FBE0020";
        ram_buffer(64309) := X"8FB0001C";
        ram_buffer(64310) := X"27BD0028";
        ram_buffer(64311) := X"03E00008";
        ram_buffer(64312) := X"00000000";
        ram_buffer(64313) := X"27BDFFF0";
        ram_buffer(64314) := X"AFBE000C";
        ram_buffer(64315) := X"03A0F021";
        ram_buffer(64316) := X"AFC40010";
        ram_buffer(64317) := X"AFC50014";
        ram_buffer(64318) := X"AFC60018";
        ram_buffer(64319) := X"AFC7001C";
        ram_buffer(64320) := X"8FC20018";
        ram_buffer(64321) := X"00000000";
        ram_buffer(64322) := X"AFC20000";
        ram_buffer(64323) := X"8FC20014";
        ram_buffer(64324) := X"00000000";
        ram_buffer(64325) := X"14400004";
        ram_buffer(64326) := X"00000000";
        ram_buffer(64327) := X"00001021";
        ram_buffer(64328) := X"10000014";
        ram_buffer(64329) := X"00000000";
        ram_buffer(64330) := X"8FC20000";
        ram_buffer(64331) := X"00000000";
        ram_buffer(64332) := X"2C420100";
        ram_buffer(64333) := X"14400007";
        ram_buffer(64334) := X"00000000";
        ram_buffer(64335) := X"8FC20010";
        ram_buffer(64336) := X"2403008A";
        ram_buffer(64337) := X"AC430000";
        ram_buffer(64338) := X"2402FFFF";
        ram_buffer(64339) := X"10000009";
        ram_buffer(64340) := X"00000000";
        ram_buffer(64341) := X"8FC20000";
        ram_buffer(64342) := X"00000000";
        ram_buffer(64343) := X"00021E00";
        ram_buffer(64344) := X"00031E03";
        ram_buffer(64345) := X"8FC20014";
        ram_buffer(64346) := X"00000000";
        ram_buffer(64347) := X"A0430000";
        ram_buffer(64348) := X"24020001";
        ram_buffer(64349) := X"03C0E821";
        ram_buffer(64350) := X"8FBE000C";
        ram_buffer(64351) := X"27BD0010";
        ram_buffer(64352) := X"03E00008";
        ram_buffer(64353) := X"00000000";
        ram_buffer(64354) := X"3C04100D";
        ram_buffer(64355) := X"27BDFFE8";
        ram_buffer(64356) := X"AFBF0014";
        ram_buffer(64357) := X"0C028186";
        ram_buffer(64358) := X"2484B390";
        ram_buffer(64359) := X"1000FFFF";
        ram_buffer(64360) := X"00000000";
        ram_buffer(64361) := X"27BDFFE8";
        ram_buffer(64362) := X"AFB00010";
        ram_buffer(64363) := X"3C10100D";
        ram_buffer(64364) := X"000420C0";
        ram_buffer(64365) := X"2610DAC4";
        ram_buffer(64366) := X"AFBF0014";
        ram_buffer(64367) := X"00908021";
        ram_buffer(64368) := X"82020000";
        ram_buffer(64369) := X"00000000";
        ram_buffer(64370) := X"1040000A";
        ram_buffer(64371) := X"00000000";
        ram_buffer(64372) := X"8E040004";
        ram_buffer(64373) := X"0C03013B";
        ram_buffer(64374) := X"00000000";
        ram_buffer(64375) := X"A2000000";
        ram_buffer(64376) := X"00001021";
        ram_buffer(64377) := X"8FBF0014";
        ram_buffer(64378) := X"8FB00010";
        ram_buffer(64379) := X"03E00008";
        ram_buffer(64380) := X"27BD0018";
        ram_buffer(64381) := X"0C030730";
        ram_buffer(64382) := X"00000000";
        ram_buffer(64383) := X"24030009";
        ram_buffer(64384) := X"AC430000";
        ram_buffer(64385) := X"1000FFF7";
        ram_buffer(64386) := X"2402FFFF";
        ram_buffer(64387) := X"27BDFFE8";
        ram_buffer(64388) := X"2C820003";
        ram_buffer(64389) := X"14400021";
        ram_buffer(64390) := X"AFBF0014";
        ram_buffer(64391) := X"3C02100D";
        ram_buffer(64392) := X"2442DAC4";
        ram_buffer(64393) := X"000420C0";
        ram_buffer(64394) := X"00822021";
        ram_buffer(64395) := X"80830000";
        ram_buffer(64396) := X"24020001";
        ram_buffer(64397) := X"1462001F";
        ram_buffer(64398) := X"00000000";
        ram_buffer(64399) := X"8C820004";
        ram_buffer(64400) := X"00000000";
        ram_buffer(64401) := X"10400021";
        ram_buffer(64402) := X"00000000";
        ram_buffer(64403) := X"94440038";
        ram_buffer(64404) := X"8C430030";
        ram_buffer(64405) := X"ACA4002C";
        ram_buffer(64406) := X"ACA30010";
        ram_buffer(64407) := X"90420034";
        ram_buffer(64408) := X"00000000";
        ram_buffer(64409) := X"14400008";
        ram_buffer(64410) := X"24024000";
        ram_buffer(64411) := X"34028000";
        ram_buffer(64412) := X"ACA20004";
        ram_buffer(64413) := X"00001021";
        ram_buffer(64414) := X"8FBF0014";
        ram_buffer(64415) := X"00000000";
        ram_buffer(64416) := X"03E00008";
        ram_buffer(64417) := X"27BD0018";
        ram_buffer(64418) := X"8FBF0014";
        ram_buffer(64419) := X"ACA20004";
        ram_buffer(64420) := X"00001021";
        ram_buffer(64421) := X"03E00008";
        ram_buffer(64422) := X"27BD0018";
        ram_buffer(64423) := X"8FBF0014";
        ram_buffer(64424) := X"24022000";
        ram_buffer(64425) := X"ACA20004";
        ram_buffer(64426) := X"00001021";
        ram_buffer(64427) := X"03E00008";
        ram_buffer(64428) := X"27BD0018";
        ram_buffer(64429) := X"0C030730";
        ram_buffer(64430) := X"00000000";
        ram_buffer(64431) := X"24030009";
        ram_buffer(64432) := X"AC430000";
        ram_buffer(64433) := X"1000FFEC";
        ram_buffer(64434) := X"2402FFFF";
        ram_buffer(64435) := X"0C030730";
        ram_buffer(64436) := X"00000000";
        ram_buffer(64437) := X"24030002";
        ram_buffer(64438) := X"AC430000";
        ram_buffer(64439) := X"1000FFE6";
        ram_buffer(64440) := X"2402FFFF";
        ram_buffer(64441) := X"03E00008";
        ram_buffer(64442) := X"24020001";
        ram_buffer(64443) := X"2C820003";
        ram_buffer(64444) := X"14400012";
        ram_buffer(64445) := X"000420C0";
        ram_buffer(64446) := X"3C02100D";
        ram_buffer(64447) := X"27BDFFE8";
        ram_buffer(64448) := X"2442DAC4";
        ram_buffer(64449) := X"00822021";
        ram_buffer(64450) := X"AFBF0014";
        ram_buffer(64451) := X"80830000";
        ram_buffer(64452) := X"24020001";
        ram_buffer(64453) := X"1062000B";
        ram_buffer(64454) := X"00000000";
        ram_buffer(64455) := X"0C030730";
        ram_buffer(64456) := X"00000000";
        ram_buffer(64457) := X"8FBF0014";
        ram_buffer(64458) := X"24030009";
        ram_buffer(64459) := X"AC430000";
        ram_buffer(64460) := X"00001021";
        ram_buffer(64461) := X"03E00008";
        ram_buffer(64462) := X"27BD0018";
        ram_buffer(64463) := X"03E00008";
        ram_buffer(64464) := X"24020001";
        ram_buffer(64465) := X"0C030730";
        ram_buffer(64466) := X"00000000";
        ram_buffer(64467) := X"8FBF0014";
        ram_buffer(64468) := X"24030019";
        ram_buffer(64469) := X"AC430000";
        ram_buffer(64470) := X"00001021";
        ram_buffer(64471) := X"03E00008";
        ram_buffer(64472) := X"27BD0018";
        ram_buffer(64473) := X"27BDFFE8";
        ram_buffer(64474) := X"2C820003";
        ram_buffer(64475) := X"14400015";
        ram_buffer(64476) := X"AFBF0014";
        ram_buffer(64477) := X"3C02100D";
        ram_buffer(64478) := X"2442DAC4";
        ram_buffer(64479) := X"000420C0";
        ram_buffer(64480) := X"00822021";
        ram_buffer(64481) := X"80830000";
        ram_buffer(64482) := X"24020001";
        ram_buffer(64483) := X"14620005";
        ram_buffer(64484) := X"00000000";
        ram_buffer(64485) := X"8FBF0014";
        ram_buffer(64486) := X"8C840004";
        ram_buffer(64487) := X"0802FFF2";
        ram_buffer(64488) := X"27BD0018";
        ram_buffer(64489) := X"0C030730";
        ram_buffer(64490) := X"00000000";
        ram_buffer(64491) := X"24030009";
        ram_buffer(64492) := X"AC430000";
        ram_buffer(64493) := X"8FBF0014";
        ram_buffer(64494) := X"2402FFFF";
        ram_buffer(64495) := X"03E00008";
        ram_buffer(64496) := X"27BD0018";
        ram_buffer(64497) := X"0C030730";
        ram_buffer(64498) := X"00000000";
        ram_buffer(64499) := X"2403001D";
        ram_buffer(64500) := X"1000FFF8";
        ram_buffer(64501) := X"AC430000";
        ram_buffer(64502) := X"27BDFFE0";
        ram_buffer(64503) := X"3C03100D";
        ram_buffer(64504) := X"2463DADC";
        ram_buffer(64505) := X"AFB00018";
        ram_buffer(64506) := X"AFA60028";
        ram_buffer(64507) := X"AFBF001C";
        ram_buffer(64508) := X"AFA7002C";
        ram_buffer(64509) := X"24100003";
        ram_buffer(64510) := X"10000004";
        ram_buffer(64511) := X"24060080";
        ram_buffer(64512) := X"26100001";
        ram_buffer(64513) := X"12060023";
        ram_buffer(64514) := X"00000000";
        ram_buffer(64515) := X"80620000";
        ram_buffer(64516) := X"00000000";
        ram_buffer(64517) := X"1440FFFA";
        ram_buffer(64518) := X"24630008";
        ram_buffer(64519) := X"30A20001";
        ram_buffer(64520) := X"1440001A";
        ram_buffer(64521) := X"24020077";
        ram_buffer(64522) := X"24020072";
        ram_buffer(64523) := X"A3A20010";
        ram_buffer(64524) := X"30A20002";
        ram_buffer(64525) := X"10400002";
        ram_buffer(64526) := X"24020077";
        ram_buffer(64527) := X"A3A20010";
        ram_buffer(64528) := X"30A50008";
        ram_buffer(64529) := X"10A00002";
        ram_buffer(64530) := X"24020061";
        ram_buffer(64531) := X"A3A20010";
        ram_buffer(64532) := X"0C0302B9";
        ram_buffer(64533) := X"27A50010";
        ram_buffer(64534) := X"10400012";
        ram_buffer(64535) := X"3C03100D";
        ram_buffer(64536) := X"001020C0";
        ram_buffer(64537) := X"2463DAC4";
        ram_buffer(64538) := X"00831821";
        ram_buffer(64539) := X"24040001";
        ram_buffer(64540) := X"A0640000";
        ram_buffer(64541) := X"8FBF001C";
        ram_buffer(64542) := X"AC620004";
        ram_buffer(64543) := X"02001021";
        ram_buffer(64544) := X"8FB00018";
        ram_buffer(64545) := X"03E00008";
        ram_buffer(64546) := X"27BD0020";
        ram_buffer(64547) := X"1000FFE8";
        ram_buffer(64548) := X"A3A20010";
        ram_buffer(64549) := X"0C030730";
        ram_buffer(64550) := X"00000000";
        ram_buffer(64551) := X"24030017";
        ram_buffer(64552) := X"AC430000";
        ram_buffer(64553) := X"8FBF001C";
        ram_buffer(64554) := X"8FB00018";
        ram_buffer(64555) := X"2402FFFF";
        ram_buffer(64556) := X"03E00008";
        ram_buffer(64557) := X"27BD0020";
        ram_buffer(64558) := X"27BDFFD8";
        ram_buffer(64559) := X"AFB20018";
        ram_buffer(64560) := X"AFB00010";
        ram_buffer(64561) := X"AFBF0024";
        ram_buffer(64562) := X"AFB40020";
        ram_buffer(64563) := X"AFB3001C";
        ram_buffer(64564) := X"AFB10014";
        ram_buffer(64565) := X"00A08021";
        ram_buffer(64566) := X"10800025";
        ram_buffer(64567) := X"00C09021";
        ram_buffer(64568) := X"04800010";
        ram_buffer(64569) := X"28820003";
        ram_buffer(64570) := X"1040000F";
        ram_buffer(64571) := X"3C02100D";
        ram_buffer(64572) := X"0C030730";
        ram_buffer(64573) := X"2414FFFF";
        ram_buffer(64574) := X"24030016";
        ram_buffer(64575) := X"AC430000";
        ram_buffer(64576) := X"8FBF0024";
        ram_buffer(64577) := X"02801021";
        ram_buffer(64578) := X"8FB3001C";
        ram_buffer(64579) := X"8FB40020";
        ram_buffer(64580) := X"8FB20018";
        ram_buffer(64581) := X"8FB10014";
        ram_buffer(64582) := X"8FB00010";
        ram_buffer(64583) := X"03E00008";
        ram_buffer(64584) := X"27BD0028";
        ram_buffer(64585) := X"3C02100D";
        ram_buffer(64586) := X"2442DAC4";
        ram_buffer(64587) := X"000420C0";
        ram_buffer(64588) := X"00822021";
        ram_buffer(64589) := X"80830000";
        ram_buffer(64590) := X"24020001";
        ram_buffer(64591) := X"14620024";
        ram_buffer(64592) := X"02403021";
        ram_buffer(64593) := X"8C870004";
        ram_buffer(64594) := X"8FBF0024";
        ram_buffer(64595) := X"8FB40020";
        ram_buffer(64596) := X"8FB3001C";
        ram_buffer(64597) := X"8FB10014";
        ram_buffer(64598) := X"02002021";
        ram_buffer(64599) := X"8FB20018";
        ram_buffer(64600) := X"8FB00010";
        ram_buffer(64601) := X"24050001";
        ram_buffer(64602) := X"0802FF53";
        ram_buffer(64603) := X"27BD0028";
        ram_buffer(64604) := X"10C0001C";
        ram_buffer(64605) := X"00008821";
        ram_buffer(64606) := X"00C0A021";
        ram_buffer(64607) := X"10000004";
        ram_buffer(64608) := X"2413000A";
        ram_buffer(64609) := X"26310001";
        ram_buffer(64610) := X"1232FFDD";
        ram_buffer(64611) := X"26100001";
        ram_buffer(64612) := X"0C030702";
        ram_buffer(64613) := X"00000000";
        ram_buffer(64614) := X"00021600";
        ram_buffer(64615) := X"00021603";
        ram_buffer(64616) := X"1453FFF8";
        ram_buffer(64617) := X"A2020000";
        ram_buffer(64618) := X"8FBF0024";
        ram_buffer(64619) := X"0220A021";
        ram_buffer(64620) := X"02801021";
        ram_buffer(64621) := X"8FB3001C";
        ram_buffer(64622) := X"8FB40020";
        ram_buffer(64623) := X"8FB20018";
        ram_buffer(64624) := X"8FB10014";
        ram_buffer(64625) := X"8FB00010";
        ram_buffer(64626) := X"03E00008";
        ram_buffer(64627) := X"27BD0028";
        ram_buffer(64628) := X"0C030730";
        ram_buffer(64629) := X"2414FFFF";
        ram_buffer(64630) := X"24030009";
        ram_buffer(64631) := X"1000FFC8";
        ram_buffer(64632) := X"AC430000";
        ram_buffer(64633) := X"1000FFC6";
        ram_buffer(64634) := X"0000A021";
        ram_buffer(64635) := X"8F8281E0";
        ram_buffer(64636) := X"27BDFFE0";
        ram_buffer(64637) := X"AFBF001C";
        ram_buffer(64638) := X"AFB10018";
        ram_buffer(64639) := X"1040001C";
        ram_buffer(64640) := X"AFB00014";
        ram_buffer(64641) := X"80430000";
        ram_buffer(64642) := X"3C050FFF";
        ram_buffer(64643) := X"34A5FFFF";
        ram_buffer(64644) := X"00641821";
        ram_buffer(64645) := X"00651824";
        ram_buffer(64646) := X"3C0501FF";
        ram_buffer(64647) := X"34A5F001";
        ram_buffer(64648) := X"0065182A";
        ram_buffer(64649) := X"10600007";
        ram_buffer(64650) := X"00442021";
        ram_buffer(64651) := X"8FBF001C";
        ram_buffer(64652) := X"8FB10018";
        ram_buffer(64653) := X"8FB00014";
        ram_buffer(64654) := X"AF8481E0";
        ram_buffer(64655) := X"03E00008";
        ram_buffer(64656) := X"27BD0020";
        ram_buffer(64657) := X"3C10100D";
        ram_buffer(64658) := X"3C11100D";
        ram_buffer(64659) := X"2610B3A0";
        ram_buffer(64660) := X"2631B3B3";
        ram_buffer(64661) := X"82040000";
        ram_buffer(64662) := X"0C0306B6";
        ram_buffer(64663) := X"26100001";
        ram_buffer(64664) := X"1611FFFC";
        ram_buffer(64665) := X"00000000";
        ram_buffer(64666) := X"1000FFFF";
        ram_buffer(64667) := X"00000000";
        ram_buffer(64668) := X"3C021020";
        ram_buffer(64669) := X"AF8281E0";
        ram_buffer(64670) := X"80420000";
        ram_buffer(64671) := X"3C030FFF";
        ram_buffer(64672) := X"3463FFFF";
        ram_buffer(64673) := X"00441021";
        ram_buffer(64674) := X"00431024";
        ram_buffer(64675) := X"3C0301FF";
        ram_buffer(64676) := X"3463F001";
        ram_buffer(64677) := X"0043102A";
        ram_buffer(64678) := X"1040FFEB";
        ram_buffer(64679) := X"3C10100D";
        ram_buffer(64680) := X"3C021020";
        ram_buffer(64681) := X"8FBF001C";
        ram_buffer(64682) := X"00442021";
        ram_buffer(64683) := X"8FB10018";
        ram_buffer(64684) := X"8FB00014";
        ram_buffer(64685) := X"AF8481E0";
        ram_buffer(64686) := X"03E00008";
        ram_buffer(64687) := X"27BD0020";
        ram_buffer(64688) := X"27BDFE70";
        ram_buffer(64689) := X"27A7015C";
        ram_buffer(64690) := X"27A60120";
        ram_buffer(64691) := X"AFB00188";
        ram_buffer(64692) := X"00A08021";
        ram_buffer(64693) := X"00802821";
        ram_buffer(64694) := X"AFBF018C";
        ram_buffer(64695) := X"0C030030";
        ram_buffer(64696) := X"27A40010";
        ram_buffer(64697) := X"14400013";
        ram_buffer(64698) := X"00000000";
        ram_buffer(64699) := X"97A40158";
        ram_buffer(64700) := X"93A30154";
        ram_buffer(64701) := X"AE04002C";
        ram_buffer(64702) := X"8FA40150";
        ram_buffer(64703) := X"14600007";
        ram_buffer(64704) := X"AE040010";
        ram_buffer(64705) := X"34038000";
        ram_buffer(64706) := X"AE030004";
        ram_buffer(64707) := X"8FBF018C";
        ram_buffer(64708) := X"8FB00188";
        ram_buffer(64709) := X"03E00008";
        ram_buffer(64710) := X"27BD0190";
        ram_buffer(64711) := X"8FBF018C";
        ram_buffer(64712) := X"24034000";
        ram_buffer(64713) := X"AE030004";
        ram_buffer(64714) := X"8FB00188";
        ram_buffer(64715) := X"03E00008";
        ram_buffer(64716) := X"27BD0190";
        ram_buffer(64717) := X"0C030730";
        ram_buffer(64718) := X"00000000";
        ram_buffer(64719) := X"24030002";
        ram_buffer(64720) := X"AC430000";
        ram_buffer(64721) := X"1000FFF1";
        ram_buffer(64722) := X"2402FFFF";
        ram_buffer(64723) := X"27BDFFE8";
        ram_buffer(64724) := X"AFBF0014";
        ram_buffer(64725) := X"0C0301F5";
        ram_buffer(64726) := X"00000000";
        ram_buffer(64727) := X"14400005";
        ram_buffer(64728) := X"00000000";
        ram_buffer(64729) := X"8FBF0014";
        ram_buffer(64730) := X"00000000";
        ram_buffer(64731) := X"03E00008";
        ram_buffer(64732) := X"27BD0018";
        ram_buffer(64733) := X"0C030730";
        ram_buffer(64734) := X"00000000";
        ram_buffer(64735) := X"24030002";
        ram_buffer(64736) := X"AC430000";
        ram_buffer(64737) := X"1000FFF7";
        ram_buffer(64738) := X"2402FFFF";
        ram_buffer(64739) := X"27BDFFE0";
        ram_buffer(64740) := X"AFBF001C";
        ram_buffer(64741) := X"AFB20018";
        ram_buffer(64742) := X"AFB10014";
        ram_buffer(64743) := X"10800026";
        ram_buffer(64744) := X"AFB00010";
        ram_buffer(64745) := X"00A08021";
        ram_buffer(64746) := X"04800012";
        ram_buffer(64747) := X"00C09021";
        ram_buffer(64748) := X"28820003";
        ram_buffer(64749) := X"10400010";
        ram_buffer(64750) := X"3C02100D";
        ram_buffer(64751) := X"10C00006";
        ram_buffer(64752) := X"00A68821";
        ram_buffer(64753) := X"82040000";
        ram_buffer(64754) := X"0C0306B6";
        ram_buffer(64755) := X"26100001";
        ram_buffer(64756) := X"1630FFFC";
        ram_buffer(64757) := X"00000000";
        ram_buffer(64758) := X"02401021";
        ram_buffer(64759) := X"8FBF001C";
        ram_buffer(64760) := X"8FB20018";
        ram_buffer(64761) := X"8FB10014";
        ram_buffer(64762) := X"8FB00010";
        ram_buffer(64763) := X"03E00008";
        ram_buffer(64764) := X"27BD0020";
        ram_buffer(64765) := X"3C02100D";
        ram_buffer(64766) := X"2442DAC4";
        ram_buffer(64767) := X"000420C0";
        ram_buffer(64768) := X"00822021";
        ram_buffer(64769) := X"80830000";
        ram_buffer(64770) := X"24020001";
        ram_buffer(64771) := X"14620015";
        ram_buffer(64772) := X"02403021";
        ram_buffer(64773) := X"8C870004";
        ram_buffer(64774) := X"8FBF001C";
        ram_buffer(64775) := X"8FB10014";
        ram_buffer(64776) := X"02002021";
        ram_buffer(64777) := X"8FB20018";
        ram_buffer(64778) := X"8FB00010";
        ram_buffer(64779) := X"24050001";
        ram_buffer(64780) := X"0802FF99";
        ram_buffer(64781) := X"27BD0020";
        ram_buffer(64782) := X"0C030730";
        ram_buffer(64783) := X"00000000";
        ram_buffer(64784) := X"8FBF001C";
        ram_buffer(64785) := X"24030016";
        ram_buffer(64786) := X"AC430000";
        ram_buffer(64787) := X"8FB20018";
        ram_buffer(64788) := X"8FB10014";
        ram_buffer(64789) := X"8FB00010";
        ram_buffer(64790) := X"2402FFFF";
        ram_buffer(64791) := X"03E00008";
        ram_buffer(64792) := X"27BD0020";
        ram_buffer(64793) := X"0C030730";
        ram_buffer(64794) := X"00000000";
        ram_buffer(64795) := X"24030009";
        ram_buffer(64796) := X"AC430000";
        ram_buffer(64797) := X"1000FFD9";
        ram_buffer(64798) := X"2402FFFF";
        ram_buffer(64799) := X"27BDFFE8";
        ram_buffer(64800) := X"AFBF0014";
        ram_buffer(64801) := X"0C030730";
        ram_buffer(64802) := X"00000000";
        ram_buffer(64803) := X"8FBF0014";
        ram_buffer(64804) := X"24030016";
        ram_buffer(64805) := X"AC430000";
        ram_buffer(64806) := X"2402FFFF";
        ram_buffer(64807) := X"03E00008";
        ram_buffer(64808) := X"27BD0018";
        ram_buffer(64809) := X"27BDFFB0";
        ram_buffer(64810) := X"AFB60040";
        ram_buffer(64811) := X"AFB5003C";
        ram_buffer(64812) := X"AFBF004C";
        ram_buffer(64813) := X"AFBE0048";
        ram_buffer(64814) := X"AFB70044";
        ram_buffer(64815) := X"AFB40038";
        ram_buffer(64816) := X"AFB30034";
        ram_buffer(64817) := X"AFB20030";
        ram_buffer(64818) := X"AFB1002C";
        ram_buffer(64819) := X"AFB00028";
        ram_buffer(64820) := X"00A0B021";
        ram_buffer(64821) := X"10A00042";
        ram_buffer(64822) := X"0080A821";
        ram_buffer(64823) := X"8C8400CC";
        ram_buffer(64824) := X"00000000";
        ram_buffer(64825) := X"10800141";
        ram_buffer(64826) := X"00000000";
        ram_buffer(64827) := X"92A2003D";
        ram_buffer(64828) := X"00000000";
        ram_buffer(64829) := X"14400034";
        ram_buffer(64830) := X"00A08021";
        ram_buffer(64831) := X"2402FFFF";
        ram_buffer(64832) := X"1202000E";
        ram_buffer(64833) := X"00000000";
        ram_buffer(64834) := X"92A20037";
        ram_buffer(64835) := X"AEB00040";
        ram_buffer(64836) := X"14400124";
        ram_buffer(64837) := X"AEA00044";
        ram_buffer(64838) := X"AEB000CC";
        ram_buffer(64839) := X"16C00007";
        ram_buffer(64840) := X"00000000";
        ram_buffer(64841) := X"96A60038";
        ram_buffer(64842) := X"8EA400CC";
        ram_buffer(64843) := X"0C02801D";
        ram_buffer(64844) := X"240500FF";
        ram_buffer(64845) := X"24020001";
        ram_buffer(64846) := X"A2A2003D";
        ram_buffer(64847) := X"8FBF004C";
        ram_buffer(64848) := X"8FBE0048";
        ram_buffer(64849) := X"8FB70044";
        ram_buffer(64850) := X"8FB60040";
        ram_buffer(64851) := X"8FB5003C";
        ram_buffer(64852) := X"8FB40038";
        ram_buffer(64853) := X"8FB30034";
        ram_buffer(64854) := X"8FB20030";
        ram_buffer(64855) := X"8FB1002C";
        ram_buffer(64856) := X"8FB00028";
        ram_buffer(64857) := X"03E00008";
        ram_buffer(64858) := X"27BD0050";
        ram_buffer(64859) := X"24020028";
        ram_buffer(64860) := X"02602021";
        ram_buffer(64861) := X"0C027A4D";
        ram_buffer(64862) := X"AF8281E4";
        ram_buffer(64863) := X"12400115";
        ram_buffer(64864) := X"00000000";
        ram_buffer(64865) := X"92A30037";
        ram_buffer(64866) := X"00000000";
        ram_buffer(64867) := X"14600028";
        ram_buffer(64868) := X"24020028";
        ram_buffer(64869) := X"96A40038";
        ram_buffer(64870) := X"0C027A3D";
        ram_buffer(64871) := X"00000000";
        ram_buffer(64872) := X"00408021";
        ram_buffer(64873) := X"1200010B";
        ram_buffer(64874) := X"00000000";
        ram_buffer(64875) := X"8EA400CC";
        ram_buffer(64876) := X"00000000";
        ram_buffer(64877) := X"1080FFD2";
        ram_buffer(64878) := X"2402FFFF";
        ram_buffer(64879) := X"24020001";
        ram_buffer(64880) := X"AC900000";
        ram_buffer(64881) := X"A2A2003D";
        ram_buffer(64882) := X"92A20037";
        ram_buffer(64883) := X"00000000";
        ram_buffer(64884) := X"144000FB";
        ram_buffer(64885) := X"24060040";
        ram_buffer(64886) := X"1000FFC8";
        ram_buffer(64887) := X"A2A0003D";
        ram_buffer(64888) := X"90820037";
        ram_buffer(64889) := X"00000000";
        ram_buffer(64890) := X"1040FFEA";
        ram_buffer(64891) := X"3C03100D";
        ram_buffer(64892) := X"00602021";
        ram_buffer(64893) := X"2490D688";
        ram_buffer(64894) := X"3C04100D";
        ram_buffer(64895) := X"AFA40014";
        ram_buffer(64896) := X"3C04100D";
        ram_buffer(64897) := X"8F8281E4";
        ram_buffer(64898) := X"AFA40018";
        ram_buffer(64899) := X"3C04100D";
        ram_buffer(64900) := X"AFA4001C";
        ram_buffer(64901) := X"3C04100D";
        ram_buffer(64902) := X"AFA30010";
        ram_buffer(64903) := X"2484DA88";
        ram_buffer(64904) := X"28432000";
        ram_buffer(64905) := X"3C1E100D";
        ram_buffer(64906) := X"10600017";
        ram_buffer(64907) := X"AFA40020";
        ram_buffer(64908) := X"000228C3";
        ram_buffer(64909) := X"02051821";
        ram_buffer(64910) := X"90670000";
        ram_buffer(64911) := X"30460007";
        ram_buffer(64912) := X"00C71807";
        ram_buffer(64913) := X"30630001";
        ram_buffer(64914) := X"02002021";
        ram_buffer(64915) := X"10600009";
        ram_buffer(64916) := X"24082000";
        ram_buffer(64917) := X"100000C1";
        ram_buffer(64918) := X"24030001";
        ram_buffer(64919) := X"90670000";
        ram_buffer(64920) := X"00000000";
        ram_buffer(64921) := X"00C71807";
        ram_buffer(64922) := X"30630001";
        ram_buffer(64923) := X"146000BB";
        ram_buffer(64924) := X"24030001";
        ram_buffer(64925) := X"24420001";
        ram_buffer(64926) := X"000228C3";
        ram_buffer(64927) := X"02051821";
        ram_buffer(64928) := X"1448FFF6";
        ram_buffer(64929) := X"30460007";
        ram_buffer(64930) := X"8FA20014";
        ram_buffer(64931) := X"0C028186";
        ram_buffer(64932) := X"2444B3B4";
        ram_buffer(64933) := X"0C027A3D";
        ram_buffer(64934) := X"24040200";
        ram_buffer(64935) := X"104000CD";
        ram_buffer(64936) := X"00409821";
        ram_buffer(64937) := X"2417000F";
        ram_buffer(64938) := X"00009021";
        ram_buffer(64939) := X"10000041";
        ram_buffer(64940) := X"24110001";
        ram_buffer(64941) := X"000210C3";
        ram_buffer(64942) := X"02021021";
        ram_buffer(64943) := X"90420000";
        ram_buffer(64944) := X"00000000";
        ram_buffer(64945) := X"30420002";
        ram_buffer(64946) := X"14400058";
        ram_buffer(64947) := X"24060040";
        ram_buffer(64948) := X"26E2FFFB";
        ram_buffer(64949) := X"000210C3";
        ram_buffer(64950) := X"02021021";
        ram_buffer(64951) := X"90420000";
        ram_buffer(64952) := X"00000000";
        ram_buffer(64953) := X"30420004";
        ram_buffer(64954) := X"1440005C";
        ram_buffer(64955) := X"24060040";
        ram_buffer(64956) := X"26E2FFFC";
        ram_buffer(64957) := X"000210C3";
        ram_buffer(64958) := X"02021021";
        ram_buffer(64959) := X"90420000";
        ram_buffer(64960) := X"00000000";
        ram_buffer(64961) := X"30420008";
        ram_buffer(64962) := X"14400060";
        ram_buffer(64963) := X"24060040";
        ram_buffer(64964) := X"26E2FFFD";
        ram_buffer(64965) := X"000210C3";
        ram_buffer(64966) := X"02021021";
        ram_buffer(64967) := X"90420000";
        ram_buffer(64968) := X"00000000";
        ram_buffer(64969) := X"30420010";
        ram_buffer(64970) := X"14400064";
        ram_buffer(64971) := X"24060040";
        ram_buffer(64972) := X"26E2FFFE";
        ram_buffer(64973) := X"000210C3";
        ram_buffer(64974) := X"02021021";
        ram_buffer(64975) := X"90420000";
        ram_buffer(64976) := X"00000000";
        ram_buffer(64977) := X"30420020";
        ram_buffer(64978) := X"14400068";
        ram_buffer(64979) := X"24060040";
        ram_buffer(64980) := X"26E2FFFF";
        ram_buffer(64981) := X"000210C3";
        ram_buffer(64982) := X"02021021";
        ram_buffer(64983) := X"90420000";
        ram_buffer(64984) := X"00000000";
        ram_buffer(64985) := X"30420040";
        ram_buffer(64986) := X"1440006C";
        ram_buffer(64987) := X"24060040";
        ram_buffer(64988) := X"001710C3";
        ram_buffer(64989) := X"02021021";
        ram_buffer(64990) := X"90420000";
        ram_buffer(64991) := X"00000000";
        ram_buffer(64992) := X"30420080";
        ram_buffer(64993) := X"14400070";
        ram_buffer(64994) := X"24060040";
        ram_buffer(64995) := X"0C03069E";
        ram_buffer(64996) := X"02802021";
        ram_buffer(64997) := X"24060200";
        ram_buffer(64998) := X"02802821";
        ram_buffer(64999) := X"0C030698";
        ram_buffer(65000) := X"02602021";
        ram_buffer(65001) := X"26310001";
        ram_buffer(65002) := X"24020400";
        ram_buffer(65003) := X"1222FF6F";
        ram_buffer(65004) := X"26F70008";
        ram_buffer(65005) := X"2404002E";
        ram_buffer(65006) := X"0C030866";
        ram_buffer(65007) := X"0011A240";
        ram_buffer(65008) := X"24060200";
        ram_buffer(65009) := X"02802821";
        ram_buffer(65010) := X"0C03068E";
        ram_buffer(65011) := X"02602021";
        ram_buffer(65012) := X"24020001";
        ram_buffer(65013) := X"12220087";
        ram_buffer(65014) := X"001110C0";
        ram_buffer(65015) := X"000210C3";
        ram_buffer(65016) := X"02021021";
        ram_buffer(65017) := X"90420000";
        ram_buffer(65018) := X"00000000";
        ram_buffer(65019) := X"30420001";
        ram_buffer(65020) := X"1040FFB0";
        ram_buffer(65021) := X"26E2FFFA";
        ram_buffer(65022) := X"24060040";
        ram_buffer(65023) := X"240500FF";
        ram_buffer(65024) := X"0C02801D";
        ram_buffer(65025) := X"02602021";
        ram_buffer(65026) := X"26E2FFFA";
        ram_buffer(65027) := X"000210C3";
        ram_buffer(65028) := X"02021021";
        ram_buffer(65029) := X"90420000";
        ram_buffer(65030) := X"00000000";
        ram_buffer(65031) := X"30420002";
        ram_buffer(65032) := X"1040FFAB";
        ram_buffer(65033) := X"26520001";
        ram_buffer(65034) := X"24060040";
        ram_buffer(65035) := X"240500FF";
        ram_buffer(65036) := X"0C02801D";
        ram_buffer(65037) := X"26640040";
        ram_buffer(65038) := X"26E2FFFB";
        ram_buffer(65039) := X"000210C3";
        ram_buffer(65040) := X"02021021";
        ram_buffer(65041) := X"90420000";
        ram_buffer(65042) := X"00000000";
        ram_buffer(65043) := X"30420004";
        ram_buffer(65044) := X"1040FFA7";
        ram_buffer(65045) := X"26520001";
        ram_buffer(65046) := X"24060040";
        ram_buffer(65047) := X"240500FF";
        ram_buffer(65048) := X"0C02801D";
        ram_buffer(65049) := X"26640080";
        ram_buffer(65050) := X"26E2FFFC";
        ram_buffer(65051) := X"000210C3";
        ram_buffer(65052) := X"02021021";
        ram_buffer(65053) := X"90420000";
        ram_buffer(65054) := X"00000000";
        ram_buffer(65055) := X"30420008";
        ram_buffer(65056) := X"1040FFA3";
        ram_buffer(65057) := X"26520001";
        ram_buffer(65058) := X"24060040";
        ram_buffer(65059) := X"240500FF";
        ram_buffer(65060) := X"0C02801D";
        ram_buffer(65061) := X"266400C0";
        ram_buffer(65062) := X"26E2FFFD";
        ram_buffer(65063) := X"000210C3";
        ram_buffer(65064) := X"02021021";
        ram_buffer(65065) := X"90420000";
        ram_buffer(65066) := X"00000000";
        ram_buffer(65067) := X"30420010";
        ram_buffer(65068) := X"1040FF9F";
        ram_buffer(65069) := X"26520001";
        ram_buffer(65070) := X"24060040";
        ram_buffer(65071) := X"240500FF";
        ram_buffer(65072) := X"0C02801D";
        ram_buffer(65073) := X"26640100";
        ram_buffer(65074) := X"26E2FFFE";
        ram_buffer(65075) := X"000210C3";
        ram_buffer(65076) := X"02021021";
        ram_buffer(65077) := X"90420000";
        ram_buffer(65078) := X"00000000";
        ram_buffer(65079) := X"30420020";
        ram_buffer(65080) := X"1040FF9B";
        ram_buffer(65081) := X"26520001";
        ram_buffer(65082) := X"24060040";
        ram_buffer(65083) := X"240500FF";
        ram_buffer(65084) := X"0C02801D";
        ram_buffer(65085) := X"26640140";
        ram_buffer(65086) := X"26E2FFFF";
        ram_buffer(65087) := X"000210C3";
        ram_buffer(65088) := X"02021021";
        ram_buffer(65089) := X"90420000";
        ram_buffer(65090) := X"00000000";
        ram_buffer(65091) := X"30420040";
        ram_buffer(65092) := X"1040FF97";
        ram_buffer(65093) := X"26520001";
        ram_buffer(65094) := X"24060040";
        ram_buffer(65095) := X"240500FF";
        ram_buffer(65096) := X"0C02801D";
        ram_buffer(65097) := X"26640180";
        ram_buffer(65098) := X"001710C3";
        ram_buffer(65099) := X"02021021";
        ram_buffer(65100) := X"90420000";
        ram_buffer(65101) := X"00000000";
        ram_buffer(65102) := X"30420080";
        ram_buffer(65103) := X"1040FF93";
        ram_buffer(65104) := X"26520001";
        ram_buffer(65105) := X"24060040";
        ram_buffer(65106) := X"240500FF";
        ram_buffer(65107) := X"0C02801D";
        ram_buffer(65108) := X"266401C0";
        ram_buffer(65109) := X"1000FF8D";
        ram_buffer(65110) := X"26520001";
        ram_buffer(65111) := X"00C33004";
        ram_buffer(65112) := X"2408FFFE";
        ram_buffer(65113) := X"00A84024";
        ram_buffer(65114) := X"00063027";
        ram_buffer(65115) := X"00851821";
        ram_buffer(65116) := X"00C73824";
        ram_buffer(65117) := X"24490001";
        ram_buffer(65118) := X"00408021";
        ram_buffer(65119) := X"24060002";
        ram_buffer(65120) := X"25050200";
        ram_buffer(65121) := X"00882021";
        ram_buffer(65122) := X"AF8981E4";
        ram_buffer(65123) := X"0C030698";
        ram_buffer(65124) := X"A0670000";
        ram_buffer(65125) := X"1600FF05";
        ram_buffer(65126) := X"00000000";
        ram_buffer(65127) := X"1000000D";
        ram_buffer(65128) := X"00000000";
        ram_buffer(65129) := X"26A400D0";
        ram_buffer(65130) := X"AEA400CC";
        ram_buffer(65131) := X"24060040";
        ram_buffer(65132) := X"0C03068E";
        ram_buffer(65133) := X"00102980";
        ram_buffer(65134) := X"1000FED8";
        ram_buffer(65135) := X"00000000";
        ram_buffer(65136) := X"8EA50040";
        ram_buffer(65137) := X"0C030698";
        ram_buffer(65138) := X"00052980";
        ram_buffer(65139) := X"1000FECB";
        ram_buffer(65140) := X"A2A0003D";
        ram_buffer(65141) := X"8EA400CC";
        ram_buffer(65142) := X"00000000";
        ram_buffer(65143) := X"1080FED7";
        ram_buffer(65144) := X"2410FFFF";
        ram_buffer(65145) := X"1000FEF6";
        ram_buffer(65146) := X"24020001";
        ram_buffer(65147) := X"1000FEC3";
        ram_buffer(65148) := X"00A08021";
        ram_buffer(65149) := X"27C2D288";
        ram_buffer(65150) := X"90450005";
        ram_buffer(65151) := X"90440006";
        ram_buffer(65152) := X"90420007";
        ram_buffer(65153) := X"92060007";
        ram_buffer(65154) := X"92080005";
        ram_buffer(65155) := X"00021027";
        ram_buffer(65156) := X"92070006";
        ram_buffer(65157) := X"00461025";
        ram_buffer(65158) := X"8FA3001C";
        ram_buffer(65159) := X"00052827";
        ram_buffer(65160) := X"00A82825";
        ram_buffer(65161) := X"00042027";
        ram_buffer(65162) := X"A2020007";
        ram_buffer(65163) := X"8FA20018";
        ram_buffer(65164) := X"00872025";
        ram_buffer(65165) := X"A2050005";
        ram_buffer(65166) := X"2465D290";
        ram_buffer(65167) := X"8FA30020";
        ram_buffer(65168) := X"A2040006";
        ram_buffer(65169) := X"2442D690";
        ram_buffer(65170) := X"8CA40000";
        ram_buffer(65171) := X"8C460000";
        ram_buffer(65172) := X"00042027";
        ram_buffer(65173) := X"00862025";
        ram_buffer(65174) := X"AC440000";
        ram_buffer(65175) := X"24420004";
        ram_buffer(65176) := X"1443FFF9";
        ram_buffer(65177) := X"24A50004";
        ram_buffer(65178) := X"8FA20010";
        ram_buffer(65179) := X"02002821";
        ram_buffer(65180) := X"02602021";
        ram_buffer(65181) := X"24060400";
        ram_buffer(65182) := X"AC40D688";
        ram_buffer(65183) := X"0C027F93";
        ram_buffer(65184) := X"A2000004";
        ram_buffer(65185) := X"27C4D288";
        ram_buffer(65186) := X"24060400";
        ram_buffer(65187) := X"0C02801D";
        ram_buffer(65188) := X"240500FF";
        ram_buffer(65189) := X"24060400";
        ram_buffer(65190) := X"240500FF";
        ram_buffer(65191) := X"0C02801D";
        ram_buffer(65192) := X"26640400";
        ram_buffer(65193) := X"1000FF4D";
        ram_buffer(65194) := X"001110C0";
        ram_buffer(65195) := X"27BDFFB8";
        ram_buffer(65196) := X"2402FFFF";
        ram_buffer(65197) := X"AFB7003C";
        ram_buffer(65198) := X"8C970048";
        ram_buffer(65199) := X"AFBE0040";
        ram_buffer(65200) := X"AFB60038";
        ram_buffer(65201) := X"AFB20028";
        ram_buffer(65202) := X"AFB10024";
        ram_buffer(65203) := X"AFB00020";
        ram_buffer(65204) := X"AFBF0044";
        ram_buffer(65205) := X"AFB50034";
        ram_buffer(65206) := X"AFB40030";
        ram_buffer(65207) := X"AFB3002C";
        ram_buffer(65208) := X"0080F021";
        ram_buffer(65209) := X"00C09021";
        ram_buffer(65210) := X"AFA5004C";
        ram_buffer(65211) := X"AFA00018";
        ram_buffer(65212) := X"AFA00014";
        ram_buffer(65213) := X"AFA20010";
        ram_buffer(65214) := X"24D0003C";
        ram_buffer(65215) := X"2411FFFF";
        ram_buffer(65216) := X"24160001";
        ram_buffer(65217) := X"8FD30040";
        ram_buffer(65218) := X"8FD40044";
        ram_buffer(65219) := X"0240A821";
        ram_buffer(65220) := X"8FC20030";
        ram_buffer(65221) := X"00000000";
        ram_buffer(65222) := X"02E2302B";
        ram_buffer(65223) := X"14C00005";
        ram_buffer(65224) := X"03C02021";
        ram_buffer(65225) := X"93C20034";
        ram_buffer(65226) := X"00000000";
        ram_buffer(65227) := X"1040002C";
        ram_buffer(65228) := X"00000000";
        ram_buffer(65229) := X"97C20038";
        ram_buffer(65230) := X"8FC50044";
        ram_buffer(65231) := X"2442FFFC";
        ram_buffer(65232) := X"00A2102B";
        ram_buffer(65233) := X"1440000A";
        ram_buffer(65234) := X"00000000";
        ram_buffer(65235) := X"8FC200CC";
        ram_buffer(65236) := X"00000000";
        ram_buffer(65237) := X"8C420000";
        ram_buffer(65238) := X"00000000";
        ram_buffer(65239) := X"10510020";
        ram_buffer(65240) := X"00402821";
        ram_buffer(65241) := X"0C02FD29";
        ram_buffer(65242) := X"00000000";
        ram_buffer(65243) := X"8FC50044";
        ram_buffer(65244) := X"8FC200CC";
        ram_buffer(65245) := X"24A40001";
        ram_buffer(65246) := X"AFC40044";
        ram_buffer(65247) := X"00452821";
        ram_buffer(65248) := X"90A20004";
        ram_buffer(65249) := X"26B50001";
        ram_buffer(65250) := X"A2A2FFFF";
        ram_buffer(65251) := X"8FC20048";
        ram_buffer(65252) := X"00000000";
        ram_buffer(65253) := X"24570001";
        ram_buffer(65254) := X"1615FFDD";
        ram_buffer(65255) := X"AFD70048";
        ram_buffer(65256) := X"8E440028";
        ram_buffer(65257) := X"00000000";
        ram_buffer(65258) := X"1091000D";
        ram_buffer(65259) := X"00000000";
        ram_buffer(65260) := X"92440036";
        ram_buffer(65261) := X"00000000";
        ram_buffer(65262) := X"10960035";
        ram_buffer(65263) := X"00000000";
        ram_buffer(65264) := X"8FA30010";
        ram_buffer(65265) := X"00000000";
        ram_buffer(65266) := X"1471FFCE";
        ram_buffer(65267) := X"2442FFC5";
        ram_buffer(65268) := X"AFA20018";
        ram_buffer(65269) := X"AFB40014";
        ram_buffer(65270) := X"1000FFCA";
        ram_buffer(65271) := X"AFB30010";
        ram_buffer(65272) := X"93C40037";
        ram_buffer(65273) := X"24020001";
        ram_buffer(65274) := X"10820013";
        ram_buffer(65275) := X"2402FFFF";
        ram_buffer(65276) := X"8FA30010";
        ram_buffer(65277) := X"00000000";
        ram_buffer(65278) := X"1062000F";
        ram_buffer(65279) := X"00000000";
        ram_buffer(65280) := X"8FC20040";
        ram_buffer(65281) := X"00000000";
        ram_buffer(65282) := X"10620003";
        ram_buffer(65283) := X"00602821";
        ram_buffer(65284) := X"0C02FD29";
        ram_buffer(65285) := X"03C02021";
        ram_buffer(65286) := X"8FA20014";
        ram_buffer(65287) := X"00000000";
        ram_buffer(65288) := X"AFC20044";
        ram_buffer(65289) := X"8FA20018";
        ram_buffer(65290) := X"00000000";
        ram_buffer(65291) := X"AFC20048";
        ram_buffer(65292) := X"1000000B";
        ram_buffer(65293) := X"2402FFFF";
        ram_buffer(65294) := X"8FC40040";
        ram_buffer(65295) := X"00000000";
        ram_buffer(65296) := X"12640006";
        ram_buffer(65297) := X"00000000";
        ram_buffer(65298) := X"02602821";
        ram_buffer(65299) := X"03C02021";
        ram_buffer(65300) := X"0C02FD29";
        ram_buffer(65301) := X"AFA20010";
        ram_buffer(65302) := X"8FA20010";
        ram_buffer(65303) := X"AFD40044";
        ram_buffer(65304) := X"8FBF0044";
        ram_buffer(65305) := X"8FBE0040";
        ram_buffer(65306) := X"8FB7003C";
        ram_buffer(65307) := X"8FB60038";
        ram_buffer(65308) := X"8FB50034";
        ram_buffer(65309) := X"8FB40030";
        ram_buffer(65310) := X"8FB3002C";
        ram_buffer(65311) := X"8FB20028";
        ram_buffer(65312) := X"8FB10024";
        ram_buffer(65313) := X"8FB00020";
        ram_buffer(65314) := X"03E00008";
        ram_buffer(65315) := X"27BD0048";
        ram_buffer(65316) := X"8FA5004C";
        ram_buffer(65317) := X"0C02CC2F";
        ram_buffer(65318) := X"02402021";
        ram_buffer(65319) := X"1440FF99";
        ram_buffer(65320) := X"00000000";
        ram_buffer(65321) := X"8FC40040";
        ram_buffer(65322) := X"00000000";
        ram_buffer(65323) := X"1664FFE6";
        ram_buffer(65324) := X"00001021";
        ram_buffer(65325) := X"1000FFEA";
        ram_buffer(65326) := X"AFD40044";
        ram_buffer(65327) := X"3C04100D";
        ram_buffer(65328) := X"27BDFFE8";
        ram_buffer(65329) := X"24060400";
        ram_buffer(65330) := X"24050200";
        ram_buffer(65331) := X"AFBF0014";
        ram_buffer(65332) := X"0C030698";
        ram_buffer(65333) := X"2484D688";
        ram_buffer(65334) := X"8FBF0014";
        ram_buffer(65335) := X"3C04100D";
        ram_buffer(65336) := X"24060400";
        ram_buffer(65337) := X"24050600";
        ram_buffer(65338) := X"2484D288";
        ram_buffer(65339) := X"08030698";
        ram_buffer(65340) := X"27BD0018";
        ram_buffer(65341) := X"27BDFFE8";
        ram_buffer(65342) := X"AFB00010";
        ram_buffer(65343) := X"3C10100D";
        ram_buffer(65344) := X"2604D688";
        ram_buffer(65345) := X"24060400";
        ram_buffer(65346) := X"AFBF0014";
        ram_buffer(65347) := X"0C03068E";
        ram_buffer(65348) := X"24050200";
        ram_buffer(65349) := X"3C04100D";
        ram_buffer(65350) := X"2610D688";
        ram_buffer(65351) := X"24060400";
        ram_buffer(65352) := X"24050600";
        ram_buffer(65353) := X"0C03068E";
        ram_buffer(65354) := X"2484D288";
        ram_buffer(65355) := X"92020005";
        ram_buffer(65356) := X"8FBF0014";
        ram_buffer(65357) := X"24030028";
        ram_buffer(65358) := X"8FB00010";
        ram_buffer(65359) := X"30420001";
        ram_buffer(65360) := X"AF8381E4";
        ram_buffer(65361) := X"03E00008";
        ram_buffer(65362) := X"27BD0018";
        ram_buffer(65363) := X"27BDFFD0";
        ram_buffer(65364) := X"AFB20018";
        ram_buffer(65365) := X"AFBF002C";
        ram_buffer(65366) := X"AFB60028";
        ram_buffer(65367) := X"AFB50024";
        ram_buffer(65368) := X"AFB40020";
        ram_buffer(65369) := X"AFB3001C";
        ram_buffer(65370) := X"AFB10014";
        ram_buffer(65371) := X"AFB00010";
        ram_buffer(65372) := X"18C00031";
        ram_buffer(65373) := X"00009021";
        ram_buffer(65374) := X"00C0A021";
        ram_buffer(65375) := X"0080A821";
        ram_buffer(65376) := X"00A09821";
        ram_buffer(65377) := X"00E08021";
        ram_buffer(65378) := X"2411FFFF";
        ram_buffer(65379) := X"1A600027";
        ram_buffer(65380) := X"00000000";
        ram_buffer(65381) := X"8E020048";
        ram_buffer(65382) := X"02B3B021";
        ram_buffer(65383) := X"8E030030";
        ram_buffer(65384) := X"26B50001";
        ram_buffer(65385) := X"0043102B";
        ram_buffer(65386) := X"14400005";
        ram_buffer(65387) := X"02002021";
        ram_buffer(65388) := X"92020034";
        ram_buffer(65389) := X"00000000";
        ram_buffer(65390) := X"1040001F";
        ram_buffer(65391) := X"00000000";
        ram_buffer(65392) := X"96020038";
        ram_buffer(65393) := X"8E030044";
        ram_buffer(65394) := X"2442FFFC";
        ram_buffer(65395) := X"0062102B";
        ram_buffer(65396) := X"1440000A";
        ram_buffer(65397) := X"00000000";
        ram_buffer(65398) := X"8E0200CC";
        ram_buffer(65399) := X"00000000";
        ram_buffer(65400) := X"8C420000";
        ram_buffer(65401) := X"00000000";
        ram_buffer(65402) := X"10510013";
        ram_buffer(65403) := X"00402821";
        ram_buffer(65404) := X"0C02FD29";
        ram_buffer(65405) := X"00000000";
        ram_buffer(65406) := X"8E030044";
        ram_buffer(65407) := X"8E0200CC";
        ram_buffer(65408) := X"24640001";
        ram_buffer(65409) := X"AE040044";
        ram_buffer(65410) := X"00431821";
        ram_buffer(65411) := X"90620004";
        ram_buffer(65412) := X"00000000";
        ram_buffer(65413) := X"A2A2FFFF";
        ram_buffer(65414) := X"8E020048";
        ram_buffer(65415) := X"00000000";
        ram_buffer(65416) := X"24420001";
        ram_buffer(65417) := X"16B6FFDD";
        ram_buffer(65418) := X"AE020048";
        ram_buffer(65419) := X"26520001";
        ram_buffer(65420) := X"1692FFD6";
        ram_buffer(65421) := X"00000000";
        ram_buffer(65422) := X"8FBF002C";
        ram_buffer(65423) := X"02401021";
        ram_buffer(65424) := X"8FB60028";
        ram_buffer(65425) := X"8FB50024";
        ram_buffer(65426) := X"8FB40020";
        ram_buffer(65427) := X"8FB3001C";
        ram_buffer(65428) := X"8FB20018";
        ram_buffer(65429) := X"8FB10014";
        ram_buffer(65430) := X"8FB00010";
        ram_buffer(65431) := X"03E00008";
        ram_buffer(65432) := X"27BD0030";
        ram_buffer(65433) := X"27BDFFC8";
        ram_buffer(65434) := X"24020001";
        ram_buffer(65435) := X"A0E2003D";
        ram_buffer(65436) := X"AFB2001C";
        ram_buffer(65437) := X"AFB00014";
        ram_buffer(65438) := X"AFBF0034";
        ram_buffer(65439) := X"AFB70030";
        ram_buffer(65440) := X"AFB6002C";
        ram_buffer(65441) := X"AFB50028";
        ram_buffer(65442) := X"AFB40024";
        ram_buffer(65443) := X"AFB30020";
        ram_buffer(65444) := X"AFB10018";
        ram_buffer(65445) := X"00E08021";
        ram_buffer(65446) := X"18C00031";
        ram_buffer(65447) := X"00009021";
        ram_buffer(65448) := X"00C0A021";
        ram_buffer(65449) := X"0080A821";
        ram_buffer(65450) := X"00A09821";
        ram_buffer(65451) := X"2417FFFF";
        ram_buffer(65452) := X"24110001";
        ram_buffer(65453) := X"1E600016";
        ram_buffer(65454) := X"02B3B021";
        ram_buffer(65455) := X"1000003D";
        ram_buffer(65456) := X"26520001";
        ram_buffer(65457) := X"0C02FD29";
        ram_buffer(65458) := X"00000000";
        ram_buffer(65459) := X"8E020040";
        ram_buffer(65460) := X"00000000";
        ram_buffer(65461) := X"10570022";
        ram_buffer(65462) := X"00000000";
        ram_buffer(65463) := X"8E030044";
        ram_buffer(65464) := X"A211003D";
        ram_buffer(65465) := X"24640001";
        ram_buffer(65466) := X"8E0200CC";
        ram_buffer(65467) := X"AE040044";
        ram_buffer(65468) := X"92A4FFFF";
        ram_buffer(65469) := X"00431821";
        ram_buffer(65470) := X"A0640004";
        ram_buffer(65471) := X"8E020048";
        ram_buffer(65472) := X"00000000";
        ram_buffer(65473) := X"24420001";
        ram_buffer(65474) := X"12D50029";
        ram_buffer(65475) := X"AE020048";
        ram_buffer(65476) := X"96020038";
        ram_buffer(65477) := X"8E030044";
        ram_buffer(65478) := X"2442FFFC";
        ram_buffer(65479) := X"0062102B";
        ram_buffer(65480) := X"26B50001";
        ram_buffer(65481) := X"1440FFEF";
        ram_buffer(65482) := X"02002021";
        ram_buffer(65483) := X"8E0200CC";
        ram_buffer(65484) := X"00000000";
        ram_buffer(65485) := X"8C450000";
        ram_buffer(65486) := X"00000000";
        ram_buffer(65487) := X"14B7FFE1";
        ram_buffer(65488) := X"00000000";
        ram_buffer(65489) := X"AC400000";
        ram_buffer(65490) := X"0C02FD29";
        ram_buffer(65491) := X"00002821";
        ram_buffer(65492) := X"8E020040";
        ram_buffer(65493) := X"00000000";
        ram_buffer(65494) := X"1457FFE0";
        ram_buffer(65495) := X"00000000";
        ram_buffer(65496) := X"8E040048";
        ram_buffer(65497) := X"8E020030";
        ram_buffer(65498) := X"24030001";
        ram_buffer(65499) := X"0044102B";
        ram_buffer(65500) := X"A203003D";
        ram_buffer(65501) := X"10400002";
        ram_buffer(65502) := X"A203003C";
        ram_buffer(65503) := X"AE040030";
        ram_buffer(65504) := X"8FBF0034";
        ram_buffer(65505) := X"02401021";
        ram_buffer(65506) := X"8FB70030";
        ram_buffer(65507) := X"8FB6002C";
        ram_buffer(65508) := X"8FB50028";
        ram_buffer(65509) := X"8FB40024";
        ram_buffer(65510) := X"8FB30020";
        ram_buffer(65511) := X"8FB2001C";
        ram_buffer(65512) := X"8FB10018";
        ram_buffer(65513) := X"8FB00014";
        ram_buffer(65514) := X"03E00008";
        ram_buffer(65515) := X"27BD0038";
        ram_buffer(65516) := X"26520001";
        ram_buffer(65517) := X"0254102A";
        ram_buffer(65518) := X"1440FFBE";
        ram_buffer(65519) := X"00000000";
        ram_buffer(65520) := X"1000FFE7";
        ram_buffer(65521) := X"00000000";
        ram_buffer(65522) := X"27BDFFE0";
        ram_buffer(65523) := X"24020001";
        ram_buffer(65524) := X"AFB10014";
        ram_buffer(65525) := X"AFB00010";
        ram_buffer(65526) := X"AFBF001C";
        ram_buffer(65527) := X"AFB20018";
        ram_buffer(65528) := X"00808021";
        ram_buffer(65529) := X"10C20011";
        ram_buffer(65530) := X"00A08821";
        ram_buffer(65531) := X"24020002";
        ram_buffer(65532) := X"10C20030";
        ram_buffer(65533) := X"00000000";
        ram_buffer(65534) := X"10C0000F";
        ram_buffer(65535) := X"00000000";
        ram_buffer(65536) := X"0C030730";
        ram_buffer(65537) := X"00000000";
        ram_buffer(65538) := X"8FBF001C";
        ram_buffer(65539) := X"24030016";
        ram_buffer(65540) := X"AC430000";
        ram_buffer(65541) := X"8FB20018";
        ram_buffer(65542) := X"8FB10014";
        ram_buffer(65543) := X"8FB00010";
        ram_buffer(65544) := X"2402FFFF";
        ram_buffer(65545) := X"03E00008";
        ram_buffer(65546) := X"27BD0020";
        ram_buffer(65547) := X"8C820048";
        ram_buffer(65548) := X"00000000";
        ram_buffer(65549) := X"00A28821";
        ram_buffer(65550) := X"8E050028";
        ram_buffer(65551) := X"AE110048";
        ram_buffer(65552) := X"0C02FD29";
        ram_buffer(65553) := X"02002021";
        ram_buffer(65554) := X"96020038";
        ram_buffer(65555) := X"00000000";
        ram_buffer(65556) := X"2442FFFD";
        ram_buffer(65557) := X"0222102A";
        ram_buffer(65558) := X"1440000E";
        ram_buffer(65559) := X"24120004";
        ram_buffer(65560) := X"8E0200CC";
        ram_buffer(65561) := X"00000000";
        ram_buffer(65562) := X"8C450000";
        ram_buffer(65563) := X"0C02FD29";
        ram_buffer(65564) := X"02002021";
        ram_buffer(65565) := X"96020038";
        ram_buffer(65566) := X"00000000";
        ram_buffer(65567) := X"02421823";
        ram_buffer(65568) := X"02238821";
        ram_buffer(65569) := X"2442FFFD";
        ram_buffer(65570) := X"0222102A";
        ram_buffer(65571) := X"1040FFF4";
        ram_buffer(65572) := X"00000000";
        ram_buffer(65573) := X"8FBF001C";
        ram_buffer(65574) := X"8E020048";
        ram_buffer(65575) := X"AE110044";
        ram_buffer(65576) := X"8FB20018";
        ram_buffer(65577) := X"8FB10014";
        ram_buffer(65578) := X"8FB00010";
        ram_buffer(65579) := X"03E00008";
        ram_buffer(65580) := X"27BD0020";
        ram_buffer(65581) := X"8C820030";
        ram_buffer(65582) := X"1000FFDF";
        ram_buffer(65583) := X"00A28821";
        ram_buffer(65584) := X"27BDFFC0";
        ram_buffer(65585) := X"AFB20020";
        ram_buffer(65586) := X"AFA50044";
        ram_buffer(65587) := X"00C09021";
        ram_buffer(65588) := X"00002821";
        ram_buffer(65589) := X"24060110";
        ram_buffer(65590) := X"AFBF003C";
        ram_buffer(65591) := X"AFBE0038";
        ram_buffer(65592) := X"AFB60030";
        ram_buffer(65593) := X"AFB5002C";
        ram_buffer(65594) := X"0080B021";
        ram_buffer(65595) := X"AFB40028";
        ram_buffer(65596) := X"AFB30024";
        ram_buffer(65597) := X"AFB1001C";
        ram_buffer(65598) := X"AFB00018";
        ram_buffer(65599) := X"00E08821";
        ram_buffer(65600) := X"0C02801D";
        ram_buffer(65601) := X"AFB70034";
        ram_buffer(65602) := X"3C02100D";
        ram_buffer(65603) := X"2442DA88";
        ram_buffer(65604) := X"00402821";
        ram_buffer(65605) := X"02C02021";
        ram_buffer(65606) := X"2406003C";
        ram_buffer(65607) := X"0C027F93";
        ram_buffer(65608) := X"AFA20010";
        ram_buffer(65609) := X"8EC50028";
        ram_buffer(65610) := X"0C02FD29";
        ram_buffer(65611) := X"02C02021";
        ram_buffer(65612) := X"8EC20040";
        ram_buffer(65613) := X"8FB00044";
        ram_buffer(65614) := X"AEC20028";
        ram_buffer(65615) := X"AEC00048";
        ram_buffer(65616) := X"82020000";
        ram_buffer(65617) := X"3C14100D";
        ram_buffer(65618) := X"241E002F";
        ram_buffer(65619) := X"24150027";
        ram_buffer(65620) := X"2694B3C4";
        ram_buffer(65621) := X"105E0042";
        ram_buffer(65622) := X"24130001";
        ram_buffer(65623) := X"02002021";
        ram_buffer(65624) := X"02202821";
        ram_buffer(65625) := X"10000006";
        ram_buffer(65626) := X"00001821";
        ram_buffer(65627) := X"105E0008";
        ram_buffer(65628) := X"24840001";
        ram_buffer(65629) := X"A0A20000";
        ram_buffer(65630) := X"1075003B";
        ram_buffer(65631) := X"24A50001";
        ram_buffer(65632) := X"80820000";
        ram_buffer(65633) := X"0060B821";
        ram_buffer(65634) := X"1440FFF8";
        ram_buffer(65635) := X"24630001";
        ram_buffer(65636) := X"02371021";
        ram_buffer(65637) := X"A0400000";
        ram_buffer(65638) := X"02403021";
        ram_buffer(65639) := X"02202821";
        ram_buffer(65640) := X"0C02FEAB";
        ram_buffer(65641) := X"02C02021";
        ram_buffer(65642) := X"14400039";
        ram_buffer(65643) := X"00000000";
        ram_buffer(65644) := X"02178021";
        ram_buffer(65645) := X"82020000";
        ram_buffer(65646) := X"00000000";
        ram_buffer(65647) := X"1040004F";
        ram_buffer(65648) := X"02202821";
        ram_buffer(65649) := X"8FA60044";
        ram_buffer(65650) := X"0C028116";
        ram_buffer(65651) := X"02802021";
        ram_buffer(65652) := X"24060110";
        ram_buffer(65653) := X"00002821";
        ram_buffer(65654) := X"0C02801D";
        ram_buffer(65655) := X"02C02021";
        ram_buffer(65656) := X"12400040";
        ram_buffer(65657) := X"2406003C";
        ram_buffer(65658) := X"92420036";
        ram_buffer(65659) := X"00000000";
        ram_buffer(65660) := X"10530035";
        ram_buffer(65661) := X"24170001";
        ram_buffer(65662) := X"02C02021";
        ram_buffer(65663) := X"2406003C";
        ram_buffer(65664) := X"00002821";
        ram_buffer(65665) := X"A2D3003C";
        ram_buffer(65666) := X"0C02801D";
        ram_buffer(65667) := X"A2D7003D";
        ram_buffer(65668) := X"02202821";
        ram_buffer(65669) := X"24060027";
        ram_buffer(65670) := X"0C02CCBF";
        ram_buffer(65671) := X"02C02021";
        ram_buffer(65672) := X"A2D70036";
        ram_buffer(65673) := X"96420038";
        ram_buffer(65674) := X"AEC00028";
        ram_buffer(65675) := X"A6C20038";
        ram_buffer(65676) := X"92420037";
        ram_buffer(65677) := X"00002821";
        ram_buffer(65678) := X"A2C20037";
        ram_buffer(65679) := X"0C02FD29";
        ram_buffer(65680) := X"02C02021";
        ram_buffer(65681) := X"8EC20040";
        ram_buffer(65682) := X"AEC00048";
        ram_buffer(65683) := X"AEC20028";
        ram_buffer(65684) := X"82020000";
        ram_buffer(65685) := X"00000000";
        ram_buffer(65686) := X"145EFFC0";
        ram_buffer(65687) := X"00000000";
        ram_buffer(65688) := X"1000FFBE";
        ram_buffer(65689) := X"26100001";
        ram_buffer(65690) := X"24170027";
        ram_buffer(65691) := X"02371021";
        ram_buffer(65692) := X"A0400000";
        ram_buffer(65693) := X"02403021";
        ram_buffer(65694) := X"02202821";
        ram_buffer(65695) := X"0C02FEAB";
        ram_buffer(65696) := X"02C02021";
        ram_buffer(65697) := X"1040FFCB";
        ram_buffer(65698) := X"02178021";
        ram_buffer(65699) := X"02178023";
        ram_buffer(65700) := X"AFA20010";
        ram_buffer(65701) := X"92C20037";
        ram_buffer(65702) := X"2405002F";
        ram_buffer(65703) := X"A2420037";
        ram_buffer(65704) := X"96C20038";
        ram_buffer(65705) := X"02002021";
        ram_buffer(65706) := X"A6420038";
        ram_buffer(65707) := X"0C03087D";
        ram_buffer(65708) := X"A2400036";
        ram_buffer(65709) := X"8FA30010";
        ram_buffer(65710) := X"1440001D";
        ram_buffer(65711) := X"00000000";
        ram_buffer(65712) := X"1000000F";
        ram_buffer(65713) := X"00601021";
        ram_buffer(65714) := X"02402821";
        ram_buffer(65715) := X"2406003C";
        ram_buffer(65716) := X"0C027F93";
        ram_buffer(65717) := X"02C02021";
        ram_buffer(65718) := X"8EC50028";
        ram_buffer(65719) := X"1000FFD7";
        ram_buffer(65720) := X"00000000";
        ram_buffer(65721) := X"8FA50010";
        ram_buffer(65722) := X"0C027F93";
        ram_buffer(65723) := X"02C02021";
        ram_buffer(65724) := X"8EC50028";
        ram_buffer(65725) := X"1000FFD1";
        ram_buffer(65726) := X"00000000";
        ram_buffer(65727) := X"00001021";
        ram_buffer(65728) := X"8FBF003C";
        ram_buffer(65729) := X"8FBE0038";
        ram_buffer(65730) := X"8FB70034";
        ram_buffer(65731) := X"8FB60030";
        ram_buffer(65732) := X"8FB5002C";
        ram_buffer(65733) := X"8FB40028";
        ram_buffer(65734) := X"8FB30024";
        ram_buffer(65735) := X"8FB20020";
        ram_buffer(65736) := X"8FB1001C";
        ram_buffer(65737) := X"8FB00018";
        ram_buffer(65738) := X"03E00008";
        ram_buffer(65739) := X"27BD0040";
        ram_buffer(65740) := X"1000FFF3";
        ram_buffer(65741) := X"2402FFFE";
        ram_buffer(65742) := X"27BDFED8";
        ram_buffer(65743) := X"27A40010";
        ram_buffer(65744) := X"24060110";
        ram_buffer(65745) := X"00002821";
        ram_buffer(65746) := X"AFBF0124";
        ram_buffer(65747) := X"0C02801D";
        ram_buffer(65748) := X"AFB00120";
        ram_buffer(65749) := X"3C10100D";
        ram_buffer(65750) := X"24020040";
        ram_buffer(65751) := X"2604D688";
        ram_buffer(65752) := X"24060400";
        ram_buffer(65753) := X"24050200";
        ram_buffer(65754) := X"A7A20048";
        ram_buffer(65755) := X"24020001";
        ram_buffer(65756) := X"0C03068E";
        ram_buffer(65757) := X"A3A20047";
        ram_buffer(65758) := X"3C04100D";
        ram_buffer(65759) := X"24060400";
        ram_buffer(65760) := X"24050600";
        ram_buffer(65761) := X"2484D288";
        ram_buffer(65762) := X"0C03068E";
        ram_buffer(65763) := X"2610D688";
        ram_buffer(65764) := X"92020005";
        ram_buffer(65765) := X"24030028";
        ram_buffer(65766) := X"30420001";
        ram_buffer(65767) := X"14400036";
        ram_buffer(65768) := X"AF8381E4";
        ram_buffer(65769) := X"8FA400DC";
        ram_buffer(65770) := X"00000000";
        ram_buffer(65771) := X"10800005";
        ram_buffer(65772) := X"00000000";
        ram_buffer(65773) := X"93A2004D";
        ram_buffer(65774) := X"00000000";
        ram_buffer(65775) := X"14400014";
        ram_buffer(65776) := X"00000000";
        ram_buffer(65777) := X"93A20047";
        ram_buffer(65778) := X"24030028";
        ram_buffer(65779) := X"AFA30050";
        ram_buffer(65780) := X"14400018";
        ram_buffer(65781) := X"AFA00054";
        ram_buffer(65782) := X"3C04100D";
        ram_buffer(65783) := X"2482DA88";
        ram_buffer(65784) := X"AC430028";
        ram_buffer(65785) := X"97A30048";
        ram_buffer(65786) := X"24052F00";
        ram_buffer(65787) := X"A4430038";
        ram_buffer(65788) := X"24030001";
        ram_buffer(65789) := X"A485DA88";
        ram_buffer(65790) := X"A0400037";
        ram_buffer(65791) := X"A0430034";
        ram_buffer(65792) := X"8FBF0124";
        ram_buffer(65793) := X"8FB00120";
        ram_buffer(65794) := X"03E00008";
        ram_buffer(65795) := X"27BD0128";
        ram_buffer(65796) := X"93A20047";
        ram_buffer(65797) := X"00000000";
        ram_buffer(65798) := X"14400011";
        ram_buffer(65799) := X"24060040";
        ram_buffer(65800) := X"A3A0004D";
        ram_buffer(65801) := X"24030028";
        ram_buffer(65802) := X"AFA30050";
        ram_buffer(65803) := X"1040FFEA";
        ram_buffer(65804) := X"AFA00054";
        ram_buffer(65805) := X"27A200E0";
        ram_buffer(65806) := X"24060040";
        ram_buffer(65807) := X"24050A00";
        ram_buffer(65808) := X"00402021";
        ram_buffer(65809) := X"0C03068E";
        ram_buffer(65810) := X"AFA200DC";
        ram_buffer(65811) := X"93A60047";
        ram_buffer(65812) := X"8FA50050";
        ram_buffer(65813) := X"8FA400DC";
        ram_buffer(65814) := X"1000000E";
        ram_buffer(65815) := X"3C03100D";
        ram_buffer(65816) := X"8FA50050";
        ram_buffer(65817) := X"0C030698";
        ram_buffer(65818) := X"00052980";
        ram_buffer(65819) := X"93A20047";
        ram_buffer(65820) := X"1000FFEC";
        ram_buffer(65821) := X"A3A0004D";
        ram_buffer(65822) := X"00002821";
        ram_buffer(65823) := X"0C02FD29";
        ram_buffer(65824) := X"27A40010";
        ram_buffer(65825) := X"93A60047";
        ram_buffer(65826) := X"8FA50050";
        ram_buffer(65827) := X"8FA400DC";
        ram_buffer(65828) := X"3C03100D";
        ram_buffer(65829) := X"24072F00";
        ram_buffer(65830) := X"2462DA88";
        ram_buffer(65831) := X"A467DA88";
        ram_buffer(65832) := X"97A30048";
        ram_buffer(65833) := X"A0460037";
        ram_buffer(65834) := X"A4430038";
        ram_buffer(65835) := X"24030001";
        ram_buffer(65836) := X"AC450028";
        ram_buffer(65837) := X"1080FFD2";
        ram_buffer(65838) := X"A0430034";
        ram_buffer(65839) := X"93A2004D";
        ram_buffer(65840) := X"00000000";
        ram_buffer(65841) := X"1040FFCE";
        ram_buffer(65842) := X"00000000";
        ram_buffer(65843) := X"10C0FFCC";
        ram_buffer(65844) := X"24060040";
        ram_buffer(65845) := X"0C030698";
        ram_buffer(65846) := X"00052980";
        ram_buffer(65847) := X"8FBF0124";
        ram_buffer(65848) := X"8FB00120";
        ram_buffer(65849) := X"03E00008";
        ram_buffer(65850) := X"27BD0128";
        ram_buffer(65851) := X"27BDFE60";
        ram_buffer(65852) := X"AFB20190";
        ram_buffer(65853) := X"AFBF019C";
        ram_buffer(65854) := X"AFB40198";
        ram_buffer(65855) := X"AFB30194";
        ram_buffer(65856) := X"AFB1018C";
        ram_buffer(65857) := X"AFB00188";
        ram_buffer(65858) := X"9082003C";
        ram_buffer(65859) := X"00000000";
        ram_buffer(65860) := X"1440000A";
        ram_buffer(65861) := X"00809021";
        ram_buffer(65862) := X"8FBF019C";
        ram_buffer(65863) := X"8FB40198";
        ram_buffer(65864) := X"8FB30194";
        ram_buffer(65865) := X"8FB1018C";
        ram_buffer(65866) := X"8FB00188";
        ram_buffer(65867) := X"02402021";
        ram_buffer(65868) := X"8FB20190";
        ram_buffer(65869) := X"08027A4D";
        ram_buffer(65870) := X"27BD01A0";
        ram_buffer(65871) := X"8C8400CC";
        ram_buffer(65872) := X"00000000";
        ram_buffer(65873) := X"10800005";
        ram_buffer(65874) := X"27B0015C";
        ram_buffer(65875) := X"9242003D";
        ram_buffer(65876) := X"00000000";
        ram_buffer(65877) := X"1440004D";
        ram_buffer(65878) := X"00000000";
        ram_buffer(65879) := X"27A40010";
        ram_buffer(65880) := X"02003821";
        ram_buffer(65881) := X"27A60120";
        ram_buffer(65882) := X"0C030030";
        ram_buffer(65883) := X"2645004C";
        ram_buffer(65884) := X"92430037";
        ram_buffer(65885) := X"24040001";
        ram_buffer(65886) := X"10640053";
        ram_buffer(65887) := X"00000000";
        ram_buffer(65888) := X"24020001";
        ram_buffer(65889) := X"02409821";
        ram_buffer(65890) := X"A3A2004D";
        ram_buffer(65891) := X"2650003C";
        ram_buffer(65892) := X"2414FFFF";
        ram_buffer(65893) := X"10000014";
        ram_buffer(65894) := X"24110001";
        ram_buffer(65895) := X"0C02FD29";
        ram_buffer(65896) := X"00000000";
        ram_buffer(65897) := X"8FA20050";
        ram_buffer(65898) := X"00000000";
        ram_buffer(65899) := X"10540022";
        ram_buffer(65900) := X"00000000";
        ram_buffer(65901) := X"8FA30054";
        ram_buffer(65902) := X"A3B1004D";
        ram_buffer(65903) := X"8FA200DC";
        ram_buffer(65904) := X"9264FFFF";
        ram_buffer(65905) := X"24650001";
        ram_buffer(65906) := X"00431821";
        ram_buffer(65907) := X"AFA50054";
        ram_buffer(65908) := X"A0640004";
        ram_buffer(65909) := X"8FA20058";
        ram_buffer(65910) := X"00000000";
        ram_buffer(65911) := X"24420001";
        ram_buffer(65912) := X"12700016";
        ram_buffer(65913) := X"AFA20058";
        ram_buffer(65914) := X"97A20048";
        ram_buffer(65915) := X"8FA30054";
        ram_buffer(65916) := X"2442FFFC";
        ram_buffer(65917) := X"0062102B";
        ram_buffer(65918) := X"26730001";
        ram_buffer(65919) := X"1440FFEF";
        ram_buffer(65920) := X"27A40010";
        ram_buffer(65921) := X"8FA200DC";
        ram_buffer(65922) := X"00000000";
        ram_buffer(65923) := X"8C450000";
        ram_buffer(65924) := X"00000000";
        ram_buffer(65925) := X"14B4FFE1";
        ram_buffer(65926) := X"00000000";
        ram_buffer(65927) := X"AC400000";
        ram_buffer(65928) := X"0C02FD29";
        ram_buffer(65929) := X"00002821";
        ram_buffer(65930) := X"8FA20050";
        ram_buffer(65931) := X"00000000";
        ram_buffer(65932) := X"1454FFE0";
        ram_buffer(65933) := X"00000000";
        ram_buffer(65934) := X"8FA20058";
        ram_buffer(65935) := X"8FA30040";
        ram_buffer(65936) := X"24040001";
        ram_buffer(65937) := X"0062182B";
        ram_buffer(65938) := X"A3A4004D";
        ram_buffer(65939) := X"10600002";
        ram_buffer(65940) := X"A3A4004C";
        ram_buffer(65941) := X"AFA20040";
        ram_buffer(65942) := X"8FA400DC";
        ram_buffer(65943) := X"00000000";
        ram_buffer(65944) := X"1080FFAD";
        ram_buffer(65945) := X"00000000";
        ram_buffer(65946) := X"93A20047";
        ram_buffer(65947) := X"00000000";
        ram_buffer(65948) := X"1040FFA9";
        ram_buffer(65949) := X"24060040";
        ram_buffer(65950) := X"8FA50050";
        ram_buffer(65951) := X"0C030698";
        ram_buffer(65952) := X"00052980";
        ram_buffer(65953) := X"1000FFA4";
        ram_buffer(65954) := X"00000000";
        ram_buffer(65955) := X"92420037";
        ram_buffer(65956) := X"00000000";
        ram_buffer(65957) := X"1440004A";
        ram_buffer(65958) := X"24060040";
        ram_buffer(65959) := X"A240003D";
        ram_buffer(65960) := X"27B0015C";
        ram_buffer(65961) := X"27A40010";
        ram_buffer(65962) := X"02003821";
        ram_buffer(65963) := X"27A60120";
        ram_buffer(65964) := X"0C030030";
        ram_buffer(65965) := X"2645004C";
        ram_buffer(65966) := X"92430037";
        ram_buffer(65967) := X"24040001";
        ram_buffer(65968) := X"1464FFAF";
        ram_buffer(65969) := X"00000000";
        ram_buffer(65970) := X"1440FFAE";
        ram_buffer(65971) := X"24020001";
        ram_buffer(65972) := X"A3A00156";
        ram_buffer(65973) := X"A3A3004D";
        ram_buffer(65974) := X"27B30120";
        ram_buffer(65975) := X"2414FFFF";
        ram_buffer(65976) := X"10000014";
        ram_buffer(65977) := X"24110001";
        ram_buffer(65978) := X"0C02FD29";
        ram_buffer(65979) := X"00000000";
        ram_buffer(65980) := X"8FA20050";
        ram_buffer(65981) := X"00000000";
        ram_buffer(65982) := X"10540022";
        ram_buffer(65983) := X"00000000";
        ram_buffer(65984) := X"8FA30054";
        ram_buffer(65985) := X"A3B1004D";
        ram_buffer(65986) := X"8FA200DC";
        ram_buffer(65987) := X"9264FFFF";
        ram_buffer(65988) := X"24650001";
        ram_buffer(65989) := X"00431821";
        ram_buffer(65990) := X"AFA50054";
        ram_buffer(65991) := X"A0640004";
        ram_buffer(65992) := X"8FA20058";
        ram_buffer(65993) := X"00000000";
        ram_buffer(65994) := X"24420001";
        ram_buffer(65995) := X"12700016";
        ram_buffer(65996) := X"AFA20058";
        ram_buffer(65997) := X"97A20048";
        ram_buffer(65998) := X"8FA30054";
        ram_buffer(65999) := X"2442FFFC";
        ram_buffer(66000) := X"0062102B";
        ram_buffer(66001) := X"26730001";
        ram_buffer(66002) := X"1440FFEF";
        ram_buffer(66003) := X"27A40010";
        ram_buffer(66004) := X"8FA200DC";
        ram_buffer(66005) := X"00000000";
        ram_buffer(66006) := X"8C450000";
        ram_buffer(66007) := X"00000000";
        ram_buffer(66008) := X"14B4FFE1";
        ram_buffer(66009) := X"00000000";
        ram_buffer(66010) := X"AC400000";
        ram_buffer(66011) := X"0C02FD29";
        ram_buffer(66012) := X"00002821";
        ram_buffer(66013) := X"8FA20050";
        ram_buffer(66014) := X"00000000";
        ram_buffer(66015) := X"1454FFE0";
        ram_buffer(66016) := X"00000000";
        ram_buffer(66017) := X"8FA20058";
        ram_buffer(66018) := X"8FA30040";
        ram_buffer(66019) := X"24040001";
        ram_buffer(66020) := X"0062182B";
        ram_buffer(66021) := X"A3A4004D";
        ram_buffer(66022) := X"10600002";
        ram_buffer(66023) := X"A3A4004C";
        ram_buffer(66024) := X"AFA20040";
        ram_buffer(66025) := X"3C05100D";
        ram_buffer(66026) := X"27A60120";
        ram_buffer(66027) := X"24A5B3E4";
        ram_buffer(66028) := X"0C02FEAB";
        ram_buffer(66029) := X"27A40010";
        ram_buffer(66030) := X"1000FF72";
        ram_buffer(66031) := X"24020001";
        ram_buffer(66032) := X"8E450040";
        ram_buffer(66033) := X"0C030698";
        ram_buffer(66034) := X"00052980";
        ram_buffer(66035) := X"1000FFB4";
        ram_buffer(66036) := X"A240003D";
        ram_buffer(66037) := X"27BDFD48";
        ram_buffer(66038) := X"AFB00298";
        ram_buffer(66039) := X"27B0026C";
        ram_buffer(66040) := X"00802821";
        ram_buffer(66041) := X"02003821";
        ram_buffer(66042) := X"27A60230";
        ram_buffer(66043) := X"27A40120";
        ram_buffer(66044) := X"AFB202A0";
        ram_buffer(66045) := X"AFBF02B4";
        ram_buffer(66046) := X"AFB602B0";
        ram_buffer(66047) := X"AFB502AC";
        ram_buffer(66048) := X"AFB402A8";
        ram_buffer(66049) := X"AFB302A4";
        ram_buffer(66050) := X"0C030030";
        ram_buffer(66051) := X"AFB1029C";
        ram_buffer(66052) := X"1040000C";
        ram_buffer(66053) := X"00409021";
        ram_buffer(66054) := X"8FBF02B4";
        ram_buffer(66055) := X"02401021";
        ram_buffer(66056) := X"8FB602B0";
        ram_buffer(66057) := X"8FB502AC";
        ram_buffer(66058) := X"8FB402A8";
        ram_buffer(66059) := X"8FB302A4";
        ram_buffer(66060) := X"8FB202A0";
        ram_buffer(66061) := X"8FB1029C";
        ram_buffer(66062) := X"8FB00298";
        ram_buffer(66063) := X"03E00008";
        ram_buffer(66064) := X"27BD02B8";
        ram_buffer(66065) := X"24060110";
        ram_buffer(66066) := X"00002821";
        ram_buffer(66067) := X"0C02801D";
        ram_buffer(66068) := X"27A40010";
        ram_buffer(66069) := X"93A20266";
        ram_buffer(66070) := X"24110001";
        ram_buffer(66071) := X"1051009A";
        ram_buffer(66072) := X"27A40010";
        ram_buffer(66073) := X"2406003C";
        ram_buffer(66074) := X"00002821";
        ram_buffer(66075) := X"A3B1004C";
        ram_buffer(66076) := X"0C02801D";
        ram_buffer(66077) := X"A3B1004D";
        ram_buffer(66078) := X"00002821";
        ram_buffer(66079) := X"24060027";
        ram_buffer(66080) := X"0C02CCBF";
        ram_buffer(66081) := X"27A40010";
        ram_buffer(66082) := X"97A20268";
        ram_buffer(66083) := X"A3B10046";
        ram_buffer(66084) := X"A7A20048";
        ram_buffer(66085) := X"93A20267";
        ram_buffer(66086) := X"00002821";
        ram_buffer(66087) := X"A3A20047";
        ram_buffer(66088) := X"0C02FD29";
        ram_buffer(66089) := X"27A40010";
        ram_buffer(66090) := X"8FA200DC";
        ram_buffer(66091) := X"8FB60050";
        ram_buffer(66092) := X"8C450000";
        ram_buffer(66093) := X"2402FFFF";
        ram_buffer(66094) := X"AFB60038";
        ram_buffer(66095) := X"10A20027";
        ram_buffer(66096) := X"AFA00058";
        ram_buffer(66097) := X"3C11100D";
        ram_buffer(66098) := X"2631D288";
        ram_buffer(66099) := X"24150001";
        ram_buffer(66100) := X"2414FFFE";
        ram_buffer(66101) := X"10000009";
        ram_buffer(66102) := X"2413FFFF";
        ram_buffer(66103) := X"0C027A4D";
        ram_buffer(66104) := X"00000000";
        ram_buffer(66105) := X"8FA200DC";
        ram_buffer(66106) := X"8FB60050";
        ram_buffer(66107) := X"8C450000";
        ram_buffer(66108) := X"00000000";
        ram_buffer(66109) := X"10B30019";
        ram_buffer(66110) := X"00000000";
        ram_buffer(66111) := X"0C02FD29";
        ram_buffer(66112) := X"27A40010";
        ram_buffer(66113) := X"001618C3";
        ram_buffer(66114) := X"32C20007";
        ram_buffer(66115) := X"93A80047";
        ram_buffer(66116) := X"00713821";
        ram_buffer(66117) := X"00551004";
        ram_buffer(66118) := X"00741824";
        ram_buffer(66119) := X"00021027";
        ram_buffer(66120) := X"02C02021";
        ram_buffer(66121) := X"24060002";
        ram_buffer(66122) := X"1100FFEC";
        ram_buffer(66123) := X"24650600";
        ram_buffer(66124) := X"90E80000";
        ram_buffer(66125) := X"02232021";
        ram_buffer(66126) := X"00481024";
        ram_buffer(66127) := X"0C030698";
        ram_buffer(66128) := X"A0E20000";
        ram_buffer(66129) := X"8FA200DC";
        ram_buffer(66130) := X"8FB60050";
        ram_buffer(66131) := X"8C450000";
        ram_buffer(66132) := X"00000000";
        ram_buffer(66133) := X"14B3FFE9";
        ram_buffer(66134) := X"00000000";
        ram_buffer(66135) := X"93A20047";
        ram_buffer(66136) := X"00000000";
        ram_buffer(66137) := X"14400046";
        ram_buffer(66138) := X"001618C3";
        ram_buffer(66139) := X"0C027A4D";
        ram_buffer(66140) := X"02C02021";
        ram_buffer(66141) := X"24020001";
        ram_buffer(66142) := X"A3A00266";
        ram_buffer(66143) := X"A3A2015D";
        ram_buffer(66144) := X"27B30230";
        ram_buffer(66145) := X"2414FFFF";
        ram_buffer(66146) := X"10000014";
        ram_buffer(66147) := X"24110001";
        ram_buffer(66148) := X"0C02FD29";
        ram_buffer(66149) := X"00000000";
        ram_buffer(66150) := X"8FA20160";
        ram_buffer(66151) := X"00000000";
        ram_buffer(66152) := X"10540022";
        ram_buffer(66153) := X"00000000";
        ram_buffer(66154) := X"8FA30164";
        ram_buffer(66155) := X"A3B1015D";
        ram_buffer(66156) := X"8FA201EC";
        ram_buffer(66157) := X"9264FFFF";
        ram_buffer(66158) := X"24650001";
        ram_buffer(66159) := X"00431821";
        ram_buffer(66160) := X"AFA50164";
        ram_buffer(66161) := X"A0640004";
        ram_buffer(66162) := X"8FA20168";
        ram_buffer(66163) := X"00000000";
        ram_buffer(66164) := X"24420001";
        ram_buffer(66165) := X"12700016";
        ram_buffer(66166) := X"AFA20168";
        ram_buffer(66167) := X"97A20158";
        ram_buffer(66168) := X"8FA30164";
        ram_buffer(66169) := X"2442FFFC";
        ram_buffer(66170) := X"0062102B";
        ram_buffer(66171) := X"26730001";
        ram_buffer(66172) := X"1440FFEF";
        ram_buffer(66173) := X"27A40120";
        ram_buffer(66174) := X"8FA201EC";
        ram_buffer(66175) := X"00000000";
        ram_buffer(66176) := X"8C450000";
        ram_buffer(66177) := X"00000000";
        ram_buffer(66178) := X"14B4FFE1";
        ram_buffer(66179) := X"00000000";
        ram_buffer(66180) := X"AC400000";
        ram_buffer(66181) := X"0C02FD29";
        ram_buffer(66182) := X"00002821";
        ram_buffer(66183) := X"8FA20160";
        ram_buffer(66184) := X"00000000";
        ram_buffer(66185) := X"1454FFE0";
        ram_buffer(66186) := X"00000000";
        ram_buffer(66187) := X"8FA20168";
        ram_buffer(66188) := X"8FA30150";
        ram_buffer(66189) := X"24040001";
        ram_buffer(66190) := X"0062182B";
        ram_buffer(66191) := X"A3A4015D";
        ram_buffer(66192) := X"10600002";
        ram_buffer(66193) := X"A3A4015C";
        ram_buffer(66194) := X"AFA20150";
        ram_buffer(66195) := X"8FA401EC";
        ram_buffer(66196) := X"00000000";
        ram_buffer(66197) := X"1080FF70";
        ram_buffer(66198) := X"00000000";
        ram_buffer(66199) := X"93A20157";
        ram_buffer(66200) := X"00000000";
        ram_buffer(66201) := X"1040FF6C";
        ram_buffer(66202) := X"24060040";
        ram_buffer(66203) := X"8FA50160";
        ram_buffer(66204) := X"0C030698";
        ram_buffer(66205) := X"00052980";
        ram_buffer(66206) := X"1000FF67";
        ram_buffer(66207) := X"00000000";
        ram_buffer(66208) := X"3C04100D";
        ram_buffer(66209) := X"2484D288";
        ram_buffer(66210) := X"00643821";
        ram_buffer(66211) := X"24020001";
        ram_buffer(66212) := X"32D60007";
        ram_buffer(66213) := X"90E50000";
        ram_buffer(66214) := X"02C2B004";
        ram_buffer(66215) := X"2402FFFE";
        ram_buffer(66216) := X"00621824";
        ram_buffer(66217) := X"00161027";
        ram_buffer(66218) := X"00451024";
        ram_buffer(66219) := X"24060002";
        ram_buffer(66220) := X"24650600";
        ram_buffer(66221) := X"00832021";
        ram_buffer(66222) := X"0C030698";
        ram_buffer(66223) := X"A0E20000";
        ram_buffer(66224) := X"1000FFAD";
        ram_buffer(66225) := X"24020001";
        ram_buffer(66226) := X"27A50230";
        ram_buffer(66227) := X"2406003C";
        ram_buffer(66228) := X"0C027F93";
        ram_buffer(66229) := X"27A40010";
        ram_buffer(66230) := X"8FA50038";
        ram_buffer(66231) := X"1000FF70";
        ram_buffer(66232) := X"00000000";
        ram_buffer(66233) := X"27BDFE58";
        ram_buffer(66234) := X"AFB10190";
        ram_buffer(66235) := X"3C11100D";
        ram_buffer(66236) := X"2631DA88";
        ram_buffer(66237) := X"8E220028";
        ram_buffer(66238) := X"AFB30198";
        ram_buffer(66239) := X"AFB20194";
        ram_buffer(66240) := X"AFBF01A4";
        ram_buffer(66241) := X"AFB501A0";
        ram_buffer(66242) := X"AFB4019C";
        ram_buffer(66243) := X"AFB0018C";
        ram_buffer(66244) := X"00809021";
        ram_buffer(66245) := X"1040006A";
        ram_buffer(66246) := X"00A09821";
        ram_buffer(66247) := X"24050001";
        ram_buffer(66248) := X"0C03071E";
        ram_buffer(66249) := X"24040110";
        ram_buffer(66250) := X"1040009C";
        ram_buffer(66251) := X"00408021";
        ram_buffer(66252) := X"82420000";
        ram_buffer(66253) := X"00000000";
        ram_buffer(66254) := X"10400023";
        ram_buffer(66255) := X"3C05100D";
        ram_buffer(66256) := X"24A5B3F0";
        ram_buffer(66257) := X"0C02CC2F";
        ram_buffer(66258) := X"02402021";
        ram_buffer(66259) := X"1040001E";
        ram_buffer(66260) := X"24020077";
        ram_buffer(66261) := X"82630000";
        ram_buffer(66262) := X"27B1015C";
        ram_buffer(66263) := X"27B40120";
        ram_buffer(66264) := X"1062005B";
        ram_buffer(66265) := X"27B50010";
        ram_buffer(66266) := X"02203821";
        ram_buffer(66267) := X"02803021";
        ram_buffer(66268) := X"02402821";
        ram_buffer(66269) := X"0C030030";
        ram_buffer(66270) := X"02A02021";
        ram_buffer(66271) := X"2403FFFE";
        ram_buffer(66272) := X"1043007E";
        ram_buffer(66273) := X"00000000";
        ram_buffer(66274) := X"14400023";
        ram_buffer(66275) := X"24020072";
        ram_buffer(66276) := X"93B50156";
        ram_buffer(66277) := X"24060110";
        ram_buffer(66278) := X"00002821";
        ram_buffer(66279) := X"0C02801D";
        ram_buffer(66280) := X"02002021";
        ram_buffer(66281) := X"24020001";
        ram_buffer(66282) := X"16A20023";
        ram_buffer(66283) := X"02802821";
        ram_buffer(66284) := X"2406003C";
        ram_buffer(66285) := X"0C027F93";
        ram_buffer(66286) := X"02002021";
        ram_buffer(66287) := X"8E050028";
        ram_buffer(66288) := X"1000002F";
        ram_buffer(66289) := X"00000000";
        ram_buffer(66290) := X"02202821";
        ram_buffer(66291) := X"02002021";
        ram_buffer(66292) := X"0C027F93";
        ram_buffer(66293) := X"2406003C";
        ram_buffer(66294) := X"8E050028";
        ram_buffer(66295) := X"0C02FD29";
        ram_buffer(66296) := X"02002021";
        ram_buffer(66297) := X"8E020040";
        ram_buffer(66298) := X"AE000048";
        ram_buffer(66299) := X"AE020028";
        ram_buffer(66300) := X"02001021";
        ram_buffer(66301) := X"8FBF01A4";
        ram_buffer(66302) := X"8FB501A0";
        ram_buffer(66303) := X"8FB4019C";
        ram_buffer(66304) := X"8FB30198";
        ram_buffer(66305) := X"8FB20194";
        ram_buffer(66306) := X"8FB10190";
        ram_buffer(66307) := X"8FB0018C";
        ram_buffer(66308) := X"03E00008";
        ram_buffer(66309) := X"27BD01A8";
        ram_buffer(66310) := X"82630000";
        ram_buffer(66311) := X"00000000";
        ram_buffer(66312) := X"10620056";
        ram_buffer(66313) := X"24060110";
        ram_buffer(66314) := X"00002821";
        ram_buffer(66315) := X"02002021";
        ram_buffer(66316) := X"0C02801D";
        ram_buffer(66317) := X"A3A00156";
        ram_buffer(66318) := X"24140001";
        ram_buffer(66319) := X"02002021";
        ram_buffer(66320) := X"2406003C";
        ram_buffer(66321) := X"00002821";
        ram_buffer(66322) := X"A214003C";
        ram_buffer(66323) := X"0C02801D";
        ram_buffer(66324) := X"A214003D";
        ram_buffer(66325) := X"02202821";
        ram_buffer(66326) := X"24060027";
        ram_buffer(66327) := X"0C02CCBF";
        ram_buffer(66328) := X"02002021";
        ram_buffer(66329) := X"97A20158";
        ram_buffer(66330) := X"AE000028";
        ram_buffer(66331) := X"A6020038";
        ram_buffer(66332) := X"93A20157";
        ram_buffer(66333) := X"A2140036";
        ram_buffer(66334) := X"A2020037";
        ram_buffer(66335) := X"00002821";
        ram_buffer(66336) := X"0C02FD29";
        ram_buffer(66337) := X"02002021";
        ram_buffer(66338) := X"8E140040";
        ram_buffer(66339) := X"24060080";
        ram_buffer(66340) := X"02402821";
        ram_buffer(66341) := X"2604004C";
        ram_buffer(66342) := X"AE140028";
        ram_buffer(66343) := X"AE000048";
        ram_buffer(66344) := X"0C030956";
        ram_buffer(66345) := X"A200004C";
        ram_buffer(66346) := X"82630000";
        ram_buffer(66347) := X"24020061";
        ram_buffer(66348) := X"10620017";
        ram_buffer(66349) := X"02001021";
        ram_buffer(66350) := X"1000FFCE";
        ram_buffer(66351) := X"00000000";
        ram_buffer(66352) := X"0C0300CE";
        ram_buffer(66353) := X"00000000";
        ram_buffer(66354) := X"1000FF95";
        ram_buffer(66355) := X"24050001";
        ram_buffer(66356) := X"02203821";
        ram_buffer(66357) := X"02803021";
        ram_buffer(66358) := X"02402821";
        ram_buffer(66359) := X"02A02021";
        ram_buffer(66360) := X"0C030030";
        ram_buffer(66361) := X"A3A00154";
        ram_buffer(66362) := X"1440FFA0";
        ram_buffer(66363) := X"02203821";
        ram_buffer(66364) := X"93A20154";
        ram_buffer(66365) := X"00000000";
        ram_buffer(66366) := X"1440002E";
        ram_buffer(66367) := X"00000000";
        ram_buffer(66368) := X"0C0301F5";
        ram_buffer(66369) := X"02402021";
        ram_buffer(66370) := X"1000FF98";
        ram_buffer(66371) := X"02203821";
        ram_buffer(66372) := X"8E110030";
        ram_buffer(66373) := X"02802821";
        ram_buffer(66374) := X"02002021";
        ram_buffer(66375) := X"0C02FD29";
        ram_buffer(66376) := X"AE110048";
        ram_buffer(66377) := X"96020038";
        ram_buffer(66378) := X"00000000";
        ram_buffer(66379) := X"2442FFFD";
        ram_buffer(66380) := X"0222102A";
        ram_buffer(66381) := X"1440000E";
        ram_buffer(66382) := X"24120004";
        ram_buffer(66383) := X"8E0200CC";
        ram_buffer(66384) := X"00000000";
        ram_buffer(66385) := X"8C450000";
        ram_buffer(66386) := X"0C02FD29";
        ram_buffer(66387) := X"02002021";
        ram_buffer(66388) := X"96020038";
        ram_buffer(66389) := X"00000000";
        ram_buffer(66390) := X"02421823";
        ram_buffer(66391) := X"02238821";
        ram_buffer(66392) := X"2442FFFD";
        ram_buffer(66393) := X"0222102A";
        ram_buffer(66394) := X"1040FFF4";
        ram_buffer(66395) := X"00000000";
        ram_buffer(66396) := X"AE110044";
        ram_buffer(66397) := X"1000FF9F";
        ram_buffer(66398) := X"02001021";
        ram_buffer(66399) := X"0C027A4D";
        ram_buffer(66400) := X"02002021";
        ram_buffer(66401) := X"0C030730";
        ram_buffer(66402) := X"00000000";
        ram_buffer(66403) := X"24030002";
        ram_buffer(66404) := X"AC430000";
        ram_buffer(66405) := X"1000FF97";
        ram_buffer(66406) := X"00001021";
        ram_buffer(66407) := X"0C030730";
        ram_buffer(66408) := X"00000000";
        ram_buffer(66409) := X"2403000C";
        ram_buffer(66410) := X"AC430000";
        ram_buffer(66411) := X"1000FF91";
        ram_buffer(66412) := X"00001021";
        ram_buffer(66413) := X"0C027A4D";
        ram_buffer(66414) := X"02002021";
        ram_buffer(66415) := X"0C030730";
        ram_buffer(66416) := X"00000000";
        ram_buffer(66417) := X"24030015";
        ram_buffer(66418) := X"AC430000";
        ram_buffer(66419) := X"1000FF89";
        ram_buffer(66420) := X"00001021";
        ram_buffer(66421) := X"3C05100D";
        ram_buffer(66422) := X"27BDFFE8";
        ram_buffer(66423) := X"AFBF0014";
        ram_buffer(66424) := X"0C0302B9";
        ram_buffer(66425) := X"24A5B3F4";
        ram_buffer(66426) := X"10400009";
        ram_buffer(66427) := X"24030001";
        ram_buffer(66428) := X"A0430034";
        ram_buffer(66429) := X"0C03013B";
        ram_buffer(66430) := X"00402021";
        ram_buffer(66431) := X"00001021";
        ram_buffer(66432) := X"8FBF0014";
        ram_buffer(66433) := X"00000000";
        ram_buffer(66434) := X"03E00008";
        ram_buffer(66435) := X"27BD0018";
        ram_buffer(66436) := X"1000FFFB";
        ram_buffer(66437) := X"2402FFFF";
        ram_buffer(66438) := X"8C820030";
        ram_buffer(66439) := X"03E00008";
        ram_buffer(66440) := X"00000000";
        ram_buffer(66441) := X"27BDFFD0";
        ram_buffer(66442) := X"8C820048";
        ram_buffer(66443) := X"AFB50028";
        ram_buffer(66444) := X"AFB30020";
        ram_buffer(66445) := X"AFB2001C";
        ram_buffer(66446) := X"AFB10018";
        ram_buffer(66447) := X"AFB00014";
        ram_buffer(66448) := X"AFBF002C";
        ram_buffer(66449) := X"AFB40024";
        ram_buffer(66450) := X"00808021";
        ram_buffer(66451) := X"00A09021";
        ram_buffer(66452) := X"24B5003C";
        ram_buffer(66453) := X"2411FFFF";
        ram_buffer(66454) := X"24130001";
        ram_buffer(66455) := X"0240A021";
        ram_buffer(66456) := X"8E030030";
        ram_buffer(66457) := X"00000000";
        ram_buffer(66458) := X"0043102B";
        ram_buffer(66459) := X"14400005";
        ram_buffer(66460) := X"02002021";
        ram_buffer(66461) := X"92020034";
        ram_buffer(66462) := X"00000000";
        ram_buffer(66463) := X"10400027";
        ram_buffer(66464) := X"2402FFFF";
        ram_buffer(66465) := X"96020038";
        ram_buffer(66466) := X"8E030044";
        ram_buffer(66467) := X"2442FFFC";
        ram_buffer(66468) := X"0062102B";
        ram_buffer(66469) := X"1440000A";
        ram_buffer(66470) := X"00000000";
        ram_buffer(66471) := X"8E0200CC";
        ram_buffer(66472) := X"00000000";
        ram_buffer(66473) := X"8C420000";
        ram_buffer(66474) := X"00000000";
        ram_buffer(66475) := X"1051001A";
        ram_buffer(66476) := X"00402821";
        ram_buffer(66477) := X"0C02FD29";
        ram_buffer(66478) := X"00000000";
        ram_buffer(66479) := X"8E030044";
        ram_buffer(66480) := X"8E0200CC";
        ram_buffer(66481) := X"24640001";
        ram_buffer(66482) := X"AE040044";
        ram_buffer(66483) := X"00431821";
        ram_buffer(66484) := X"90620004";
        ram_buffer(66485) := X"26940001";
        ram_buffer(66486) := X"A282FFFF";
        ram_buffer(66487) := X"8E020048";
        ram_buffer(66488) := X"00000000";
        ram_buffer(66489) := X"24420001";
        ram_buffer(66490) := X"16B4FFDD";
        ram_buffer(66491) := X"AE020048";
        ram_buffer(66492) := X"8E430028";
        ram_buffer(66493) := X"00000000";
        ram_buffer(66494) := X"10710007";
        ram_buffer(66495) := X"00000000";
        ram_buffer(66496) := X"92430036";
        ram_buffer(66497) := X"00000000";
        ram_buffer(66498) := X"1473FFD5";
        ram_buffer(66499) := X"0240A021";
        ram_buffer(66500) := X"10000002";
        ram_buffer(66501) := X"00001021";
        ram_buffer(66502) := X"2402FFFF";
        ram_buffer(66503) := X"8FBF002C";
        ram_buffer(66504) := X"8FB50028";
        ram_buffer(66505) := X"8FB40024";
        ram_buffer(66506) := X"8FB30020";
        ram_buffer(66507) := X"8FB2001C";
        ram_buffer(66508) := X"8FB10018";
        ram_buffer(66509) := X"8FB00014";
        ram_buffer(66510) := X"03E00008";
        ram_buffer(66511) := X"27BD0030";
        ram_buffer(66512) := X"27BDFFC0";
        ram_buffer(66513) := X"AFB0001C";
        ram_buffer(66514) := X"3C10100C";
        ram_buffer(66515) := X"AFB50030";
        ram_buffer(66516) := X"00A0A821";
        ram_buffer(66517) := X"26057BF0";
        ram_buffer(66518) := X"AFB70038";
        ram_buffer(66519) := X"AFB60034";
        ram_buffer(66520) := X"AFBF003C";
        ram_buffer(66521) := X"AFB4002C";
        ram_buffer(66522) := X"AFB30028";
        ram_buffer(66523) := X"AFB20024";
        ram_buffer(66524) := X"AFB10020";
        ram_buffer(66525) := X"0080B821";
        ram_buffer(66526) := X"0C02716A";
        ram_buffer(66527) := X"00C0B021";
        ram_buffer(66528) := X"1040005B";
        ram_buffer(66529) := X"26057BF0";
        ram_buffer(66530) := X"02A02021";
        ram_buffer(66531) := X"0C02716A";
        ram_buffer(66532) := X"00408821";
        ram_buffer(66533) := X"1040005D";
        ram_buffer(66534) := X"00409021";
        ram_buffer(66535) := X"24060002";
        ram_buffer(66536) := X"00002821";
        ram_buffer(66537) := X"0C02758D";
        ram_buffer(66538) := X"02202021";
        ram_buffer(66539) := X"0C03074B";
        ram_buffer(66540) := X"02202021";
        ram_buffer(66541) := X"00408021";
        ram_buffer(66542) := X"00002821";
        ram_buffer(66543) := X"00003021";
        ram_buffer(66544) := X"0C02758D";
        ram_buffer(66545) := X"02202021";
        ram_buffer(66546) := X"0C027A3D";
        ram_buffer(66547) := X"02002021";
        ram_buffer(66548) := X"00409821";
        ram_buffer(66549) := X"0C027A3D";
        ram_buffer(66550) := X"02002021";
        ram_buffer(66551) := X"02203821";
        ram_buffer(66552) := X"02003021";
        ram_buffer(66553) := X"24050001";
        ram_buffer(66554) := X"02602021";
        ram_buffer(66555) := X"0C0272E9";
        ram_buffer(66556) := X"0040A021";
        ram_buffer(66557) := X"16020023";
        ram_buffer(66558) := X"3C05100D";
        ram_buffer(66559) := X"0C026DBB";
        ram_buffer(66560) := X"02202021";
        ram_buffer(66561) := X"02403821";
        ram_buffer(66562) := X"02003021";
        ram_buffer(66563) := X"24050001";
        ram_buffer(66564) := X"0C0272E9";
        ram_buffer(66565) := X"02802021";
        ram_buffer(66566) := X"16020024";
        ram_buffer(66567) := X"3C05100D";
        ram_buffer(66568) := X"0C026DBB";
        ram_buffer(66569) := X"02402021";
        ram_buffer(66570) := X"02003021";
        ram_buffer(66571) := X"02802821";
        ram_buffer(66572) := X"0C0307E3";
        ram_buffer(66573) := X"02602021";
        ram_buffer(66574) := X"14400026";
        ram_buffer(66575) := X"00408021";
        ram_buffer(66576) := X"3C05100D";
        ram_buffer(66577) := X"2406000A";
        ram_buffer(66578) := X"24A5B46C";
        ram_buffer(66579) := X"0C027F93";
        ram_buffer(66580) := X"02C02021";
        ram_buffer(66581) := X"8FBF003C";
        ram_buffer(66582) := X"02001021";
        ram_buffer(66583) := X"8FB70038";
        ram_buffer(66584) := X"8FB60034";
        ram_buffer(66585) := X"8FB50030";
        ram_buffer(66586) := X"8FB4002C";
        ram_buffer(66587) := X"8FB30028";
        ram_buffer(66588) := X"8FB20024";
        ram_buffer(66589) := X"8FB10020";
        ram_buffer(66590) := X"8FB0001C";
        ram_buffer(66591) := X"03E00008";
        ram_buffer(66592) := X"27BD0040";
        ram_buffer(66593) := X"AFB00010";
        ram_buffer(66594) := X"00403821";
        ram_buffer(66595) := X"02E03021";
        ram_buffer(66596) := X"24A5B414";
        ram_buffer(66597) := X"0C0283DB";
        ram_buffer(66598) := X"02C02021";
        ram_buffer(66599) := X"0C026DBB";
        ram_buffer(66600) := X"02202021";
        ram_buffer(66601) := X"1000FFEB";
        ram_buffer(66602) := X"2410FFFF";
        ram_buffer(66603) := X"AFB00010";
        ram_buffer(66604) := X"00403821";
        ram_buffer(66605) := X"02A03021";
        ram_buffer(66606) := X"24A5B414";
        ram_buffer(66607) := X"0C0283DB";
        ram_buffer(66608) := X"02C02021";
        ram_buffer(66609) := X"0C026DBB";
        ram_buffer(66610) := X"02402021";
        ram_buffer(66611) := X"1000FFE1";
        ram_buffer(66612) := X"2410FFFF";
        ram_buffer(66613) := X"3C05100D";
        ram_buffer(66614) := X"2406001A";
        ram_buffer(66615) := X"24A5B450";
        ram_buffer(66616) := X"0C027F93";
        ram_buffer(66617) := X"02C02021";
        ram_buffer(66618) := X"1000FFDA";
        ram_buffer(66619) := X"2410FFFF";
        ram_buffer(66620) := X"3C05100D";
        ram_buffer(66621) := X"02E03021";
        ram_buffer(66622) := X"24A5B3F8";
        ram_buffer(66623) := X"0C0283DB";
        ram_buffer(66624) := X"02C02021";
        ram_buffer(66625) := X"1000FFD3";
        ram_buffer(66626) := X"2410FFFF";
        ram_buffer(66627) := X"3C05100D";
        ram_buffer(66628) := X"02C02021";
        ram_buffer(66629) := X"02A03021";
        ram_buffer(66630) := X"0C0283DB";
        ram_buffer(66631) := X"24A5B3F8";
        ram_buffer(66632) := X"0C026DBB";
        ram_buffer(66633) := X"00002021";
        ram_buffer(66634) := X"1000FFCA";
        ram_buffer(66635) := X"2410FFFF";
        ram_buffer(66636) := X"27BDFEF8";
        ram_buffer(66637) := X"00802821";
        ram_buffer(66638) := X"AFB200E8";
        ram_buffer(66639) := X"00809021";
        ram_buffer(66640) := X"3C04100D";
        ram_buffer(66641) := X"2484B478";
        ram_buffer(66642) := X"AFBF0104";
        ram_buffer(66643) := X"AFBE0100";
        ram_buffer(66644) := X"AFB700FC";
        ram_buffer(66645) := X"AFB600F8";
        ram_buffer(66646) := X"AFB500F4";
        ram_buffer(66647) := X"AFB400F0";
        ram_buffer(66648) := X"AFB300EC";
        ram_buffer(66649) := X"AFB100E4";
        ram_buffer(66650) := X"0C028116";
        ram_buffer(66651) := X"AFB000E0";
        ram_buffer(66652) := X"3C05100D";
        ram_buffer(66653) := X"24A58F90";
        ram_buffer(66654) := X"0C0302B9";
        ram_buffer(66655) := X"02402021";
        ram_buffer(66656) := X"10400074";
        ram_buffer(66657) := X"3C16100D";
        ram_buffer(66658) := X"0040B821";
        ram_buffer(66659) := X"3C15100D";
        ram_buffer(66660) := X"26C2B3F0";
        ram_buffer(66661) := X"AFA200D0";
        ram_buffer(66662) := X"26A2B4BC";
        ram_buffer(66663) := X"3C13100D";
        ram_buffer(66664) := X"AFA200D4";
        ram_buffer(66665) := X"3C02100D";
        ram_buffer(66666) := X"3C14100D";
        ram_buffer(66667) := X"2673B4E4";
        ram_buffer(66668) := X"3C1E100D";
        ram_buffer(66669) := X"AFA200D8";
        ram_buffer(66670) := X"2410FFFF";
        ram_buffer(66671) := X"27B500CC";
        ram_buffer(66672) := X"24110001";
        ram_buffer(66673) := X"8EE20048";
        ram_buffer(66674) := X"27B60090";
        ram_buffer(66675) := X"8EE50030";
        ram_buffer(66676) := X"00000000";
        ram_buffer(66677) := X"0045102B";
        ram_buffer(66678) := X"14400005";
        ram_buffer(66679) := X"02E02021";
        ram_buffer(66680) := X"92E20034";
        ram_buffer(66681) := X"00000000";
        ram_buffer(66682) := X"10400040";
        ram_buffer(66683) := X"00000000";
        ram_buffer(66684) := X"96E20038";
        ram_buffer(66685) := X"8EE50044";
        ram_buffer(66686) := X"2442FFFC";
        ram_buffer(66687) := X"00A2102B";
        ram_buffer(66688) := X"1440000A";
        ram_buffer(66689) := X"00000000";
        ram_buffer(66690) := X"8EE200CC";
        ram_buffer(66691) := X"00000000";
        ram_buffer(66692) := X"8C420000";
        ram_buffer(66693) := X"00000000";
        ram_buffer(66694) := X"10500034";
        ram_buffer(66695) := X"00402821";
        ram_buffer(66696) := X"0C02FD29";
        ram_buffer(66697) := X"00000000";
        ram_buffer(66698) := X"8EE50044";
        ram_buffer(66699) := X"8EE200CC";
        ram_buffer(66700) := X"24A40001";
        ram_buffer(66701) := X"AEE40044";
        ram_buffer(66702) := X"00452821";
        ram_buffer(66703) := X"90A20004";
        ram_buffer(66704) := X"26D60001";
        ram_buffer(66705) := X"A2C2FFFF";
        ram_buffer(66706) := X"8EE20048";
        ram_buffer(66707) := X"00000000";
        ram_buffer(66708) := X"24420001";
        ram_buffer(66709) := X"16D5FFDD";
        ram_buffer(66710) := X"AEE20048";
        ram_buffer(66711) := X"8FA400B8";
        ram_buffer(66712) := X"00000000";
        ram_buffer(66713) := X"10900022";
        ram_buffer(66714) := X"2684B4A0";
        ram_buffer(66715) := X"93A400C6";
        ram_buffer(66716) := X"00000000";
        ram_buffer(66717) := X"1491FFD4";
        ram_buffer(66718) := X"02402821";
        ram_buffer(66719) := X"00003021";
        ram_buffer(66720) := X"0C028116";
        ram_buffer(66721) := X"2684B4A0";
        ram_buffer(66722) := X"8FA600C0";
        ram_buffer(66723) := X"27A50090";
        ram_buffer(66724) := X"0C028116";
        ram_buffer(66725) := X"02602021";
        ram_buffer(66726) := X"93A200C4";
        ram_buffer(66727) := X"00000000";
        ram_buffer(66728) := X"1040FFC8";
        ram_buffer(66729) := X"00000000";
        ram_buffer(66730) := X"8FA500D0";
        ram_buffer(66731) := X"0C02CC2F";
        ram_buffer(66732) := X"02402021";
        ram_buffer(66733) := X"14400020";
        ram_buffer(66734) := X"27B00010";
        ram_buffer(66735) := X"8FA500D4";
        ram_buffer(66736) := X"27A60090";
        ram_buffer(66737) := X"0C0283DB";
        ram_buffer(66738) := X"02002021";
        ram_buffer(66739) := X"8FA200D8";
        ram_buffer(66740) := X"02002821";
        ram_buffer(66741) := X"0C028116";
        ram_buffer(66742) := X"2444B4C8";
        ram_buffer(66743) := X"0C03044C";
        ram_buffer(66744) := X"02002021";
        ram_buffer(66745) := X"1000FFB5";
        ram_buffer(66746) := X"2410FFFF";
        ram_buffer(66747) := X"2684B4A0";
        ram_buffer(66748) := X"2406FFFF";
        ram_buffer(66749) := X"0C028116";
        ram_buffer(66750) := X"02402821";
        ram_buffer(66751) := X"0C03013B";
        ram_buffer(66752) := X"02E02021";
        ram_buffer(66753) := X"8FBF0104";
        ram_buffer(66754) := X"8FBE0100";
        ram_buffer(66755) := X"8FB700FC";
        ram_buffer(66756) := X"8FB600F8";
        ram_buffer(66757) := X"8FB500F4";
        ram_buffer(66758) := X"8FB400F0";
        ram_buffer(66759) := X"8FB300EC";
        ram_buffer(66760) := X"8FB200E8";
        ram_buffer(66761) := X"8FB100E4";
        ram_buffer(66762) := X"8FB000E0";
        ram_buffer(66763) := X"00001021";
        ram_buffer(66764) := X"03E00008";
        ram_buffer(66765) := X"27BD0108";
        ram_buffer(66766) := X"27A70090";
        ram_buffer(66767) := X"02403021";
        ram_buffer(66768) := X"27C5B4C0";
        ram_buffer(66769) := X"0C0283DB";
        ram_buffer(66770) := X"02002021";
        ram_buffer(66771) := X"1000FFDF";
        ram_buffer(66772) := X"00000000";
        ram_buffer(66773) := X"3C04100D";
        ram_buffer(66774) := X"02402821";
        ram_buffer(66775) := X"0C028116";
        ram_buffer(66776) := X"2484B48C";
        ram_buffer(66777) := X"1000FFE7";
        ram_buffer(66778) := X"00000000";
        ram_buffer(66779) := X"27BDFF98";
        ram_buffer(66780) := X"24050001";
        ram_buffer(66781) := X"24041388";
        ram_buffer(66782) := X"AFBF0064";
        ram_buffer(66783) := X"AFBE0060";
        ram_buffer(66784) := X"AFB7005C";
        ram_buffer(66785) := X"AFB60058";
        ram_buffer(66786) := X"AFB50054";
        ram_buffer(66787) := X"AFB40050";
        ram_buffer(66788) := X"AFB3004C";
        ram_buffer(66789) := X"AFB20048";
        ram_buffer(66790) := X"AFB10044";
        ram_buffer(66791) := X"0C03071E";
        ram_buffer(66792) := X"AFB00040";
        ram_buffer(66793) := X"104001A2";
        ram_buffer(66794) := X"00408021";
        ram_buffer(66795) := X"00402021";
        ram_buffer(66796) := X"2405001A";
        ram_buffer(66797) := X"00001021";
        ram_buffer(66798) := X"24060FA0";
        ram_buffer(66799) := X"14A00002";
        ram_buffer(66800) := X"0045001A";
        ram_buffer(66801) := X"0007000D";
        ram_buffer(66802) := X"24840001";
        ram_buffer(66803) := X"24420001";
        ram_buffer(66804) := X"00001810";
        ram_buffer(66805) := X"24630041";
        ram_buffer(66806) := X"1446FFF8";
        ram_buffer(66807) := X"A083FFFF";
        ram_buffer(66808) := X"3C02100D";
        ram_buffer(66809) := X"3C04100D";
        ram_buffer(66810) := X"2445B3F4";
        ram_buffer(66811) := X"2484B4F4";
        ram_buffer(66812) := X"0C0302B9";
        ram_buffer(66813) := X"AFA20034";
        ram_buffer(66814) := X"10400004";
        ram_buffer(66815) := X"24030001";
        ram_buffer(66816) := X"A0430034";
        ram_buffer(66817) := X"0C03013B";
        ram_buffer(66818) := X"00402021";
        ram_buffer(66819) := X"8FA30034";
        ram_buffer(66820) := X"3C02100D";
        ram_buffer(66821) := X"2465B3F4";
        ram_buffer(66822) := X"2444B4EC";
        ram_buffer(66823) := X"0C0302B9";
        ram_buffer(66824) := X"AFA2003C";
        ram_buffer(66825) := X"10400004";
        ram_buffer(66826) := X"24030001";
        ram_buffer(66827) := X"A0430034";
        ram_buffer(66828) := X"0C03013B";
        ram_buffer(66829) := X"00402021";
        ram_buffer(66830) := X"3C02100D";
        ram_buffer(66831) := X"3C03100D";
        ram_buffer(66832) := X"2445B4F8";
        ram_buffer(66833) := X"2464B4FC";
        ram_buffer(66834) := X"AFA20020";
        ram_buffer(66835) := X"0C0302B9";
        ram_buffer(66836) := X"AFA30024";
        ram_buffer(66837) := X"10400176";
        ram_buffer(66838) := X"00408821";
        ram_buffer(66839) := X"24020001";
        ram_buffer(66840) := X"A222003D";
        ram_buffer(66841) := X"02009821";
        ram_buffer(66842) := X"0000A021";
        ram_buffer(66843) := X"2415FFFF";
        ram_buffer(66844) := X"10000016";
        ram_buffer(66845) := X"24120001";
        ram_buffer(66846) := X"0C02FD29";
        ram_buffer(66847) := X"02202021";
        ram_buffer(66848) := X"8E220040";
        ram_buffer(66849) := X"00000000";
        ram_buffer(66850) := X"10550024";
        ram_buffer(66851) := X"00000000";
        ram_buffer(66852) := X"8E230044";
        ram_buffer(66853) := X"A232003D";
        ram_buffer(66854) := X"24640001";
        ram_buffer(66855) := X"8E2200CC";
        ram_buffer(66856) := X"AE240044";
        ram_buffer(66857) := X"92640000";
        ram_buffer(66858) := X"00431821";
        ram_buffer(66859) := X"A0640004";
        ram_buffer(66860) := X"8E220048";
        ram_buffer(66861) := X"26940001";
        ram_buffer(66862) := X"24420001";
        ram_buffer(66863) := X"2A830FA0";
        ram_buffer(66864) := X"26730001";
        ram_buffer(66865) := X"10600016";
        ram_buffer(66866) := X"AE220048";
        ram_buffer(66867) := X"96220038";
        ram_buffer(66868) := X"8E230044";
        ram_buffer(66869) := X"2442FFFC";
        ram_buffer(66870) := X"0062102B";
        ram_buffer(66871) := X"1440FFEF";
        ram_buffer(66872) := X"24640001";
        ram_buffer(66873) := X"8E2200CC";
        ram_buffer(66874) := X"00000000";
        ram_buffer(66875) := X"8C450000";
        ram_buffer(66876) := X"00000000";
        ram_buffer(66877) := X"14B5FFE0";
        ram_buffer(66878) := X"00000000";
        ram_buffer(66879) := X"AC400000";
        ram_buffer(66880) := X"00002821";
        ram_buffer(66881) := X"0C02FD29";
        ram_buffer(66882) := X"02202021";
        ram_buffer(66883) := X"8E220040";
        ram_buffer(66884) := X"00000000";
        ram_buffer(66885) := X"1455FFDE";
        ram_buffer(66886) := X"00000000";
        ram_buffer(66887) := X"8E220048";
        ram_buffer(66888) := X"8E230030";
        ram_buffer(66889) := X"24040001";
        ram_buffer(66890) := X"0062182B";
        ram_buffer(66891) := X"A224003D";
        ram_buffer(66892) := X"10600002";
        ram_buffer(66893) := X"A224003C";
        ram_buffer(66894) := X"AE220030";
        ram_buffer(66895) := X"0C03013B";
        ram_buffer(66896) := X"02202021";
        ram_buffer(66897) := X"02002021";
        ram_buffer(66898) := X"24061388";
        ram_buffer(66899) := X"0C02801D";
        ram_buffer(66900) := X"00002821";
        ram_buffer(66901) := X"3C02100D";
        ram_buffer(66902) := X"AFA20038";
        ram_buffer(66903) := X"24458F90";
        ram_buffer(66904) := X"8FA20024";
        ram_buffer(66905) := X"0C0302B9";
        ram_buffer(66906) := X"2444B4FC";
        ram_buffer(66907) := X"10400130";
        ram_buffer(66908) := X"00408821";
        ram_buffer(66909) := X"8C420048";
        ram_buffer(66910) := X"26141388";
        ram_buffer(66911) := X"02009021";
        ram_buffer(66912) := X"1000001C";
        ram_buffer(66913) := X"2413FFFF";
        ram_buffer(66914) := X"96220038";
        ram_buffer(66915) := X"8E230044";
        ram_buffer(66916) := X"2442FFFC";
        ram_buffer(66917) := X"0062102B";
        ram_buffer(66918) := X"1440000A";
        ram_buffer(66919) := X"00000000";
        ram_buffer(66920) := X"8E2200CC";
        ram_buffer(66921) := X"00000000";
        ram_buffer(66922) := X"8C420000";
        ram_buffer(66923) := X"00000000";
        ram_buffer(66924) := X"10530019";
        ram_buffer(66925) := X"00402821";
        ram_buffer(66926) := X"0C02FD29";
        ram_buffer(66927) := X"00000000";
        ram_buffer(66928) := X"8E230044";
        ram_buffer(66929) := X"8E2200CC";
        ram_buffer(66930) := X"24640001";
        ram_buffer(66931) := X"AE240044";
        ram_buffer(66932) := X"00431821";
        ram_buffer(66933) := X"90620004";
        ram_buffer(66934) := X"00000000";
        ram_buffer(66935) := X"A242FFFF";
        ram_buffer(66936) := X"8E220048";
        ram_buffer(66937) := X"00000000";
        ram_buffer(66938) := X"24420001";
        ram_buffer(66939) := X"1292000A";
        ram_buffer(66940) := X"AE220048";
        ram_buffer(66941) := X"8E230030";
        ram_buffer(66942) := X"26520001";
        ram_buffer(66943) := X"0043102B";
        ram_buffer(66944) := X"1440FFE1";
        ram_buffer(66945) := X"02202021";
        ram_buffer(66946) := X"92220034";
        ram_buffer(66947) := X"00000000";
        ram_buffer(66948) := X"1440FFDD";
        ram_buffer(66949) := X"00000000";
        ram_buffer(66950) := X"0C03013B";
        ram_buffer(66951) := X"02202021";
        ram_buffer(66952) := X"3C04100D";
        ram_buffer(66953) := X"02002821";
        ram_buffer(66954) := X"0C028116";
        ram_buffer(66955) := X"2484B514";
        ram_buffer(66956) := X"3C02100D";
        ram_buffer(66957) := X"2444B3F0";
        ram_buffer(66958) := X"0C03044C";
        ram_buffer(66959) := X"AFA20030";
        ram_buffer(66960) := X"3C02100D";
        ram_buffer(66961) := X"AFA2002C";
        ram_buffer(66962) := X"2455B524";
        ram_buffer(66963) := X"8FA20020";
        ram_buffer(66964) := X"3C16100D";
        ram_buffer(66965) := X"2442B4F8";
        ram_buffer(66966) := X"3C03100D";
        ram_buffer(66967) := X"AFA20018";
        ram_buffer(66968) := X"26C2B534";
        ram_buffer(66969) := X"00009821";
        ram_buffer(66970) := X"AFA30028";
        ram_buffer(66971) := X"24110001";
        ram_buffer(66972) := X"AFA2001C";
        ram_buffer(66973) := X"8FA20028";
        ram_buffer(66974) := X"02002021";
        ram_buffer(66975) := X"2445B51C";
        ram_buffer(66976) := X"0C0283DB";
        ram_buffer(66977) := X"02603021";
        ram_buffer(66978) := X"8FA20034";
        ram_buffer(66979) := X"02002021";
        ram_buffer(66980) := X"0C0302B9";
        ram_buffer(66981) := X"2445B3F4";
        ram_buffer(66982) := X"10400005";
        ram_buffer(66983) := X"00009021";
        ram_buffer(66984) := X"A0510034";
        ram_buffer(66985) := X"0C03013B";
        ram_buffer(66986) := X"00402021";
        ram_buffer(66987) := X"00009021";
        ram_buffer(66988) := X"02603821";
        ram_buffer(66989) := X"02603021";
        ram_buffer(66990) := X"02A02821";
        ram_buffer(66991) := X"02002021";
        ram_buffer(66992) := X"0C0283DB";
        ram_buffer(66993) := X"AFB20010";
        ram_buffer(66994) := X"8FA50018";
        ram_buffer(66995) := X"0C0302B9";
        ram_buffer(66996) := X"02002021";
        ram_buffer(66997) := X"1040003E";
        ram_buffer(66998) := X"0040B821";
        ram_buffer(66999) := X"8FA5001C";
        ram_buffer(67000) := X"02403821";
        ram_buffer(67001) := X"02603021";
        ram_buffer(67002) := X"0C0283DB";
        ram_buffer(67003) := X"02002021";
        ram_buffer(67004) := X"0200A021";
        ram_buffer(67005) := X"A2F1003D";
        ram_buffer(67006) := X"0000B021";
        ram_buffer(67007) := X"10000017";
        ram_buffer(67008) := X"241EFFFF";
        ram_buffer(67009) := X"0C02FD29";
        ram_buffer(67010) := X"02E02021";
        ram_buffer(67011) := X"8EE20040";
        ram_buffer(67012) := X"00000000";
        ram_buffer(67013) := X"105E0025";
        ram_buffer(67014) := X"00000000";
        ram_buffer(67015) := X"8EE40044";
        ram_buffer(67016) := X"A2F1003D";
        ram_buffer(67017) := X"24850001";
        ram_buffer(67018) := X"8EE200CC";
        ram_buffer(67019) := X"AEE50044";
        ram_buffer(67020) := X"92850000";
        ram_buffer(67021) := X"00442021";
        ram_buffer(67022) := X"A0850004";
        ram_buffer(67023) := X"8EE20048";
        ram_buffer(67024) := X"26D60001";
        ram_buffer(67025) := X"24420001";
        ram_buffer(67026) := X"2AC40008";
        ram_buffer(67027) := X"26860001";
        ram_buffer(67028) := X"10800017";
        ram_buffer(67029) := X"AEE20048";
        ram_buffer(67030) := X"00C0A021";
        ram_buffer(67031) := X"96E20038";
        ram_buffer(67032) := X"8EE40044";
        ram_buffer(67033) := X"2442FFFC";
        ram_buffer(67034) := X"0082102B";
        ram_buffer(67035) := X"1440FFEE";
        ram_buffer(67036) := X"24850001";
        ram_buffer(67037) := X"8EE200CC";
        ram_buffer(67038) := X"00000000";
        ram_buffer(67039) := X"8C450000";
        ram_buffer(67040) := X"00000000";
        ram_buffer(67041) := X"14BEFFDF";
        ram_buffer(67042) := X"00000000";
        ram_buffer(67043) := X"AC400000";
        ram_buffer(67044) := X"00002821";
        ram_buffer(67045) := X"0C02FD29";
        ram_buffer(67046) := X"02E02021";
        ram_buffer(67047) := X"8EE20040";
        ram_buffer(67048) := X"00000000";
        ram_buffer(67049) := X"145EFFDD";
        ram_buffer(67050) := X"00000000";
        ram_buffer(67051) := X"8EE20048";
        ram_buffer(67052) := X"8EE40030";
        ram_buffer(67053) := X"A2F1003D";
        ram_buffer(67054) := X"0082202B";
        ram_buffer(67055) := X"10800002";
        ram_buffer(67056) := X"A2F1003C";
        ram_buffer(67057) := X"AEE20030";
        ram_buffer(67058) := X"0C03013B";
        ram_buffer(67059) := X"02E02021";
        ram_buffer(67060) := X"26520001";
        ram_buffer(67061) := X"24020005";
        ram_buffer(67062) := X"1642FFB6";
        ram_buffer(67063) := X"02603821";
        ram_buffer(67064) := X"26730001";
        ram_buffer(67065) := X"1672FFA3";
        ram_buffer(67066) := X"3C04100D";
        ram_buffer(67067) := X"0C0301F5";
        ram_buffer(67068) := X"2484B540";
        ram_buffer(67069) := X"8FA20030";
        ram_buffer(67070) := X"0C03044C";
        ram_buffer(67071) := X"2444B3F0";
        ram_buffer(67072) := X"8FA20020";
        ram_buffer(67073) := X"3C04100D";
        ram_buffer(67074) := X"2445B4F8";
        ram_buffer(67075) := X"0C0302B9";
        ram_buffer(67076) := X"2484B550";
        ram_buffer(67077) := X"10400004";
        ram_buffer(67078) := X"00000000";
        ram_buffer(67079) := X"3C04100D";
        ram_buffer(67080) := X"0C028186";
        ram_buffer(67081) := X"2484B564";
        ram_buffer(67082) := X"8FA2002C";
        ram_buffer(67083) := X"3C14100D";
        ram_buffer(67084) := X"2453B524";
        ram_buffer(67085) := X"8FA20038";
        ram_buffer(67086) := X"00008821";
        ram_buffer(67087) := X"24528F90";
        ram_buffer(67088) := X"2682B56C";
        ram_buffer(67089) := X"AFA20018";
        ram_buffer(67090) := X"0000B821";
        ram_buffer(67091) := X"02203821";
        ram_buffer(67092) := X"02203021";
        ram_buffer(67093) := X"02602821";
        ram_buffer(67094) := X"02002021";
        ram_buffer(67095) := X"0C0283DB";
        ram_buffer(67096) := X"AFB70010";
        ram_buffer(67097) := X"02402821";
        ram_buffer(67098) := X"0C0302B9";
        ram_buffer(67099) := X"02002021";
        ram_buffer(67100) := X"10400031";
        ram_buffer(67101) := X"0040B021";
        ram_buffer(67102) := X"8C420048";
        ram_buffer(67103) := X"0200A821";
        ram_buffer(67104) := X"0000F021";
        ram_buffer(67105) := X"241401F4";
        ram_buffer(67106) := X"8EC30030";
        ram_buffer(67107) := X"00000000";
        ram_buffer(67108) := X"0043102B";
        ram_buffer(67109) := X"14400005";
        ram_buffer(67110) := X"02C02021";
        ram_buffer(67111) := X"92C20034";
        ram_buffer(67112) := X"00000000";
        ram_buffer(67113) := X"1040001C";
        ram_buffer(67114) := X"00000000";
        ram_buffer(67115) := X"96C20038";
        ram_buffer(67116) := X"8EC30044";
        ram_buffer(67117) := X"2442FFFC";
        ram_buffer(67118) := X"0062102B";
        ram_buffer(67119) := X"1440000A";
        ram_buffer(67120) := X"00000000";
        ram_buffer(67121) := X"8EC200CC";
        ram_buffer(67122) := X"2403FFFF";
        ram_buffer(67123) := X"8C420000";
        ram_buffer(67124) := X"00000000";
        ram_buffer(67125) := X"10430010";
        ram_buffer(67126) := X"00402821";
        ram_buffer(67127) := X"0C02FD29";
        ram_buffer(67128) := X"00000000";
        ram_buffer(67129) := X"8EC30044";
        ram_buffer(67130) := X"8EC200CC";
        ram_buffer(67131) := X"24640001";
        ram_buffer(67132) := X"AEC40044";
        ram_buffer(67133) := X"00431821";
        ram_buffer(67134) := X"90620004";
        ram_buffer(67135) := X"27DE0001";
        ram_buffer(67136) := X"A2A20000";
        ram_buffer(67137) := X"8EC20048";
        ram_buffer(67138) := X"26B50001";
        ram_buffer(67139) := X"24420001";
        ram_buffer(67140) := X"17D4FFDD";
        ram_buffer(67141) := X"AEC20048";
        ram_buffer(67142) := X"8FA40018";
        ram_buffer(67143) := X"AFB00010";
        ram_buffer(67144) := X"03C03821";
        ram_buffer(67145) := X"02E03021";
        ram_buffer(67146) := X"0C028116";
        ram_buffer(67147) := X"02202821";
        ram_buffer(67148) := X"0C03013B";
        ram_buffer(67149) := X"02C02021";
        ram_buffer(67150) := X"26F70001";
        ram_buffer(67151) := X"24020005";
        ram_buffer(67152) := X"16E2FFC3";
        ram_buffer(67153) := X"02203821";
        ram_buffer(67154) := X"26310001";
        ram_buffer(67155) := X"1637FFBF";
        ram_buffer(67156) := X"0000B821";
        ram_buffer(67157) := X"8FA20024";
        ram_buffer(67158) := X"00009021";
        ram_buffer(67159) := X"0C0301F5";
        ram_buffer(67160) := X"2444B4FC";
        ram_buffer(67161) := X"8FA2003C";
        ram_buffer(67162) := X"24140005";
        ram_buffer(67163) := X"0C0301F5";
        ram_buffer(67164) := X"2444B4EC";
        ram_buffer(67165) := X"3C04100D";
        ram_buffer(67166) := X"0C0301F5";
        ram_buffer(67167) := X"2484B588";
        ram_buffer(67168) := X"8FA2002C";
        ram_buffer(67169) := X"00000000";
        ram_buffer(67170) := X"2453B524";
        ram_buffer(67171) := X"8FA20028";
        ram_buffer(67172) := X"00000000";
        ram_buffer(67173) := X"2455B51C";
        ram_buffer(67174) := X"00008821";
        ram_buffer(67175) := X"AFB10010";
        ram_buffer(67176) := X"02002021";
        ram_buffer(67177) := X"02403821";
        ram_buffer(67178) := X"02403021";
        ram_buffer(67179) := X"0C0283DB";
        ram_buffer(67180) := X"02602821";
        ram_buffer(67181) := X"26310001";
        ram_buffer(67182) := X"0C0301F5";
        ram_buffer(67183) := X"02002021";
        ram_buffer(67184) := X"1634FFF6";
        ram_buffer(67185) := X"02403021";
        ram_buffer(67186) := X"02002021";
        ram_buffer(67187) := X"0C0283DB";
        ram_buffer(67188) := X"02A02821";
        ram_buffer(67189) := X"26520001";
        ram_buffer(67190) := X"0C0301F5";
        ram_buffer(67191) := X"02002021";
        ram_buffer(67192) := X"1651FFEE";
        ram_buffer(67193) := X"00008821";
        ram_buffer(67194) := X"8FA20030";
        ram_buffer(67195) := X"0C03044C";
        ram_buffer(67196) := X"2444B3F0";
        ram_buffer(67197) := X"0C027A4D";
        ram_buffer(67198) := X"02002021";
        ram_buffer(67199) := X"00001021";
        ram_buffer(67200) := X"8FBF0064";
        ram_buffer(67201) := X"8FBE0060";
        ram_buffer(67202) := X"8FB7005C";
        ram_buffer(67203) := X"8FB60058";
        ram_buffer(67204) := X"8FB50054";
        ram_buffer(67205) := X"8FB40050";
        ram_buffer(67206) := X"8FB3004C";
        ram_buffer(67207) := X"8FB20048";
        ram_buffer(67208) := X"8FB10044";
        ram_buffer(67209) := X"8FB00040";
        ram_buffer(67210) := X"03E00008";
        ram_buffer(67211) := X"27BD0068";
        ram_buffer(67212) := X"1000FFF3";
        ram_buffer(67213) := X"2402FFFF";
        ram_buffer(67214) := X"8F8281E8";
        ram_buffer(67215) := X"00000000";
        ram_buffer(67216) := X"10400003";
        ram_buffer(67217) := X"00000000";
        ram_buffer(67218) := X"08027F93";
        ram_buffer(67219) := X"00452821";
        ram_buffer(67220) := X"3C021000";
        ram_buffer(67221) := X"00452821";
        ram_buffer(67222) := X"08027F93";
        ram_buffer(67223) := X"AF8281E8";
        ram_buffer(67224) := X"8F8281E8";
        ram_buffer(67225) := X"00000000";
        ram_buffer(67226) := X"00451021";
        ram_buffer(67227) := X"00802821";
        ram_buffer(67228) := X"08027F93";
        ram_buffer(67229) := X"00402021";
        ram_buffer(67230) := X"8F8281E8";
        ram_buffer(67231) := X"24060200";
        ram_buffer(67232) := X"240500FF";
        ram_buffer(67233) := X"0802801D";
        ram_buffer(67234) := X"00442021";
        ram_buffer(67235) := X"27BDFFE0";
        ram_buffer(67236) := X"AFB10018";
        ram_buffer(67237) := X"AFB00014";
        ram_buffer(67238) := X"AFBF001C";
        ram_buffer(67239) := X"00008021";
        ram_buffer(67240) := X"3C110008";
        ram_buffer(67241) := X"8F8281E8";
        ram_buffer(67242) := X"00000000";
        ram_buffer(67243) := X"00501021";
        ram_buffer(67244) := X"90440000";
        ram_buffer(67245) := X"0C0306B6";
        ram_buffer(67246) := X"26100001";
        ram_buffer(67247) := X"1611FFF9";
        ram_buffer(67248) := X"00000000";
        ram_buffer(67249) := X"8FBF001C";
        ram_buffer(67250) := X"8FB10018";
        ram_buffer(67251) := X"8FB00014";
        ram_buffer(67252) := X"03E00008";
        ram_buffer(67253) := X"27BD0020";
        ram_buffer(67254) := X"3C032000";
        ram_buffer(67255) := X"8C620020";
        ram_buffer(67256) := X"00000000";
        ram_buffer(67257) := X"30420002";
        ram_buffer(67258) := X"1040FFFB";
        ram_buffer(67259) := X"00000000";
        ram_buffer(67260) := X"AC640000";
        ram_buffer(67261) := X"03E00008";
        ram_buffer(67262) := X"00001021";
        ram_buffer(67263) := X"80820000";
        ram_buffer(67264) := X"00000000";
        ram_buffer(67265) := X"10400010";
        ram_buffer(67266) := X"2406000A";
        ram_buffer(67267) := X"2407000D";
        ram_buffer(67268) := X"1046000F";
        ram_buffer(67269) := X"00402821";
        ram_buffer(67270) := X"24840001";
        ram_buffer(67271) := X"3C032000";
        ram_buffer(67272) := X"8C620020";
        ram_buffer(67273) := X"00000000";
        ram_buffer(67274) := X"30420002";
        ram_buffer(67275) := X"1040FFFB";
        ram_buffer(67276) := X"00000000";
        ram_buffer(67277) := X"AC650000";
        ram_buffer(67278) := X"80820000";
        ram_buffer(67279) := X"00000000";
        ram_buffer(67280) := X"1440FFF3";
        ram_buffer(67281) := X"00000000";
        ram_buffer(67282) := X"03E00008";
        ram_buffer(67283) := X"00001021";
        ram_buffer(67284) := X"3C032000";
        ram_buffer(67285) := X"8C620020";
        ram_buffer(67286) := X"00000000";
        ram_buffer(67287) := X"30420002";
        ram_buffer(67288) := X"1040FFFB";
        ram_buffer(67289) := X"00000000";
        ram_buffer(67290) := X"AC670000";
        ram_buffer(67291) := X"80850000";
        ram_buffer(67292) := X"1000FFEA";
        ram_buffer(67293) := X"24840001";
        ram_buffer(67294) := X"2406001C";
        ram_buffer(67295) := X"2407FFFC";
        ram_buffer(67296) := X"00C41006";
        ram_buffer(67297) := X"3042000F";
        ram_buffer(67298) := X"2C43000A";
        ram_buffer(67299) := X"1060000E";
        ram_buffer(67300) := X"24450057";
        ram_buffer(67301) := X"24450030";
        ram_buffer(67302) := X"3C032000";
        ram_buffer(67303) := X"8C620020";
        ram_buffer(67304) := X"00000000";
        ram_buffer(67305) := X"30420002";
        ram_buffer(67306) := X"1040FFFB";
        ram_buffer(67307) := X"00000000";
        ram_buffer(67308) := X"24C6FFFC";
        ram_buffer(67309) := X"AC650000";
        ram_buffer(67310) := X"14C7FFF2";
        ram_buffer(67311) := X"00C41006";
        ram_buffer(67312) := X"03E00008";
        ram_buffer(67313) := X"00000000";
        ram_buffer(67314) := X"3C032000";
        ram_buffer(67315) := X"8C620020";
        ram_buffer(67316) := X"00000000";
        ram_buffer(67317) := X"30420002";
        ram_buffer(67318) := X"1040FFFB";
        ram_buffer(67319) := X"00000000";
        ram_buffer(67320) := X"24C6FFFC";
        ram_buffer(67321) := X"AC650000";
        ram_buffer(67322) := X"14C7FFE6";
        ram_buffer(67323) := X"00C41006";
        ram_buffer(67324) := X"1000FFF3";
        ram_buffer(67325) := X"00000000";
        ram_buffer(67326) := X"3C022000";
        ram_buffer(67327) := X"8C420020";
        ram_buffer(67328) := X"03E00008";
        ram_buffer(67329) := X"30420001";
        ram_buffer(67330) := X"3C032000";
        ram_buffer(67331) := X"8C620020";
        ram_buffer(67332) := X"00000000";
        ram_buffer(67333) := X"30420001";
        ram_buffer(67334) := X"1040FFFB";
        ram_buffer(67335) := X"00000000";
        ram_buffer(67336) := X"8C620000";
        ram_buffer(67337) := X"03E00008";
        ram_buffer(67338) := X"00000000";
        ram_buffer(67339) := X"3C022000";
        ram_buffer(67340) := X"8C430068";
        ram_buffer(67341) := X"8C420060";
        ram_buffer(67342) := X"03E00008";
        ram_buffer(67343) := X"00000000";
        ram_buffer(67344) := X"3C04100D";
        ram_buffer(67345) := X"27BDFFE8";
        ram_buffer(67346) := X"AFBF0014";
        ram_buffer(67347) := X"0C0306BF";
        ram_buffer(67348) := X"2484B590";
        ram_buffer(67349) := X"3C032000";
        ram_buffer(67350) := X"8C620020";
        ram_buffer(67351) := X"00000000";
        ram_buffer(67352) := X"30420002";
        ram_buffer(67353) := X"1040FFFC";
        ram_buffer(67354) := X"2402000A";
        ram_buffer(67355) := X"AC620000";
        ram_buffer(67356) := X"1000FFFF";
        ram_buffer(67357) := X"00000000";
        ram_buffer(67358) := X"27BDFFE8";
        ram_buffer(67359) := X"AFBF0014";
        ram_buffer(67360) := X"AFBE0010";
        ram_buffer(67361) := X"03A0F021";
        ram_buffer(67362) := X"AFC40018";
        ram_buffer(67363) := X"AFC5001C";
        ram_buffer(67364) := X"8F828098";
        ram_buffer(67365) := X"8FC6001C";
        ram_buffer(67366) := X"8FC50018";
        ram_buffer(67367) := X"00402021";
        ram_buffer(67368) := X"0C02F251";
        ram_buffer(67369) := X"00000000";
        ram_buffer(67370) := X"03C0E821";
        ram_buffer(67371) := X"8FBF0014";
        ram_buffer(67372) := X"8FBE0010";
        ram_buffer(67373) := X"27BD0018";
        ram_buffer(67374) := X"03E00008";
        ram_buffer(67375) := X"00000000";
        ram_buffer(67376) := X"27BDFFF8";
        ram_buffer(67377) := X"AFBE0004";
        ram_buffer(67378) := X"03A0F021";
        ram_buffer(67379) := X"8F828098";
        ram_buffer(67380) := X"03C0E821";
        ram_buffer(67381) := X"8FBE0004";
        ram_buffer(67382) := X"27BD0008";
        ram_buffer(67383) := X"03E00008";
        ram_buffer(67384) := X"00000000";
        ram_buffer(67385) := X"27BDFFE0";
        ram_buffer(67386) := X"AFBF001C";
        ram_buffer(67387) := X"AFBE0018";
        ram_buffer(67388) := X"03A0F021";
        ram_buffer(67389) := X"AFC40020";
        ram_buffer(67390) := X"00A01021";
        ram_buffer(67391) := X"00402821";
        ram_buffer(67392) := X"8FC40020";
        ram_buffer(67393) := X"0C03075B";
        ram_buffer(67394) := X"00000000";
        ram_buffer(67395) := X"AFC20010";
        ram_buffer(67396) := X"8FC20010";
        ram_buffer(67397) := X"03C0E821";
        ram_buffer(67398) := X"8FBF001C";
        ram_buffer(67399) := X"8FBE0018";
        ram_buffer(67400) := X"27BD0020";
        ram_buffer(67401) := X"03E00008";
        ram_buffer(67402) := X"00000000";
        ram_buffer(67403) := X"27BDFFE8";
        ram_buffer(67404) := X"AFBF0014";
        ram_buffer(67405) := X"AFBE0010";
        ram_buffer(67406) := X"03A0F021";
        ram_buffer(67407) := X"00801821";
        ram_buffer(67408) := X"8F828098";
        ram_buffer(67409) := X"00602821";
        ram_buffer(67410) := X"00402021";
        ram_buffer(67411) := X"0C030739";
        ram_buffer(67412) := X"00000000";
        ram_buffer(67413) := X"03C0E821";
        ram_buffer(67414) := X"8FBF0014";
        ram_buffer(67415) := X"8FBE0010";
        ram_buffer(67416) := X"27BD0018";
        ram_buffer(67417) := X"03E00008";
        ram_buffer(67418) := X"00000000";
        ram_buffer(67419) := X"27BDFFD8";
        ram_buffer(67420) := X"AFBF0024";
        ram_buffer(67421) := X"AFBE0020";
        ram_buffer(67422) := X"AFB0001C";
        ram_buffer(67423) := X"03A0F021";
        ram_buffer(67424) := X"AFC40028";
        ram_buffer(67425) := X"00A08021";
        ram_buffer(67426) := X"8FC20028";
        ram_buffer(67427) := X"00000000";
        ram_buffer(67428) := X"AFC20014";
        ram_buffer(67429) := X"8FC20014";
        ram_buffer(67430) := X"00000000";
        ram_buffer(67431) := X"1040000A";
        ram_buffer(67432) := X"00000000";
        ram_buffer(67433) := X"8FC20014";
        ram_buffer(67434) := X"00000000";
        ram_buffer(67435) := X"8C420038";
        ram_buffer(67436) := X"00000000";
        ram_buffer(67437) := X"14400004";
        ram_buffer(67438) := X"00000000";
        ram_buffer(67439) := X"8FC40014";
        ram_buffer(67440) := X"0C027069";
        ram_buffer(67441) := X"00000000";
        ram_buffer(67442) := X"8E020028";
        ram_buffer(67443) := X"00000000";
        ram_buffer(67444) := X"14400007";
        ram_buffer(67445) := X"00000000";
        ram_buffer(67446) := X"8FC20028";
        ram_buffer(67447) := X"2403001D";
        ram_buffer(67448) := X"AC430000";
        ram_buffer(67449) := X"2402FFFF";
        ram_buffer(67450) := X"10000051";
        ram_buffer(67451) := X"00000000";
        ram_buffer(67452) := X"8602000C";
        ram_buffer(67453) := X"00000000";
        ram_buffer(67454) := X"3042FFFF";
        ram_buffer(67455) := X"30420008";
        ram_buffer(67456) := X"10400005";
        ram_buffer(67457) := X"00000000";
        ram_buffer(67458) := X"02002821";
        ram_buffer(67459) := X"8FC40028";
        ram_buffer(67460) := X"0C026EE1";
        ram_buffer(67461) := X"00000000";
        ram_buffer(67462) := X"8602000C";
        ram_buffer(67463) := X"00000000";
        ram_buffer(67464) := X"3042FFFF";
        ram_buffer(67465) := X"30421000";
        ram_buffer(67466) := X"10400006";
        ram_buffer(67467) := X"00000000";
        ram_buffer(67468) := X"8E020050";
        ram_buffer(67469) := X"00000000";
        ram_buffer(67470) := X"AFC20010";
        ram_buffer(67471) := X"10000011";
        ram_buffer(67472) := X"00000000";
        ram_buffer(67473) := X"8E020028";
        ram_buffer(67474) := X"8E03001C";
        ram_buffer(67475) := X"24070001";
        ram_buffer(67476) := X"00003021";
        ram_buffer(67477) := X"00602821";
        ram_buffer(67478) := X"8FC40028";
        ram_buffer(67479) := X"0040F809";
        ram_buffer(67480) := X"00000000";
        ram_buffer(67481) := X"AFC20010";
        ram_buffer(67482) := X"8FC30010";
        ram_buffer(67483) := X"2402FFFF";
        ram_buffer(67484) := X"14620004";
        ram_buffer(67485) := X"00000000";
        ram_buffer(67486) := X"8FC20010";
        ram_buffer(67487) := X"1000002C";
        ram_buffer(67488) := X"00000000";
        ram_buffer(67489) := X"8602000C";
        ram_buffer(67490) := X"00000000";
        ram_buffer(67491) := X"3042FFFF";
        ram_buffer(67492) := X"30420004";
        ram_buffer(67493) := X"10400011";
        ram_buffer(67494) := X"00000000";
        ram_buffer(67495) := X"8E020004";
        ram_buffer(67496) := X"8FC30010";
        ram_buffer(67497) := X"00000000";
        ram_buffer(67498) := X"00621023";
        ram_buffer(67499) := X"AFC20010";
        ram_buffer(67500) := X"8E020030";
        ram_buffer(67501) := X"00000000";
        ram_buffer(67502) := X"1040001C";
        ram_buffer(67503) := X"00000000";
        ram_buffer(67504) := X"8E02003C";
        ram_buffer(67505) := X"8FC30010";
        ram_buffer(67506) := X"00000000";
        ram_buffer(67507) := X"00621023";
        ram_buffer(67508) := X"AFC20010";
        ram_buffer(67509) := X"10000015";
        ram_buffer(67510) := X"00000000";
        ram_buffer(67511) := X"8602000C";
        ram_buffer(67512) := X"00000000";
        ram_buffer(67513) := X"3042FFFF";
        ram_buffer(67514) := X"30420008";
        ram_buffer(67515) := X"1040000F";
        ram_buffer(67516) := X"00000000";
        ram_buffer(67517) := X"8E020000";
        ram_buffer(67518) := X"00000000";
        ram_buffer(67519) := X"1040000B";
        ram_buffer(67520) := X"00000000";
        ram_buffer(67521) := X"8E020000";
        ram_buffer(67522) := X"00000000";
        ram_buffer(67523) := X"00401821";
        ram_buffer(67524) := X"8E020010";
        ram_buffer(67525) := X"00000000";
        ram_buffer(67526) := X"00621023";
        ram_buffer(67527) := X"8FC30010";
        ram_buffer(67528) := X"00000000";
        ram_buffer(67529) := X"00621021";
        ram_buffer(67530) := X"AFC20010";
        ram_buffer(67531) := X"8FC20010";
        ram_buffer(67532) := X"03C0E821";
        ram_buffer(67533) := X"8FBF0024";
        ram_buffer(67534) := X"8FBE0020";
        ram_buffer(67535) := X"8FB0001C";
        ram_buffer(67536) := X"27BD0028";
        ram_buffer(67537) := X"03E00008";
        ram_buffer(67538) := X"00000000";
        ram_buffer(67539) := X"27BDFFE8";
        ram_buffer(67540) := X"AFBF0014";
        ram_buffer(67541) := X"AFBE0010";
        ram_buffer(67542) := X"03A0F021";
        ram_buffer(67543) := X"00801821";
        ram_buffer(67544) := X"8F828098";
        ram_buffer(67545) := X"00602821";
        ram_buffer(67546) := X"00402021";
        ram_buffer(67547) := X"0C03075B";
        ram_buffer(67548) := X"00000000";
        ram_buffer(67549) := X"03C0E821";
        ram_buffer(67550) := X"8FBF0014";
        ram_buffer(67551) := X"8FBE0010";
        ram_buffer(67552) := X"27BD0018";
        ram_buffer(67553) := X"03E00008";
        ram_buffer(67554) := X"00000000";
        ram_buffer(67555) := X"27BDFFE8";
        ram_buffer(67556) := X"AFBE0014";
        ram_buffer(67557) := X"03A0F021";
        ram_buffer(67558) := X"AFC40018";
        ram_buffer(67559) := X"AFC5001C";
        ram_buffer(67560) := X"AFC60020";
        ram_buffer(67561) := X"8FC20018";
        ram_buffer(67562) := X"00000000";
        ram_buffer(67563) := X"AFC20000";
        ram_buffer(67564) := X"8FC2001C";
        ram_buffer(67565) := X"00000000";
        ram_buffer(67566) := X"AFC20004";
        ram_buffer(67567) := X"8FC20020";
        ram_buffer(67568) := X"00000000";
        ram_buffer(67569) := X"2C420004";
        ram_buffer(67570) := X"14400052";
        ram_buffer(67571) := X"00000000";
        ram_buffer(67572) := X"8FC30000";
        ram_buffer(67573) := X"8FC20004";
        ram_buffer(67574) := X"00000000";
        ram_buffer(67575) := X"00621025";
        ram_buffer(67576) := X"30420003";
        ram_buffer(67577) := X"1440004B";
        ram_buffer(67578) := X"00000000";
        ram_buffer(67579) := X"8FC20000";
        ram_buffer(67580) := X"00000000";
        ram_buffer(67581) := X"AFC20008";
        ram_buffer(67582) := X"8FC20004";
        ram_buffer(67583) := X"00000000";
        ram_buffer(67584) := X"AFC2000C";
        ram_buffer(67585) := X"10000016";
        ram_buffer(67586) := X"00000000";
        ram_buffer(67587) := X"8FC20008";
        ram_buffer(67588) := X"00000000";
        ram_buffer(67589) := X"8C430000";
        ram_buffer(67590) := X"8FC2000C";
        ram_buffer(67591) := X"00000000";
        ram_buffer(67592) := X"8C420000";
        ram_buffer(67593) := X"00000000";
        ram_buffer(67594) := X"14620014";
        ram_buffer(67595) := X"00000000";
        ram_buffer(67596) := X"8FC20008";
        ram_buffer(67597) := X"00000000";
        ram_buffer(67598) := X"24420004";
        ram_buffer(67599) := X"AFC20008";
        ram_buffer(67600) := X"8FC2000C";
        ram_buffer(67601) := X"00000000";
        ram_buffer(67602) := X"24420004";
        ram_buffer(67603) := X"AFC2000C";
        ram_buffer(67604) := X"8FC20020";
        ram_buffer(67605) := X"00000000";
        ram_buffer(67606) := X"2442FFFC";
        ram_buffer(67607) := X"AFC20020";
        ram_buffer(67608) := X"8FC20020";
        ram_buffer(67609) := X"00000000";
        ram_buffer(67610) := X"2C420004";
        ram_buffer(67611) := X"1040FFE7";
        ram_buffer(67612) := X"00000000";
        ram_buffer(67613) := X"10000002";
        ram_buffer(67614) := X"00000000";
        ram_buffer(67615) := X"00000000";
        ram_buffer(67616) := X"8FC20008";
        ram_buffer(67617) := X"00000000";
        ram_buffer(67618) := X"AFC20000";
        ram_buffer(67619) := X"8FC2000C";
        ram_buffer(67620) := X"00000000";
        ram_buffer(67621) := X"AFC20004";
        ram_buffer(67622) := X"1000001E";
        ram_buffer(67623) := X"00000000";
        ram_buffer(67624) := X"8FC20000";
        ram_buffer(67625) := X"00000000";
        ram_buffer(67626) := X"90430000";
        ram_buffer(67627) := X"8FC20004";
        ram_buffer(67628) := X"00000000";
        ram_buffer(67629) := X"90420000";
        ram_buffer(67630) := X"00000000";
        ram_buffer(67631) := X"1062000D";
        ram_buffer(67632) := X"00000000";
        ram_buffer(67633) := X"8FC20000";
        ram_buffer(67634) := X"00000000";
        ram_buffer(67635) := X"90420000";
        ram_buffer(67636) := X"00000000";
        ram_buffer(67637) := X"00401821";
        ram_buffer(67638) := X"8FC20004";
        ram_buffer(67639) := X"00000000";
        ram_buffer(67640) := X"90420000";
        ram_buffer(67641) := X"00000000";
        ram_buffer(67642) := X"00621023";
        ram_buffer(67643) := X"10000010";
        ram_buffer(67644) := X"00000000";
        ram_buffer(67645) := X"8FC20000";
        ram_buffer(67646) := X"00000000";
        ram_buffer(67647) := X"24420001";
        ram_buffer(67648) := X"AFC20000";
        ram_buffer(67649) := X"8FC20004";
        ram_buffer(67650) := X"00000000";
        ram_buffer(67651) := X"24420001";
        ram_buffer(67652) := X"AFC20004";
        ram_buffer(67653) := X"8FC20020";
        ram_buffer(67654) := X"00000000";
        ram_buffer(67655) := X"2443FFFF";
        ram_buffer(67656) := X"AFC30020";
        ram_buffer(67657) := X"1440FFDE";
        ram_buffer(67658) := X"00000000";
        ram_buffer(67659) := X"00001021";
        ram_buffer(67660) := X"03C0E821";
        ram_buffer(67661) := X"8FBE0014";
        ram_buffer(67662) := X"27BD0018";
        ram_buffer(67663) := X"03E00008";
        ram_buffer(67664) := X"00000000";
        ram_buffer(67665) := X"27BDFFE8";
        ram_buffer(67666) := X"AFBF0014";
        ram_buffer(67667) := X"AFBE0010";
        ram_buffer(67668) := X"03A0F021";
        ram_buffer(67669) := X"AFC40018";
        ram_buffer(67670) := X"AFC5001C";
        ram_buffer(67671) := X"8FC20018";
        ram_buffer(67672) := X"00000000";
        ram_buffer(67673) := X"8C420008";
        ram_buffer(67674) := X"00000000";
        ram_buffer(67675) := X"00403021";
        ram_buffer(67676) := X"8FC5001C";
        ram_buffer(67677) := X"8FC40018";
        ram_buffer(67678) := X"0C0309B1";
        ram_buffer(67679) := X"00000000";
        ram_buffer(67680) := X"03C0E821";
        ram_buffer(67681) := X"8FBF0014";
        ram_buffer(67682) := X"8FBE0010";
        ram_buffer(67683) := X"27BD0018";
        ram_buffer(67684) := X"03E00008";
        ram_buffer(67685) := X"00000000";
        ram_buffer(67686) := X"27BDFFE0";
        ram_buffer(67687) := X"AFBF001C";
        ram_buffer(67688) := X"AFBE0018";
        ram_buffer(67689) := X"03A0F021";
        ram_buffer(67690) := X"AFC40020";
        ram_buffer(67691) := X"8F828098";
        ram_buffer(67692) := X"00000000";
        ram_buffer(67693) := X"AFC20010";
        ram_buffer(67694) := X"8FC20010";
        ram_buffer(67695) := X"00000000";
        ram_buffer(67696) := X"8C420008";
        ram_buffer(67697) := X"00000000";
        ram_buffer(67698) := X"00403021";
        ram_buffer(67699) := X"8FC50020";
        ram_buffer(67700) := X"8FC40010";
        ram_buffer(67701) := X"0C0309B1";
        ram_buffer(67702) := X"00000000";
        ram_buffer(67703) := X"03C0E821";
        ram_buffer(67704) := X"8FBF001C";
        ram_buffer(67705) := X"8FBE0018";
        ram_buffer(67706) := X"27BD0020";
        ram_buffer(67707) := X"03E00008";
        ram_buffer(67708) := X"00000000";
        ram_buffer(67709) := X"27BDFFE0";
        ram_buffer(67710) := X"AFBE001C";
        ram_buffer(67711) := X"03A0F021";
        ram_buffer(67712) := X"AFC40020";
        ram_buffer(67713) := X"AFC50024";
        ram_buffer(67714) := X"8FC20020";
        ram_buffer(67715) := X"00000000";
        ram_buffer(67716) := X"AFC20000";
        ram_buffer(67717) := X"8FC20024";
        ram_buffer(67718) := X"00000000";
        ram_buffer(67719) := X"A3C20010";
        ram_buffer(67720) := X"93C20010";
        ram_buffer(67721) := X"00000000";
        ram_buffer(67722) := X"14400058";
        ram_buffer(67723) := X"00000000";
        ram_buffer(67724) := X"1000000E";
        ram_buffer(67725) := X"00000000";
        ram_buffer(67726) := X"8FC20000";
        ram_buffer(67727) := X"00000000";
        ram_buffer(67728) := X"90420000";
        ram_buffer(67729) := X"00000000";
        ram_buffer(67730) := X"14400004";
        ram_buffer(67731) := X"00000000";
        ram_buffer(67732) := X"8FC20000";
        ram_buffer(67733) := X"100000BB";
        ram_buffer(67734) := X"00000000";
        ram_buffer(67735) := X"8FC20000";
        ram_buffer(67736) := X"00000000";
        ram_buffer(67737) := X"24420001";
        ram_buffer(67738) := X"AFC20000";
        ram_buffer(67739) := X"8FC20000";
        ram_buffer(67740) := X"00000000";
        ram_buffer(67741) := X"30420003";
        ram_buffer(67742) := X"1440FFEF";
        ram_buffer(67743) := X"00000000";
        ram_buffer(67744) := X"8FC20000";
        ram_buffer(67745) := X"00000000";
        ram_buffer(67746) := X"AFC2000C";
        ram_buffer(67747) := X"10000005";
        ram_buffer(67748) := X"00000000";
        ram_buffer(67749) := X"8FC2000C";
        ram_buffer(67750) := X"00000000";
        ram_buffer(67751) := X"24420004";
        ram_buffer(67752) := X"AFC2000C";
        ram_buffer(67753) := X"8FC2000C";
        ram_buffer(67754) := X"00000000";
        ram_buffer(67755) := X"8C430000";
        ram_buffer(67756) := X"3C02FEFE";
        ram_buffer(67757) := X"3442FEFF";
        ram_buffer(67758) := X"00621821";
        ram_buffer(67759) := X"8FC2000C";
        ram_buffer(67760) := X"00000000";
        ram_buffer(67761) := X"8C420000";
        ram_buffer(67762) := X"00000000";
        ram_buffer(67763) := X"00021027";
        ram_buffer(67764) := X"00621824";
        ram_buffer(67765) := X"3C028080";
        ram_buffer(67766) := X"34428080";
        ram_buffer(67767) := X"00621024";
        ram_buffer(67768) := X"1040FFEC";
        ram_buffer(67769) := X"00000000";
        ram_buffer(67770) := X"8FC2000C";
        ram_buffer(67771) := X"00000000";
        ram_buffer(67772) := X"AFC20000";
        ram_buffer(67773) := X"10000005";
        ram_buffer(67774) := X"00000000";
        ram_buffer(67775) := X"8FC20000";
        ram_buffer(67776) := X"00000000";
        ram_buffer(67777) := X"24420001";
        ram_buffer(67778) := X"AFC20000";
        ram_buffer(67779) := X"8FC20000";
        ram_buffer(67780) := X"00000000";
        ram_buffer(67781) := X"90420000";
        ram_buffer(67782) := X"00000000";
        ram_buffer(67783) := X"1440FFF7";
        ram_buffer(67784) := X"00000000";
        ram_buffer(67785) := X"8FC20000";
        ram_buffer(67786) := X"10000086";
        ram_buffer(67787) := X"00000000";
        ram_buffer(67788) := X"8FC20000";
        ram_buffer(67789) := X"00000000";
        ram_buffer(67790) := X"90420000";
        ram_buffer(67791) := X"00000000";
        ram_buffer(67792) := X"14400004";
        ram_buffer(67793) := X"00000000";
        ram_buffer(67794) := X"00001021";
        ram_buffer(67795) := X"1000007D";
        ram_buffer(67796) := X"00000000";
        ram_buffer(67797) := X"8FC20000";
        ram_buffer(67798) := X"00000000";
        ram_buffer(67799) := X"90420000";
        ram_buffer(67800) := X"93C30010";
        ram_buffer(67801) := X"00000000";
        ram_buffer(67802) := X"14620004";
        ram_buffer(67803) := X"00000000";
        ram_buffer(67804) := X"8FC20000";
        ram_buffer(67805) := X"10000073";
        ram_buffer(67806) := X"00000000";
        ram_buffer(67807) := X"8FC20000";
        ram_buffer(67808) := X"00000000";
        ram_buffer(67809) := X"24420001";
        ram_buffer(67810) := X"AFC20000";
        ram_buffer(67811) := X"8FC20000";
        ram_buffer(67812) := X"00000000";
        ram_buffer(67813) := X"30420003";
        ram_buffer(67814) := X"1440FFE5";
        ram_buffer(67815) := X"00000000";
        ram_buffer(67816) := X"93C20010";
        ram_buffer(67817) := X"00000000";
        ram_buffer(67818) := X"AFC20004";
        ram_buffer(67819) := X"24020008";
        ram_buffer(67820) := X"AFC20008";
        ram_buffer(67821) := X"1000000D";
        ram_buffer(67822) := X"00000000";
        ram_buffer(67823) := X"8FC30004";
        ram_buffer(67824) := X"8FC20008";
        ram_buffer(67825) := X"00000000";
        ram_buffer(67826) := X"00431004";
        ram_buffer(67827) := X"8FC30004";
        ram_buffer(67828) := X"00000000";
        ram_buffer(67829) := X"00621025";
        ram_buffer(67830) := X"AFC20004";
        ram_buffer(67831) := X"8FC20008";
        ram_buffer(67832) := X"00000000";
        ram_buffer(67833) := X"00021040";
        ram_buffer(67834) := X"AFC20008";
        ram_buffer(67835) := X"8FC20008";
        ram_buffer(67836) := X"00000000";
        ram_buffer(67837) := X"2C420020";
        ram_buffer(67838) := X"1440FFF0";
        ram_buffer(67839) := X"00000000";
        ram_buffer(67840) := X"8FC20000";
        ram_buffer(67841) := X"00000000";
        ram_buffer(67842) := X"AFC2000C";
        ram_buffer(67843) := X"10000005";
        ram_buffer(67844) := X"00000000";
        ram_buffer(67845) := X"8FC2000C";
        ram_buffer(67846) := X"00000000";
        ram_buffer(67847) := X"24420004";
        ram_buffer(67848) := X"AFC2000C";
        ram_buffer(67849) := X"8FC2000C";
        ram_buffer(67850) := X"00000000";
        ram_buffer(67851) := X"8C430000";
        ram_buffer(67852) := X"3C02FEFE";
        ram_buffer(67853) := X"3442FEFF";
        ram_buffer(67854) := X"00621821";
        ram_buffer(67855) := X"8FC2000C";
        ram_buffer(67856) := X"00000000";
        ram_buffer(67857) := X"8C420000";
        ram_buffer(67858) := X"00000000";
        ram_buffer(67859) := X"00021027";
        ram_buffer(67860) := X"00621824";
        ram_buffer(67861) := X"3C028080";
        ram_buffer(67862) := X"34428080";
        ram_buffer(67863) := X"00621024";
        ram_buffer(67864) := X"14400017";
        ram_buffer(67865) := X"00000000";
        ram_buffer(67866) := X"8FC2000C";
        ram_buffer(67867) := X"00000000";
        ram_buffer(67868) := X"8C430000";
        ram_buffer(67869) := X"8FC20004";
        ram_buffer(67870) := X"00000000";
        ram_buffer(67871) := X"00621826";
        ram_buffer(67872) := X"3C02FEFE";
        ram_buffer(67873) := X"3442FEFF";
        ram_buffer(67874) := X"00621821";
        ram_buffer(67875) := X"8FC2000C";
        ram_buffer(67876) := X"00000000";
        ram_buffer(67877) := X"8C440000";
        ram_buffer(67878) := X"8FC20004";
        ram_buffer(67879) := X"00000000";
        ram_buffer(67880) := X"00821026";
        ram_buffer(67881) := X"00021027";
        ram_buffer(67882) := X"00621824";
        ram_buffer(67883) := X"3C028080";
        ram_buffer(67884) := X"34428080";
        ram_buffer(67885) := X"00621024";
        ram_buffer(67886) := X"1040FFD6";
        ram_buffer(67887) := X"00000000";
        ram_buffer(67888) := X"8FC2000C";
        ram_buffer(67889) := X"00000000";
        ram_buffer(67890) := X"AFC20000";
        ram_buffer(67891) := X"10000005";
        ram_buffer(67892) := X"00000000";
        ram_buffer(67893) := X"8FC20000";
        ram_buffer(67894) := X"00000000";
        ram_buffer(67895) := X"24420001";
        ram_buffer(67896) := X"AFC20000";
        ram_buffer(67897) := X"8FC20000";
        ram_buffer(67898) := X"00000000";
        ram_buffer(67899) := X"90420000";
        ram_buffer(67900) := X"00000000";
        ram_buffer(67901) := X"10400008";
        ram_buffer(67902) := X"00000000";
        ram_buffer(67903) := X"8FC20000";
        ram_buffer(67904) := X"00000000";
        ram_buffer(67905) := X"90420000";
        ram_buffer(67906) := X"93C30010";
        ram_buffer(67907) := X"00000000";
        ram_buffer(67908) := X"1462FFF0";
        ram_buffer(67909) := X"00000000";
        ram_buffer(67910) := X"8FC20000";
        ram_buffer(67911) := X"00000000";
        ram_buffer(67912) := X"90420000";
        ram_buffer(67913) := X"93C30010";
        ram_buffer(67914) := X"00000000";
        ram_buffer(67915) := X"14620004";
        ram_buffer(67916) := X"00000000";
        ram_buffer(67917) := X"8FC20000";
        ram_buffer(67918) := X"10000002";
        ram_buffer(67919) := X"00000000";
        ram_buffer(67920) := X"00001021";
        ram_buffer(67921) := X"03C0E821";
        ram_buffer(67922) := X"8FBE001C";
        ram_buffer(67923) := X"27BD0020";
        ram_buffer(67924) := X"03E00008";
        ram_buffer(67925) := X"00000000";
        ram_buffer(67926) := X"27BDFFF0";
        ram_buffer(67927) := X"AFBE000C";
        ram_buffer(67928) := X"03A0F021";
        ram_buffer(67929) := X"AFC40010";
        ram_buffer(67930) := X"AFC50014";
        ram_buffer(67931) := X"AFC60018";
        ram_buffer(67932) := X"8FC20010";
        ram_buffer(67933) := X"00000000";
        ram_buffer(67934) := X"AFC20004";
        ram_buffer(67935) := X"8FC20010";
        ram_buffer(67936) := X"00000000";
        ram_buffer(67937) := X"30420003";
        ram_buffer(67938) := X"14400024";
        ram_buffer(67939) := X"00000000";
        ram_buffer(67940) := X"8FC20010";
        ram_buffer(67941) := X"00000000";
        ram_buffer(67942) := X"AFC20000";
        ram_buffer(67943) := X"10000005";
        ram_buffer(67944) := X"00000000";
        ram_buffer(67945) := X"8FC20000";
        ram_buffer(67946) := X"00000000";
        ram_buffer(67947) := X"24420004";
        ram_buffer(67948) := X"AFC20000";
        ram_buffer(67949) := X"8FC20000";
        ram_buffer(67950) := X"00000000";
        ram_buffer(67951) := X"8C430000";
        ram_buffer(67952) := X"3C02FEFE";
        ram_buffer(67953) := X"3442FEFF";
        ram_buffer(67954) := X"00621821";
        ram_buffer(67955) := X"8FC20000";
        ram_buffer(67956) := X"00000000";
        ram_buffer(67957) := X"8C420000";
        ram_buffer(67958) := X"00000000";
        ram_buffer(67959) := X"00021027";
        ram_buffer(67960) := X"00621824";
        ram_buffer(67961) := X"3C028080";
        ram_buffer(67962) := X"34428080";
        ram_buffer(67963) := X"00621024";
        ram_buffer(67964) := X"1040FFEC";
        ram_buffer(67965) := X"00000000";
        ram_buffer(67966) := X"8FC20000";
        ram_buffer(67967) := X"00000000";
        ram_buffer(67968) := X"AFC20010";
        ram_buffer(67969) := X"10000005";
        ram_buffer(67970) := X"00000000";
        ram_buffer(67971) := X"8FC20010";
        ram_buffer(67972) := X"00000000";
        ram_buffer(67973) := X"24420001";
        ram_buffer(67974) := X"AFC20010";
        ram_buffer(67975) := X"8FC20010";
        ram_buffer(67976) := X"00000000";
        ram_buffer(67977) := X"80420000";
        ram_buffer(67978) := X"00000000";
        ram_buffer(67979) := X"1440FFF7";
        ram_buffer(67980) := X"00000000";
        ram_buffer(67981) := X"10000008";
        ram_buffer(67982) := X"00000000";
        ram_buffer(67983) := X"8FC20018";
        ram_buffer(67984) := X"00000000";
        ram_buffer(67985) := X"14400004";
        ram_buffer(67986) := X"00000000";
        ram_buffer(67987) := X"8FC20010";
        ram_buffer(67988) := X"00000000";
        ram_buffer(67989) := X"A0400000";
        ram_buffer(67990) := X"8FC20018";
        ram_buffer(67991) := X"00000000";
        ram_buffer(67992) := X"2443FFFF";
        ram_buffer(67993) := X"AFC30018";
        ram_buffer(67994) := X"10400010";
        ram_buffer(67995) := X"00000000";
        ram_buffer(67996) := X"8FC20010";
        ram_buffer(67997) := X"00000000";
        ram_buffer(67998) := X"24430001";
        ram_buffer(67999) := X"AFC30010";
        ram_buffer(68000) := X"8FC30014";
        ram_buffer(68001) := X"00000000";
        ram_buffer(68002) := X"24640001";
        ram_buffer(68003) := X"AFC40014";
        ram_buffer(68004) := X"80630000";
        ram_buffer(68005) := X"00000000";
        ram_buffer(68006) := X"A0430000";
        ram_buffer(68007) := X"80420000";
        ram_buffer(68008) := X"00000000";
        ram_buffer(68009) := X"1440FFE5";
        ram_buffer(68010) := X"00000000";
        ram_buffer(68011) := X"8FC20004";
        ram_buffer(68012) := X"03C0E821";
        ram_buffer(68013) := X"8FBE000C";
        ram_buffer(68014) := X"27BD0010";
        ram_buffer(68015) := X"03E00008";
        ram_buffer(68016) := X"00000000";
        ram_buffer(68017) := X"27BDFFD8";
        ram_buffer(68018) := X"AFBF0024";
        ram_buffer(68019) := X"AFBE0020";
        ram_buffer(68020) := X"AFB0001C";
        ram_buffer(68021) := X"03A0F021";
        ram_buffer(68022) := X"AFC40028";
        ram_buffer(68023) := X"AFC5002C";
        ram_buffer(68024) := X"00C08021";
        ram_buffer(68025) := X"8FC20028";
        ram_buffer(68026) := X"00000000";
        ram_buffer(68027) := X"AFC20010";
        ram_buffer(68028) := X"8FC20010";
        ram_buffer(68029) := X"00000000";
        ram_buffer(68030) := X"1040000A";
        ram_buffer(68031) := X"00000000";
        ram_buffer(68032) := X"8FC20010";
        ram_buffer(68033) := X"00000000";
        ram_buffer(68034) := X"8C420038";
        ram_buffer(68035) := X"00000000";
        ram_buffer(68036) := X"14400004";
        ram_buffer(68037) := X"00000000";
        ram_buffer(68038) := X"8FC40010";
        ram_buffer(68039) := X"0C027069";
        ram_buffer(68040) := X"00000000";
        ram_buffer(68041) := X"8E020008";
        ram_buffer(68042) := X"00000000";
        ram_buffer(68043) := X"2442FFFF";
        ram_buffer(68044) := X"AE020008";
        ram_buffer(68045) := X"8E020008";
        ram_buffer(68046) := X"00000000";
        ram_buffer(68047) := X"04410027";
        ram_buffer(68048) := X"00000000";
        ram_buffer(68049) := X"8E030008";
        ram_buffer(68050) := X"8E020018";
        ram_buffer(68051) := X"00000000";
        ram_buffer(68052) := X"0062102A";
        ram_buffer(68053) := X"1440001A";
        ram_buffer(68054) := X"00000000";
        ram_buffer(68055) := X"8E020000";
        ram_buffer(68056) := X"8FC3002C";
        ram_buffer(68057) := X"00000000";
        ram_buffer(68058) := X"306300FF";
        ram_buffer(68059) := X"A0430000";
        ram_buffer(68060) := X"8E020000";
        ram_buffer(68061) := X"00000000";
        ram_buffer(68062) := X"90430000";
        ram_buffer(68063) := X"2402000A";
        ram_buffer(68064) := X"10620008";
        ram_buffer(68065) := X"00000000";
        ram_buffer(68066) := X"8E020000";
        ram_buffer(68067) := X"00000000";
        ram_buffer(68068) := X"24430001";
        ram_buffer(68069) := X"AE030000";
        ram_buffer(68070) := X"90420000";
        ram_buffer(68071) := X"1000001A";
        ram_buffer(68072) := X"00000000";
        ram_buffer(68073) := X"02003021";
        ram_buffer(68074) := X"2405000A";
        ram_buffer(68075) := X"8FC40028";
        ram_buffer(68076) := X"0C02FA03";
        ram_buffer(68077) := X"00000000";
        ram_buffer(68078) := X"10000013";
        ram_buffer(68079) := X"00000000";
        ram_buffer(68080) := X"02003021";
        ram_buffer(68081) := X"8FC5002C";
        ram_buffer(68082) := X"8FC40028";
        ram_buffer(68083) := X"0C02FA03";
        ram_buffer(68084) := X"00000000";
        ram_buffer(68085) := X"1000000C";
        ram_buffer(68086) := X"00000000";
        ram_buffer(68087) := X"8E020000";
        ram_buffer(68088) := X"8FC3002C";
        ram_buffer(68089) := X"00000000";
        ram_buffer(68090) := X"306300FF";
        ram_buffer(68091) := X"A0430000";
        ram_buffer(68092) := X"8E020000";
        ram_buffer(68093) := X"00000000";
        ram_buffer(68094) := X"24430001";
        ram_buffer(68095) := X"AE030000";
        ram_buffer(68096) := X"90420000";
        ram_buffer(68097) := X"00000000";
        ram_buffer(68098) := X"AFC20014";
        ram_buffer(68099) := X"8FC20014";
        ram_buffer(68100) := X"03C0E821";
        ram_buffer(68101) := X"8FBF0024";
        ram_buffer(68102) := X"8FBE0020";
        ram_buffer(68103) := X"8FB0001C";
        ram_buffer(68104) := X"27BD0028";
        ram_buffer(68105) := X"03E00008";
        ram_buffer(68106) := X"00000000";
        ram_buffer(68107) := X"27BDFFD0";
        ram_buffer(68108) := X"AFBF002C";
        ram_buffer(68109) := X"AFBE0028";
        ram_buffer(68110) := X"AFB00024";
        ram_buffer(68111) := X"03A0F021";
        ram_buffer(68112) := X"AFC40030";
        ram_buffer(68113) := X"00A08021";
        ram_buffer(68114) := X"8F828098";
        ram_buffer(68115) := X"00000000";
        ram_buffer(68116) := X"AFC20010";
        ram_buffer(68117) := X"8FC20010";
        ram_buffer(68118) := X"00000000";
        ram_buffer(68119) := X"AFC20014";
        ram_buffer(68120) := X"8FC20014";
        ram_buffer(68121) := X"00000000";
        ram_buffer(68122) := X"1040000A";
        ram_buffer(68123) := X"00000000";
        ram_buffer(68124) := X"8FC20014";
        ram_buffer(68125) := X"00000000";
        ram_buffer(68126) := X"8C420038";
        ram_buffer(68127) := X"00000000";
        ram_buffer(68128) := X"14400004";
        ram_buffer(68129) := X"00000000";
        ram_buffer(68130) := X"8FC40014";
        ram_buffer(68131) := X"0C027069";
        ram_buffer(68132) := X"00000000";
        ram_buffer(68133) := X"8E020008";
        ram_buffer(68134) := X"00000000";
        ram_buffer(68135) := X"2442FFFF";
        ram_buffer(68136) := X"AE020008";
        ram_buffer(68137) := X"8E020008";
        ram_buffer(68138) := X"00000000";
        ram_buffer(68139) := X"04410027";
        ram_buffer(68140) := X"00000000";
        ram_buffer(68141) := X"8E030008";
        ram_buffer(68142) := X"8E020018";
        ram_buffer(68143) := X"00000000";
        ram_buffer(68144) := X"0062102A";
        ram_buffer(68145) := X"1440001A";
        ram_buffer(68146) := X"00000000";
        ram_buffer(68147) := X"8E020000";
        ram_buffer(68148) := X"8FC30030";
        ram_buffer(68149) := X"00000000";
        ram_buffer(68150) := X"306300FF";
        ram_buffer(68151) := X"A0430000";
        ram_buffer(68152) := X"8E020000";
        ram_buffer(68153) := X"00000000";
        ram_buffer(68154) := X"90430000";
        ram_buffer(68155) := X"2402000A";
        ram_buffer(68156) := X"10620008";
        ram_buffer(68157) := X"00000000";
        ram_buffer(68158) := X"8E020000";
        ram_buffer(68159) := X"00000000";
        ram_buffer(68160) := X"24430001";
        ram_buffer(68161) := X"AE030000";
        ram_buffer(68162) := X"90420000";
        ram_buffer(68163) := X"1000001A";
        ram_buffer(68164) := X"00000000";
        ram_buffer(68165) := X"02003021";
        ram_buffer(68166) := X"2405000A";
        ram_buffer(68167) := X"8FC40010";
        ram_buffer(68168) := X"0C02FA03";
        ram_buffer(68169) := X"00000000";
        ram_buffer(68170) := X"10000013";
        ram_buffer(68171) := X"00000000";
        ram_buffer(68172) := X"02003021";
        ram_buffer(68173) := X"8FC50030";
        ram_buffer(68174) := X"8FC40010";
        ram_buffer(68175) := X"0C02FA03";
        ram_buffer(68176) := X"00000000";
        ram_buffer(68177) := X"1000000C";
        ram_buffer(68178) := X"00000000";
        ram_buffer(68179) := X"8E020000";
        ram_buffer(68180) := X"8FC30030";
        ram_buffer(68181) := X"00000000";
        ram_buffer(68182) := X"306300FF";
        ram_buffer(68183) := X"A0430000";
        ram_buffer(68184) := X"8E020000";
        ram_buffer(68185) := X"00000000";
        ram_buffer(68186) := X"24430001";
        ram_buffer(68187) := X"AE030000";
        ram_buffer(68188) := X"90420000";
        ram_buffer(68189) := X"00000000";
        ram_buffer(68190) := X"AFC20018";
        ram_buffer(68191) := X"8FC20018";
        ram_buffer(68192) := X"03C0E821";
        ram_buffer(68193) := X"8FBF002C";
        ram_buffer(68194) := X"8FBE0028";
        ram_buffer(68195) := X"8FB00024";
        ram_buffer(68196) := X"27BD0030";
        ram_buffer(68197) := X"03E00008";
        ram_buffer(68198) := X"00000000";
        ram_buffer(68199) := X"00E04021";
        ram_buffer(68200) := X"00A04821";
        ram_buffer(68201) := X"14C00053";
        ram_buffer(68202) := X"00805021";
        ram_buffer(68203) := X"0087102B";
        ram_buffer(68204) := X"1040006E";
        ram_buffer(68205) := X"3C020001";
        ram_buffer(68206) := X"00E2102B";
        ram_buffer(68207) := X"10400162";
        ram_buffer(68208) := X"3C020100";
        ram_buffer(68209) := X"2CE30100";
        ram_buffer(68210) := X"2C630001";
        ram_buffer(68211) := X"000318C0";
        ram_buffer(68212) := X"3C02100D";
        ram_buffer(68213) := X"00673006";
        ram_buffer(68214) := X"2442B660";
        ram_buffer(68215) := X"00C21021";
        ram_buffer(68216) := X"90420000";
        ram_buffer(68217) := X"00000000";
        ram_buffer(68218) := X"00431821";
        ram_buffer(68219) := X"24020020";
        ram_buffer(68220) := X"00431023";
        ram_buffer(68221) := X"10400007";
        ram_buffer(68222) := X"00085C02";
        ram_buffer(68223) := X"00443004";
        ram_buffer(68224) := X"00651806";
        ram_buffer(68225) := X"00474004";
        ram_buffer(68226) := X"00665025";
        ram_buffer(68227) := X"00454804";
        ram_buffer(68228) := X"00085C02";
        ram_buffer(68229) := X"15600002";
        ram_buffer(68230) := X"014B001B";
        ram_buffer(68231) := X"0007000D";
        ram_buffer(68232) := X"3105FFFF";
        ram_buffer(68233) := X"00091C02";
        ram_buffer(68234) := X"00001012";
        ram_buffer(68235) := X"00003010";
        ram_buffer(68236) := X"00063400";
        ram_buffer(68237) := X"00661825";
        ram_buffer(68238) := X"00A20018";
        ram_buffer(68239) := X"00002012";
        ram_buffer(68240) := X"0064382B";
        ram_buffer(68241) := X"00000000";
        ram_buffer(68242) := X"15600002";
        ram_buffer(68243) := X"014B001B";
        ram_buffer(68244) := X"0007000D";
        ram_buffer(68245) := X"10E00009";
        ram_buffer(68246) := X"00000000";
        ram_buffer(68247) := X"00681821";
        ram_buffer(68248) := X"0068302B";
        ram_buffer(68249) := X"14C00004";
        ram_buffer(68250) := X"2447FFFF";
        ram_buffer(68251) := X"0064302B";
        ram_buffer(68252) := X"14C0015F";
        ram_buffer(68253) := X"2442FFFE";
        ram_buffer(68254) := X"00E01021";
        ram_buffer(68255) := X"00642023";
        ram_buffer(68256) := X"3129FFFF";
        ram_buffer(68257) := X"15600002";
        ram_buffer(68258) := X"008B001B";
        ram_buffer(68259) := X"0007000D";
        ram_buffer(68260) := X"00001812";
        ram_buffer(68261) := X"00003010";
        ram_buffer(68262) := X"00063400";
        ram_buffer(68263) := X"01264825";
        ram_buffer(68264) := X"00A30018";
        ram_buffer(68265) := X"00002812";
        ram_buffer(68266) := X"0125302B";
        ram_buffer(68267) := X"00000000";
        ram_buffer(68268) := X"15600002";
        ram_buffer(68269) := X"008B001B";
        ram_buffer(68270) := X"0007000D";
        ram_buffer(68271) := X"10C00008";
        ram_buffer(68272) := X"01094821";
        ram_buffer(68273) := X"0128402B";
        ram_buffer(68274) := X"15000128";
        ram_buffer(68275) := X"2464FFFF";
        ram_buffer(68276) := X"0125482B";
        ram_buffer(68277) := X"11200125";
        ram_buffer(68278) := X"00000000";
        ram_buffer(68279) := X"2463FFFE";
        ram_buffer(68280) := X"00021400";
        ram_buffer(68281) := X"00431825";
        ram_buffer(68282) := X"00001021";
        ram_buffer(68283) := X"03E00008";
        ram_buffer(68284) := X"00000000";
        ram_buffer(68285) := X"0086102B";
        ram_buffer(68286) := X"14400070";
        ram_buffer(68287) := X"00001821";
        ram_buffer(68288) := X"3C020001";
        ram_buffer(68289) := X"00C2102B";
        ram_buffer(68290) := X"1440006F";
        ram_buffer(68291) := X"2CC80100";
        ram_buffer(68292) := X"3C020100";
        ram_buffer(68293) := X"00C2102B";
        ram_buffer(68294) := X"10400002";
        ram_buffer(68295) := X"24080018";
        ram_buffer(68296) := X"24080010";
        ram_buffer(68297) := X"3C02100D";
        ram_buffer(68298) := X"01061806";
        ram_buffer(68299) := X"2442B660";
        ram_buffer(68300) := X"00621021";
        ram_buffer(68301) := X"90420000";
        ram_buffer(68302) := X"240B0020";
        ram_buffer(68303) := X"00484021";
        ram_buffer(68304) := X"01685823";
        ram_buffer(68305) := X"1560006C";
        ram_buffer(68306) := X"01071006";
        ram_buffer(68307) := X"00C4302B";
        ram_buffer(68308) := X"14C00114";
        ram_buffer(68309) := X"00000000";
        ram_buffer(68310) := X"00A7182B";
        ram_buffer(68311) := X"38630001";
        ram_buffer(68312) := X"00001021";
        ram_buffer(68313) := X"03E00008";
        ram_buffer(68314) := X"00000000";
        ram_buffer(68315) := X"14E00008";
        ram_buffer(68316) := X"0102102B";
        ram_buffer(68317) := X"24020001";
        ram_buffer(68318) := X"14E00002";
        ram_buffer(68319) := X"0047001B";
        ram_buffer(68320) := X"0007000D";
        ram_buffer(68321) := X"00004012";
        ram_buffer(68322) := X"3C020001";
        ram_buffer(68323) := X"0102102B";
        ram_buffer(68324) := X"1440009C";
        ram_buffer(68325) := X"2D070100";
        ram_buffer(68326) := X"3C020100";
        ram_buffer(68327) := X"0102102B";
        ram_buffer(68328) := X"10400002";
        ram_buffer(68329) := X"24070018";
        ram_buffer(68330) := X"24070010";
        ram_buffer(68331) := X"3C02100D";
        ram_buffer(68332) := X"00E81806";
        ram_buffer(68333) := X"2442B660";
        ram_buffer(68334) := X"00621021";
        ram_buffer(68335) := X"90420000";
        ram_buffer(68336) := X"240C0020";
        ram_buffer(68337) := X"00473821";
        ram_buffer(68338) := X"01876023";
        ram_buffer(68339) := X"15800099";
        ram_buffer(68340) := X"00000000";
        ram_buffer(68341) := X"00882023";
        ram_buffer(68342) := X"00085402";
        ram_buffer(68343) := X"3105FFFF";
        ram_buffer(68344) := X"24020001";
        ram_buffer(68345) := X"15400002";
        ram_buffer(68346) := X"008A001B";
        ram_buffer(68347) := X"0007000D";
        ram_buffer(68348) := X"00091C02";
        ram_buffer(68349) := X"00003012";
        ram_buffer(68350) := X"00003810";
        ram_buffer(68351) := X"00073C00";
        ram_buffer(68352) := X"00671825";
        ram_buffer(68353) := X"00C50018";
        ram_buffer(68354) := X"00005812";
        ram_buffer(68355) := X"006B382B";
        ram_buffer(68356) := X"00000000";
        ram_buffer(68357) := X"15400002";
        ram_buffer(68358) := X"008A001B";
        ram_buffer(68359) := X"0007000D";
        ram_buffer(68360) := X"10E0000A";
        ram_buffer(68361) := X"006B2023";
        ram_buffer(68362) := X"00681821";
        ram_buffer(68363) := X"0068202B";
        ram_buffer(68364) := X"14800004";
        ram_buffer(68365) := X"24C7FFFF";
        ram_buffer(68366) := X"006B202B";
        ram_buffer(68367) := X"148000EA";
        ram_buffer(68368) := X"24C6FFFE";
        ram_buffer(68369) := X"00E03021";
        ram_buffer(68370) := X"006B2023";
        ram_buffer(68371) := X"3129FFFF";
        ram_buffer(68372) := X"15400002";
        ram_buffer(68373) := X"008A001B";
        ram_buffer(68374) := X"0007000D";
        ram_buffer(68375) := X"00001812";
        ram_buffer(68376) := X"00003810";
        ram_buffer(68377) := X"00073C00";
        ram_buffer(68378) := X"01274825";
        ram_buffer(68379) := X"00650018";
        ram_buffer(68380) := X"00002812";
        ram_buffer(68381) := X"0125382B";
        ram_buffer(68382) := X"00000000";
        ram_buffer(68383) := X"15400002";
        ram_buffer(68384) := X"008A001B";
        ram_buffer(68385) := X"0007000D";
        ram_buffer(68386) := X"10E00008";
        ram_buffer(68387) := X"01094821";
        ram_buffer(68388) := X"0128402B";
        ram_buffer(68389) := X"150000B1";
        ram_buffer(68390) := X"2464FFFF";
        ram_buffer(68391) := X"0125482B";
        ram_buffer(68392) := X"112000AE";
        ram_buffer(68393) := X"00000000";
        ram_buffer(68394) := X"2463FFFE";
        ram_buffer(68395) := X"00063400";
        ram_buffer(68396) := X"00C31825";
        ram_buffer(68397) := X"03E00008";
        ram_buffer(68398) := X"00000000";
        ram_buffer(68399) := X"00001021";
        ram_buffer(68400) := X"03E00008";
        ram_buffer(68401) := X"00000000";
        ram_buffer(68402) := X"2D080001";
        ram_buffer(68403) := X"000840C0";
        ram_buffer(68404) := X"3C02100D";
        ram_buffer(68405) := X"01061806";
        ram_buffer(68406) := X"2442B660";
        ram_buffer(68407) := X"00621021";
        ram_buffer(68408) := X"90420000";
        ram_buffer(68409) := X"240B0020";
        ram_buffer(68410) := X"00484021";
        ram_buffer(68411) := X"01685823";
        ram_buffer(68412) := X"1160FF96";
        ram_buffer(68413) := X"01071006";
        ram_buffer(68414) := X"01663004";
        ram_buffer(68415) := X"00C23025";
        ram_buffer(68416) := X"01046806";
        ram_buffer(68417) := X"00066402";
        ram_buffer(68418) := X"15800002";
        ram_buffer(68419) := X"01AC001B";
        ram_buffer(68420) := X"0007000D";
        ram_buffer(68421) := X"30CEFFFF";
        ram_buffer(68422) := X"01054006";
        ram_buffer(68423) := X"01642004";
        ram_buffer(68424) := X"01042025";
        ram_buffer(68425) := X"00045402";
        ram_buffer(68426) := X"00001012";
        ram_buffer(68427) := X"00007810";
        ram_buffer(68428) := X"000F4400";
        ram_buffer(68429) := X"01484025";
        ram_buffer(68430) := X"01C20018";
        ram_buffer(68431) := X"00004812";
        ram_buffer(68432) := X"0109182B";
        ram_buffer(68433) := X"00000000";
        ram_buffer(68434) := X"15800002";
        ram_buffer(68435) := X"01AC001B";
        ram_buffer(68436) := X"0007000D";
        ram_buffer(68437) := X"10600006";
        ram_buffer(68438) := X"01673804";
        ram_buffer(68439) := X"01064021";
        ram_buffer(68440) := X"0106182B";
        ram_buffer(68441) := X"10600097";
        ram_buffer(68442) := X"244AFFFF";
        ram_buffer(68443) := X"01401021";
        ram_buffer(68444) := X"01094823";
        ram_buffer(68445) := X"3088FFFF";
        ram_buffer(68446) := X"15800002";
        ram_buffer(68447) := X"012C001B";
        ram_buffer(68448) := X"0007000D";
        ram_buffer(68449) := X"00001812";
        ram_buffer(68450) := X"00006810";
        ram_buffer(68451) := X"000D2400";
        ram_buffer(68452) := X"01042025";
        ram_buffer(68453) := X"01C30018";
        ram_buffer(68454) := X"00005012";
        ram_buffer(68455) := X"008A402B";
        ram_buffer(68456) := X"00000000";
        ram_buffer(68457) := X"15800002";
        ram_buffer(68458) := X"012C001B";
        ram_buffer(68459) := X"0007000D";
        ram_buffer(68460) := X"11000006";
        ram_buffer(68461) := X"00000000";
        ram_buffer(68462) := X"00862021";
        ram_buffer(68463) := X"0086402B";
        ram_buffer(68464) := X"1100007B";
        ram_buffer(68465) := X"2469FFFF";
        ram_buffer(68466) := X"01201821";
        ram_buffer(68467) := X"00021400";
        ram_buffer(68468) := X"00431825";
        ram_buffer(68469) := X"008A2023";
        ram_buffer(68470) := X"00670019";
        ram_buffer(68471) := X"00003010";
        ram_buffer(68472) := X"0086102B";
        ram_buffer(68473) := X"00003812";
        ram_buffer(68474) := X"14400066";
        ram_buffer(68475) := X"00000000";
        ram_buffer(68476) := X"10860060";
        ram_buffer(68477) := X"00000000";
        ram_buffer(68478) := X"00001021";
        ram_buffer(68479) := X"03E00008";
        ram_buffer(68480) := X"00000000";
        ram_buffer(68481) := X"2CE70001";
        ram_buffer(68482) := X"000738C0";
        ram_buffer(68483) := X"3C02100D";
        ram_buffer(68484) := X"00E81806";
        ram_buffer(68485) := X"2442B660";
        ram_buffer(68486) := X"00621021";
        ram_buffer(68487) := X"90420000";
        ram_buffer(68488) := X"240C0020";
        ram_buffer(68489) := X"00473821";
        ram_buffer(68490) := X"01876023";
        ram_buffer(68491) := X"1180FF69";
        ram_buffer(68492) := X"00000000";
        ram_buffer(68493) := X"01884004";
        ram_buffer(68494) := X"00E46806";
        ram_buffer(68495) := X"00085402";
        ram_buffer(68496) := X"15400002";
        ram_buffer(68497) := X"01AA001B";
        ram_buffer(68498) := X"0007000D";
        ram_buffer(68499) := X"310BFFFF";
        ram_buffer(68500) := X"01843004";
        ram_buffer(68501) := X"01854804";
        ram_buffer(68502) := X"00E53806";
        ram_buffer(68503) := X"00E63025";
        ram_buffer(68504) := X"00062402";
        ram_buffer(68505) := X"00001012";
        ram_buffer(68506) := X"00001810";
        ram_buffer(68507) := X"00031C00";
        ram_buffer(68508) := X"00831825";
        ram_buffer(68509) := X"00006012";
        ram_buffer(68510) := X"00000000";
        ram_buffer(68511) := X"00000000";
        ram_buffer(68512) := X"01620018";
        ram_buffer(68513) := X"00002812";
        ram_buffer(68514) := X"0065102B";
        ram_buffer(68515) := X"00000000";
        ram_buffer(68516) := X"15400002";
        ram_buffer(68517) := X"01AA001B";
        ram_buffer(68518) := X"0007000D";
        ram_buffer(68519) := X"1040000A";
        ram_buffer(68520) := X"00000000";
        ram_buffer(68521) := X"00681821";
        ram_buffer(68522) := X"0068102B";
        ram_buffer(68523) := X"1440004C";
        ram_buffer(68524) := X"2584FFFF";
        ram_buffer(68525) := X"0065102B";
        ram_buffer(68526) := X"10400049";
        ram_buffer(68527) := X"00000000";
        ram_buffer(68528) := X"258CFFFE";
        ram_buffer(68529) := X"00681821";
        ram_buffer(68530) := X"00652823";
        ram_buffer(68531) := X"30C7FFFF";
        ram_buffer(68532) := X"15400002";
        ram_buffer(68533) := X"00AA001B";
        ram_buffer(68534) := X"0007000D";
        ram_buffer(68535) := X"00001012";
        ram_buffer(68536) := X"00001810";
        ram_buffer(68537) := X"00031C00";
        ram_buffer(68538) := X"00E31825";
        ram_buffer(68539) := X"01620018";
        ram_buffer(68540) := X"00002012";
        ram_buffer(68541) := X"0064302B";
        ram_buffer(68542) := X"00000000";
        ram_buffer(68543) := X"15400002";
        ram_buffer(68544) := X"00AA001B";
        ram_buffer(68545) := X"0007000D";
        ram_buffer(68546) := X"10C0000A";
        ram_buffer(68547) := X"00000000";
        ram_buffer(68548) := X"00681821";
        ram_buffer(68549) := X"0068282B";
        ram_buffer(68550) := X"14A0002F";
        ram_buffer(68551) := X"2446FFFF";
        ram_buffer(68552) := X"0064282B";
        ram_buffer(68553) := X"10A0002C";
        ram_buffer(68554) := X"00000000";
        ram_buffer(68555) := X"2442FFFE";
        ram_buffer(68556) := X"00681821";
        ram_buffer(68557) := X"000C6400";
        ram_buffer(68558) := X"00642023";
        ram_buffer(68559) := X"01821025";
        ram_buffer(68560) := X"1000FF28";
        ram_buffer(68561) := X"01602821";
        ram_buffer(68562) := X"00E2102B";
        ram_buffer(68563) := X"10400013";
        ram_buffer(68564) := X"00000000";
        ram_buffer(68565) := X"1000FE9E";
        ram_buffer(68566) := X"24030010";
        ram_buffer(68567) := X"00801821";
        ram_buffer(68568) := X"00063400";
        ram_buffer(68569) := X"1000FF53";
        ram_buffer(68570) := X"00C31825";
        ram_buffer(68571) := X"1000FEDC";
        ram_buffer(68572) := X"00801821";
        ram_buffer(68573) := X"01652804";
        ram_buffer(68574) := X"00A7282B";
        ram_buffer(68575) := X"10A0FF9E";
        ram_buffer(68576) := X"00000000";
        ram_buffer(68577) := X"2463FFFF";
        ram_buffer(68578) := X"00001021";
        ram_buffer(68579) := X"03E00008";
        ram_buffer(68580) := X"00000000";
        ram_buffer(68581) := X"1000FF05";
        ram_buffer(68582) := X"24070018";
        ram_buffer(68583) := X"1000FE8C";
        ram_buffer(68584) := X"24030018";
        ram_buffer(68585) := X"24030001";
        ram_buffer(68586) := X"1000FF94";
        ram_buffer(68587) := X"00001021";
        ram_buffer(68588) := X"008A402B";
        ram_buffer(68589) := X"1100FF84";
        ram_buffer(68590) := X"2463FFFE";
        ram_buffer(68591) := X"1000FF83";
        ram_buffer(68592) := X"00862021";
        ram_buffer(68593) := X"0109182B";
        ram_buffer(68594) := X"1060FF68";
        ram_buffer(68595) := X"2442FFFE";
        ram_buffer(68596) := X"1000FF67";
        ram_buffer(68597) := X"01064021";
        ram_buffer(68598) := X"1000FFD6";
        ram_buffer(68599) := X"00C01021";
        ram_buffer(68600) := X"1000FFB9";
        ram_buffer(68601) := X"00806021";
        ram_buffer(68602) := X"1000FF17";
        ram_buffer(68603) := X"00681821";
        ram_buffer(68604) := X"1000FEA2";
        ram_buffer(68605) := X"00681821";
        ram_buffer(68606) := X"00E04021";
        ram_buffer(68607) := X"00A06821";
        ram_buffer(68608) := X"14C00052";
        ram_buffer(68609) := X"00801021";
        ram_buffer(68610) := X"0087182B";
        ram_buffer(68611) := X"10600071";
        ram_buffer(68612) := X"3C030001";
        ram_buffer(68613) := X"00E3182B";
        ram_buffer(68614) := X"10600164";
        ram_buffer(68615) := X"3C030100";
        ram_buffer(68616) := X"2CEB0100";
        ram_buffer(68617) := X"2D6B0001";
        ram_buffer(68618) := X"000B58C0";
        ram_buffer(68619) := X"3C03100D";
        ram_buffer(68620) := X"01673006";
        ram_buffer(68621) := X"2463B660";
        ram_buffer(68622) := X"00C31821";
        ram_buffer(68623) := X"906A0000";
        ram_buffer(68624) := X"24030020";
        ram_buffer(68625) := X"014B4821";
        ram_buffer(68626) := X"00695823";
        ram_buffer(68627) := X"11600007";
        ram_buffer(68628) := X"00086402";
        ram_buffer(68629) := X"01642004";
        ram_buffer(68630) := X"01254806";
        ram_buffer(68631) := X"01674004";
        ram_buffer(68632) := X"01241025";
        ram_buffer(68633) := X"01656804";
        ram_buffer(68634) := X"00086402";
        ram_buffer(68635) := X"15800002";
        ram_buffer(68636) := X"004C001B";
        ram_buffer(68637) := X"0007000D";
        ram_buffer(68638) := X"3107FFFF";
        ram_buffer(68639) := X"000D5402";
        ram_buffer(68640) := X"00007012";
        ram_buffer(68641) := X"00004810";
        ram_buffer(68642) := X"00094C00";
        ram_buffer(68643) := X"01495025";
        ram_buffer(68644) := X"00EE0018";
        ram_buffer(68645) := X"00007012";
        ram_buffer(68646) := X"014E782B";
        ram_buffer(68647) := X"00000000";
        ram_buffer(68648) := X"15800002";
        ram_buffer(68649) := X"004C001B";
        ram_buffer(68650) := X"0007000D";
        ram_buffer(68651) := X"11E00009";
        ram_buffer(68652) := X"014E4823";
        ram_buffer(68653) := X"01485021";
        ram_buffer(68654) := X"0148102B";
        ram_buffer(68655) := X"14400005";
        ram_buffer(68656) := X"014E4823";
        ram_buffer(68657) := X"014E102B";
        ram_buffer(68658) := X"14400153";
        ram_buffer(68659) := X"00000000";
        ram_buffer(68660) := X"014E4823";
        ram_buffer(68661) := X"31A6FFFF";
        ram_buffer(68662) := X"15800002";
        ram_buffer(68663) := X"012C001B";
        ram_buffer(68664) := X"0007000D";
        ram_buffer(68665) := X"00001812";
        ram_buffer(68666) := X"00002010";
        ram_buffer(68667) := X"00042400";
        ram_buffer(68668) := X"00C42025";
        ram_buffer(68669) := X"00E30018";
        ram_buffer(68670) := X"00001812";
        ram_buffer(68671) := X"0083102B";
        ram_buffer(68672) := X"00000000";
        ram_buffer(68673) := X"15800002";
        ram_buffer(68674) := X"012C001B";
        ram_buffer(68675) := X"0007000D";
        ram_buffer(68676) := X"10400009";
        ram_buffer(68677) := X"00000000";
        ram_buffer(68678) := X"00882021";
        ram_buffer(68679) := X"0088102B";
        ram_buffer(68680) := X"14400005";
        ram_buffer(68681) := X"00000000";
        ram_buffer(68682) := X"0083102B";
        ram_buffer(68683) := X"10400002";
        ram_buffer(68684) := X"00000000";
        ram_buffer(68685) := X"00882021";
        ram_buffer(68686) := X"00831823";
        ram_buffer(68687) := X"00001021";
        ram_buffer(68688) := X"01631806";
        ram_buffer(68689) := X"03E00008";
        ram_buffer(68690) := X"00000000";
        ram_buffer(68691) := X"0086182B";
        ram_buffer(68692) := X"14600073";
        ram_buffer(68693) := X"00A01821";
        ram_buffer(68694) := X"3C030001";
        ram_buffer(68695) := X"00C3182B";
        ram_buffer(68696) := X"14600072";
        ram_buffer(68697) := X"2CC80100";
        ram_buffer(68698) := X"3C030100";
        ram_buffer(68699) := X"00C3182B";
        ram_buffer(68700) := X"10600002";
        ram_buffer(68701) := X"24080018";
        ram_buffer(68702) := X"24080010";
        ram_buffer(68703) := X"3C03100D";
        ram_buffer(68704) := X"01064806";
        ram_buffer(68705) := X"2463B660";
        ram_buffer(68706) := X"01231821";
        ram_buffer(68707) := X"90630000";
        ram_buffer(68708) := X"240F0020";
        ram_buffer(68709) := X"00681821";
        ram_buffer(68710) := X"01E37823";
        ram_buffer(68711) := X"15E0006F";
        ram_buffer(68712) := X"00000000";
        ram_buffer(68713) := X"00C4182B";
        ram_buffer(68714) := X"14600005";
        ram_buffer(68715) := X"00A71823";
        ram_buffer(68716) := X"00A7182B";
        ram_buffer(68717) := X"1460011A";
        ram_buffer(68718) := X"00000000";
        ram_buffer(68719) := X"00A71823";
        ram_buffer(68720) := X"00862023";
        ram_buffer(68721) := X"00A3102B";
        ram_buffer(68722) := X"00821023";
        ram_buffer(68723) := X"03E00008";
        ram_buffer(68724) := X"00000000";
        ram_buffer(68725) := X"14E00007";
        ram_buffer(68726) := X"3C020001";
        ram_buffer(68727) := X"24020001";
        ram_buffer(68728) := X"14E00002";
        ram_buffer(68729) := X"0047001B";
        ram_buffer(68730) := X"0007000D";
        ram_buffer(68731) := X"00004012";
        ram_buffer(68732) := X"3C020001";
        ram_buffer(68733) := X"0102102B";
        ram_buffer(68734) := X"144000A5";
        ram_buffer(68735) := X"2D090100";
        ram_buffer(68736) := X"3C020100";
        ram_buffer(68737) := X"0102102B";
        ram_buffer(68738) := X"10400002";
        ram_buffer(68739) := X"24090018";
        ram_buffer(68740) := X"24090010";
        ram_buffer(68741) := X"3C02100D";
        ram_buffer(68742) := X"01281806";
        ram_buffer(68743) := X"2442B660";
        ram_buffer(68744) := X"00621021";
        ram_buffer(68745) := X"90470000";
        ram_buffer(68746) := X"24030020";
        ram_buffer(68747) := X"00E94821";
        ram_buffer(68748) := X"00695823";
        ram_buffer(68749) := X"156000A2";
        ram_buffer(68750) := X"00000000";
        ram_buffer(68751) := X"00884823";
        ram_buffer(68752) := X"00086402";
        ram_buffer(68753) := X"3102FFFF";
        ram_buffer(68754) := X"15800002";
        ram_buffer(68755) := X"012C001B";
        ram_buffer(68756) := X"0007000D";
        ram_buffer(68757) := X"000D5402";
        ram_buffer(68758) := X"00003012";
        ram_buffer(68759) := X"00001810";
        ram_buffer(68760) := X"00031C00";
        ram_buffer(68761) := X"01435025";
        ram_buffer(68762) := X"00C20018";
        ram_buffer(68763) := X"00003012";
        ram_buffer(68764) := X"0146182B";
        ram_buffer(68765) := X"00000000";
        ram_buffer(68766) := X"15800002";
        ram_buffer(68767) := X"012C001B";
        ram_buffer(68768) := X"0007000D";
        ram_buffer(68769) := X"10600009";
        ram_buffer(68770) := X"01464823";
        ram_buffer(68771) := X"01485021";
        ram_buffer(68772) := X"0148182B";
        ram_buffer(68773) := X"14600005";
        ram_buffer(68774) := X"01464823";
        ram_buffer(68775) := X"0146182B";
        ram_buffer(68776) := X"146000DB";
        ram_buffer(68777) := X"00000000";
        ram_buffer(68778) := X"01464823";
        ram_buffer(68779) := X"31AAFFFF";
        ram_buffer(68780) := X"15800002";
        ram_buffer(68781) := X"012C001B";
        ram_buffer(68782) := X"0007000D";
        ram_buffer(68783) := X"00001812";
        ram_buffer(68784) := X"00003010";
        ram_buffer(68785) := X"00063400";
        ram_buffer(68786) := X"00000000";
        ram_buffer(68787) := X"00620018";
        ram_buffer(68788) := X"01461025";
        ram_buffer(68789) := X"00001812";
        ram_buffer(68790) := X"0043202B";
        ram_buffer(68791) := X"00000000";
        ram_buffer(68792) := X"15800002";
        ram_buffer(68793) := X"012C001B";
        ram_buffer(68794) := X"0007000D";
        ram_buffer(68795) := X"10800008";
        ram_buffer(68796) := X"00000000";
        ram_buffer(68797) := X"00481021";
        ram_buffer(68798) := X"0048202B";
        ram_buffer(68799) := X"14800004";
        ram_buffer(68800) := X"0043202B";
        ram_buffer(68801) := X"10800002";
        ram_buffer(68802) := X"00000000";
        ram_buffer(68803) := X"00481021";
        ram_buffer(68804) := X"00431823";
        ram_buffer(68805) := X"01631806";
        ram_buffer(68806) := X"1000FF8A";
        ram_buffer(68807) := X"00001021";
        ram_buffer(68808) := X"00801021";
        ram_buffer(68809) := X"03E00008";
        ram_buffer(68810) := X"00000000";
        ram_buffer(68811) := X"2D080001";
        ram_buffer(68812) := X"000840C0";
        ram_buffer(68813) := X"3C03100D";
        ram_buffer(68814) := X"01064806";
        ram_buffer(68815) := X"2463B660";
        ram_buffer(68816) := X"01231821";
        ram_buffer(68817) := X"90630000";
        ram_buffer(68818) := X"240F0020";
        ram_buffer(68819) := X"00681821";
        ram_buffer(68820) := X"01E37823";
        ram_buffer(68821) := X"11E0FF93";
        ram_buffer(68822) := X"00000000";
        ram_buffer(68823) := X"01E63004";
        ram_buffer(68824) := X"00675006";
        ram_buffer(68825) := X"00CA5025";
        ram_buffer(68826) := X"0064C806";
        ram_buffer(68827) := X"000AC402";
        ram_buffer(68828) := X"17000002";
        ram_buffer(68829) := X"0338001B";
        ram_buffer(68830) := X"0007000D";
        ram_buffer(68831) := X"3142FFFF";
        ram_buffer(68832) := X"01E43004";
        ram_buffer(68833) := X"00654806";
        ram_buffer(68834) := X"01264825";
        ram_buffer(68835) := X"00097402";
        ram_buffer(68836) := X"01E73004";
        ram_buffer(68837) := X"00005812";
        ram_buffer(68838) := X"00006810";
        ram_buffer(68839) := X"000D6C00";
        ram_buffer(68840) := X"01CD6825";
        ram_buffer(68841) := X"004B0018";
        ram_buffer(68842) := X"00006012";
        ram_buffer(68843) := X"01AC202B";
        ram_buffer(68844) := X"00000000";
        ram_buffer(68845) := X"17000002";
        ram_buffer(68846) := X"0338001B";
        ram_buffer(68847) := X"0007000D";
        ram_buffer(68848) := X"10800006";
        ram_buffer(68849) := X"01E52804";
        ram_buffer(68850) := X"01AA6821";
        ram_buffer(68851) := X"01AA202B";
        ram_buffer(68852) := X"1080008A";
        ram_buffer(68853) := X"2567FFFF";
        ram_buffer(68854) := X"00E05821";
        ram_buffer(68855) := X"01AC6023";
        ram_buffer(68856) := X"3129FFFF";
        ram_buffer(68857) := X"17000002";
        ram_buffer(68858) := X"0198001B";
        ram_buffer(68859) := X"0007000D";
        ram_buffer(68860) := X"00002012";
        ram_buffer(68861) := X"00004010";
        ram_buffer(68862) := X"00084400";
        ram_buffer(68863) := X"01284025";
        ram_buffer(68864) := X"00440018";
        ram_buffer(68865) := X"00001012";
        ram_buffer(68866) := X"0102382B";
        ram_buffer(68867) := X"00000000";
        ram_buffer(68868) := X"17000002";
        ram_buffer(68869) := X"0198001B";
        ram_buffer(68870) := X"0007000D";
        ram_buffer(68871) := X"10E00006";
        ram_buffer(68872) := X"00000000";
        ram_buffer(68873) := X"010A4021";
        ram_buffer(68874) := X"010A382B";
        ram_buffer(68875) := X"10E0006E";
        ram_buffer(68876) := X"2489FFFF";
        ram_buffer(68877) := X"01202021";
        ram_buffer(68878) := X"000B4C00";
        ram_buffer(68879) := X"01245825";
        ram_buffer(68880) := X"01024023";
        ram_buffer(68881) := X"01660019";
        ram_buffer(68882) := X"00006010";
        ram_buffer(68883) := X"010C102B";
        ram_buffer(68884) := X"00006812";
        ram_buffer(68885) := X"1440005A";
        ram_buffer(68886) := X"00000000";
        ram_buffer(68887) := X"110C0073";
        ram_buffer(68888) := X"00000000";
        ram_buffer(68889) := X"010C4023";
        ram_buffer(68890) := X"00003012";
        ram_buffer(68891) := X"00A63023";
        ram_buffer(68892) := X"00A6282B";
        ram_buffer(68893) := X"01054023";
        ram_buffer(68894) := X"00682804";
        ram_buffer(68895) := X"01E63006";
        ram_buffer(68896) := X"01E81006";
        ram_buffer(68897) := X"00A61825";
        ram_buffer(68898) := X"03E00008";
        ram_buffer(68899) := X"00000000";
        ram_buffer(68900) := X"2D290001";
        ram_buffer(68901) := X"000948C0";
        ram_buffer(68902) := X"3C02100D";
        ram_buffer(68903) := X"01281806";
        ram_buffer(68904) := X"2442B660";
        ram_buffer(68905) := X"00621021";
        ram_buffer(68906) := X"90470000";
        ram_buffer(68907) := X"24030020";
        ram_buffer(68908) := X"00E94821";
        ram_buffer(68909) := X"00695823";
        ram_buffer(68910) := X"1160FF60";
        ram_buffer(68911) := X"00000000";
        ram_buffer(68912) := X"01684004";
        ram_buffer(68913) := X"01247006";
        ram_buffer(68914) := X"00086402";
        ram_buffer(68915) := X"15800002";
        ram_buffer(68916) := X"01CC001B";
        ram_buffer(68917) := X"0007000D";
        ram_buffer(68918) := X"3103FFFF";
        ram_buffer(68919) := X"01642004";
        ram_buffer(68920) := X"01254806";
        ram_buffer(68921) := X"01244825";
        ram_buffer(68922) := X"00095402";
        ram_buffer(68923) := X"00003812";
        ram_buffer(68924) := X"00003010";
        ram_buffer(68925) := X"00063400";
        ram_buffer(68926) := X"01463025";
        ram_buffer(68927) := X"00670018";
        ram_buffer(68928) := X"00003812";
        ram_buffer(68929) := X"00C7102B";
        ram_buffer(68930) := X"00000000";
        ram_buffer(68931) := X"15800002";
        ram_buffer(68932) := X"01CC001B";
        ram_buffer(68933) := X"0007000D";
        ram_buffer(68934) := X"10400008";
        ram_buffer(68935) := X"01656804";
        ram_buffer(68936) := X"00C83021";
        ram_buffer(68937) := X"00C8102B";
        ram_buffer(68938) := X"14400004";
        ram_buffer(68939) := X"00C7102B";
        ram_buffer(68940) := X"10400002";
        ram_buffer(68941) := X"00000000";
        ram_buffer(68942) := X"00C83021";
        ram_buffer(68943) := X"00C73823";
        ram_buffer(68944) := X"312AFFFF";
        ram_buffer(68945) := X"15800002";
        ram_buffer(68946) := X"00EC001B";
        ram_buffer(68947) := X"0007000D";
        ram_buffer(68948) := X"00002012";
        ram_buffer(68949) := X"00004810";
        ram_buffer(68950) := X"00094C00";
        ram_buffer(68951) := X"01495025";
        ram_buffer(68952) := X"00640018";
        ram_buffer(68953) := X"00002012";
        ram_buffer(68954) := X"0144102B";
        ram_buffer(68955) := X"00000000";
        ram_buffer(68956) := X"15800002";
        ram_buffer(68957) := X"00EC001B";
        ram_buffer(68958) := X"0007000D";
        ram_buffer(68959) := X"10400008";
        ram_buffer(68960) := X"00000000";
        ram_buffer(68961) := X"01485021";
        ram_buffer(68962) := X"0148102B";
        ram_buffer(68963) := X"14400005";
        ram_buffer(68964) := X"01444823";
        ram_buffer(68965) := X"0144102B";
        ram_buffer(68966) := X"10400002";
        ram_buffer(68967) := X"01485021";
        ram_buffer(68968) := X"01444823";
        ram_buffer(68969) := X"1000FF28";
        ram_buffer(68970) := X"00601021";
        ram_buffer(68971) := X"00E3182B";
        ram_buffer(68972) := X"1060000B";
        ram_buffer(68973) := X"00000000";
        ram_buffer(68974) := X"1000FE9C";
        ram_buffer(68975) := X"240B0010";
        ram_buffer(68976) := X"01A63023";
        ram_buffer(68977) := X"018A5023";
        ram_buffer(68978) := X"01A6102B";
        ram_buffer(68979) := X"01421023";
        ram_buffer(68980) := X"1000FFA6";
        ram_buffer(68981) := X"01024023";
        ram_buffer(68982) := X"1000FF0E";
        ram_buffer(68983) := X"24090018";
        ram_buffer(68984) := X"1000FE92";
        ram_buffer(68985) := X"240B0018";
        ram_buffer(68986) := X"0102382B";
        ram_buffer(68987) := X"10E0FF91";
        ram_buffer(68988) := X"2484FFFE";
        ram_buffer(68989) := X"1000FF90";
        ram_buffer(68990) := X"010A4021";
        ram_buffer(68991) := X"01AC202B";
        ram_buffer(68992) := X"1080FF75";
        ram_buffer(68993) := X"256BFFFE";
        ram_buffer(68994) := X"1000FF74";
        ram_buffer(68995) := X"01AA6821";
        ram_buffer(68996) := X"1000FF25";
        ram_buffer(68997) := X"01485021";
        ram_buffer(68998) := X"1000FEAD";
        ram_buffer(68999) := X"01485021";
        ram_buffer(69000) := X"00A01821";
        ram_buffer(69001) := X"03E00008";
        ram_buffer(69002) := X"00000000";
        ram_buffer(69003) := X"00AD102B";
        ram_buffer(69004) := X"1440FFE3";
        ram_buffer(69005) := X"00000000";
        ram_buffer(69006) := X"00003012";
        ram_buffer(69007) := X"1000FF8B";
        ram_buffer(69008) := X"00004021";
        ram_buffer(69009) := X"27BDFFE0";
        ram_buffer(69010) := X"3C06007F";
        ram_buffer(69011) := X"34C6FFFF";
        ram_buffer(69012) := X"00053DC2";
        ram_buffer(69013) := X"AFB00010";
        ram_buffer(69014) := X"000485C2";
        ram_buffer(69015) := X"00C41824";
        ram_buffer(69016) := X"AFB10014";
        ram_buffer(69017) := X"00C53024";
        ram_buffer(69018) := X"321000FF";
        ram_buffer(69019) := X"30E700FF";
        ram_buffer(69020) := X"00048FC2";
        ram_buffer(69021) := X"00052FC2";
        ram_buffer(69022) := X"AFBF001C";
        ram_buffer(69023) := X"AFB20018";
        ram_buffer(69024) := X"000318C0";
        ram_buffer(69025) := X"000630C0";
        ram_buffer(69026) := X"12250056";
        ram_buffer(69027) := X"02071023";
        ram_buffer(69028) := X"18400094";
        ram_buffer(69029) := X"00000000";
        ram_buffer(69030) := X"14E00020";
        ram_buffer(69031) := X"00000000";
        ram_buffer(69032) := X"14C00079";
        ram_buffer(69033) := X"2442FFFF";
        ram_buffer(69034) := X"240200FF";
        ram_buffer(69035) := X"1202007A";
        ram_buffer(69036) := X"00000000";
        ram_buffer(69037) := X"000310C2";
        ram_buffer(69038) := X"240300FF";
        ram_buffer(69039) := X"1603006C";
        ram_buffer(69040) := X"00000000";
        ram_buffer(69041) := X"10400077";
        ram_buffer(69042) := X"02202021";
        ram_buffer(69043) := X"3C05003F";
        ram_buffer(69044) := X"34A5FFFF";
        ram_buffer(69045) := X"00451824";
        ram_buffer(69046) := X"14600098";
        ram_buffer(69047) := X"00000000";
        ram_buffer(69048) := X"00002021";
        ram_buffer(69049) := X"241000FF";
        ram_buffer(69050) := X"3C03007F";
        ram_buffer(69051) := X"3463FFFF";
        ram_buffer(69052) := X"001085C0";
        ram_buffer(69053) := X"8FBF001C";
        ram_buffer(69054) := X"00A31824";
        ram_buffer(69055) := X"00701825";
        ram_buffer(69056) := X"000417C0";
        ram_buffer(69057) := X"8FB20018";
        ram_buffer(69058) := X"8FB10014";
        ram_buffer(69059) := X"8FB00010";
        ram_buffer(69060) := X"00621025";
        ram_buffer(69061) := X"03E00008";
        ram_buffer(69062) := X"27BD0020";
        ram_buffer(69063) := X"240400FF";
        ram_buffer(69064) := X"1204005D";
        ram_buffer(69065) := X"3C040400";
        ram_buffer(69066) := X"00C43025";
        ram_buffer(69067) := X"2844001C";
        ram_buffer(69068) := X"10800094";
        ram_buffer(69069) := X"00022023";
        ram_buffer(69070) := X"00862004";
        ram_buffer(69071) := X"00463006";
        ram_buffer(69072) := X"0004102B";
        ram_buffer(69073) := X"00C23025";
        ram_buffer(69074) := X"00661823";
        ram_buffer(69075) := X"3C120400";
        ram_buffer(69076) := X"00721024";
        ram_buffer(69077) := X"1040005F";
        ram_buffer(69078) := X"30620007";
        ram_buffer(69079) := X"2652FFFF";
        ram_buffer(69080) := X"00729024";
        ram_buffer(69081) := X"0C031D29";
        ram_buffer(69082) := X"02402021";
        ram_buffer(69083) := X"2442FFFB";
        ram_buffer(69084) := X"0050182A";
        ram_buffer(69085) := X"14600069";
        ram_buffer(69086) := X"00529004";
        ram_buffer(69087) := X"00501023";
        ram_buffer(69088) := X"24430001";
        ram_buffer(69089) := X"00031023";
        ram_buffer(69090) := X"00521004";
        ram_buffer(69091) := X"00729006";
        ram_buffer(69092) := X"0002182B";
        ram_buffer(69093) := X"02431825";
        ram_buffer(69094) := X"30720007";
        ram_buffer(69095) := X"00008021";
        ram_buffer(69096) := X"12400006";
        ram_buffer(69097) := X"3C020400";
        ram_buffer(69098) := X"3062000F";
        ram_buffer(69099) := X"24040004";
        ram_buffer(69100) := X"10440002";
        ram_buffer(69101) := X"3C020400";
        ram_buffer(69102) := X"24630004";
        ram_buffer(69103) := X"00621024";
        ram_buffer(69104) := X"1040FFBC";
        ram_buffer(69105) := X"240200FF";
        ram_buffer(69106) := X"26100001";
        ram_buffer(69107) := X"12020034";
        ram_buffer(69108) := X"00031980";
        ram_buffer(69109) := X"00032A42";
        ram_buffer(69110) := X"321000FF";
        ram_buffer(69111) := X"1000FFC2";
        ram_buffer(69112) := X"02202021";
        ram_buffer(69113) := X"18400059";
        ram_buffer(69114) := X"00000000";
        ram_buffer(69115) := X"10E00030";
        ram_buffer(69116) := X"240400FF";
        ram_buffer(69117) := X"12040028";
        ram_buffer(69118) := X"3C040400";
        ram_buffer(69119) := X"00C43025";
        ram_buffer(69120) := X"2844001C";
        ram_buffer(69121) := X"10800094";
        ram_buffer(69122) := X"00022023";
        ram_buffer(69123) := X"00862004";
        ram_buffer(69124) := X"00463006";
        ram_buffer(69125) := X"0004102B";
        ram_buffer(69126) := X"00C21025";
        ram_buffer(69127) := X"00621821";
        ram_buffer(69128) := X"3C020400";
        ram_buffer(69129) := X"00621024";
        ram_buffer(69130) := X"1040002A";
        ram_buffer(69131) := X"30620007";
        ram_buffer(69132) := X"26100001";
        ram_buffer(69133) := X"240200FF";
        ram_buffer(69134) := X"12020019";
        ram_buffer(69135) := X"3C02FBFF";
        ram_buffer(69136) := X"3442FFFF";
        ram_buffer(69137) := X"00621024";
        ram_buffer(69138) := X"00021042";
        ram_buffer(69139) := X"30630001";
        ram_buffer(69140) := X"00431825";
        ram_buffer(69141) := X"30620007";
        ram_buffer(69142) := X"1440FFD4";
        ram_buffer(69143) := X"3062000F";
        ram_buffer(69144) := X"000310C2";
        ram_buffer(69145) := X"240300FF";
        ram_buffer(69146) := X"1203FF96";
        ram_buffer(69147) := X"00000000";
        ram_buffer(69148) := X"3C06007F";
        ram_buffer(69149) := X"34C6FFFF";
        ram_buffer(69150) := X"00462824";
        ram_buffer(69151) := X"321000FF";
        ram_buffer(69152) := X"1000FF99";
        ram_buffer(69153) := X"02202021";
        ram_buffer(69154) := X"1040FFAF";
        ram_buffer(69155) := X"240400FF";
        ram_buffer(69156) := X"1604FFA7";
        ram_buffer(69157) := X"2844001C";
        ram_buffer(69158) := X"1460FF87";
        ram_buffer(69159) := X"000310C2";
        ram_buffer(69160) := X"02202021";
        ram_buffer(69161) := X"241000FF";
        ram_buffer(69162) := X"1000FF8F";
        ram_buffer(69163) := X"00002821";
        ram_buffer(69164) := X"10C0FF7D";
        ram_buffer(69165) := X"2442FFFF";
        ram_buffer(69166) := X"14400052";
        ram_buffer(69167) := X"240400FF";
        ram_buffer(69168) := X"1000FFD7";
        ram_buffer(69169) := X"00661821";
        ram_buffer(69170) := X"108000C9";
        ram_buffer(69171) := X"00801821";
        ram_buffer(69172) := X"30620007";
        ram_buffer(69173) := X"1440FFB4";
        ram_buffer(69174) := X"000310C2";
        ram_buffer(69175) := X"1000FF77";
        ram_buffer(69176) := X"240300FF";
        ram_buffer(69177) := X"14400029";
        ram_buffer(69178) := X"00000000";
        ram_buffer(69179) := X"26020001";
        ram_buffer(69180) := X"304200FF";
        ram_buffer(69181) := X"28420002";
        ram_buffer(69182) := X"1440004E";
        ram_buffer(69183) := X"00669023";
        ram_buffer(69184) := X"3C020400";
        ram_buffer(69185) := X"02421024";
        ram_buffer(69186) := X"10400031";
        ram_buffer(69187) := X"00000000";
        ram_buffer(69188) := X"00C39023";
        ram_buffer(69189) := X"1000FF93";
        ram_buffer(69190) := X"00A08821";
        ram_buffer(69191) := X"3C03FBFF";
        ram_buffer(69192) := X"3463FFFF";
        ram_buffer(69193) := X"02431824";
        ram_buffer(69194) := X"02028023";
        ram_buffer(69195) := X"1000FF9C";
        ram_buffer(69196) := X"32520007";
        ram_buffer(69197) := X"00008821";
        ram_buffer(69198) := X"3443FFFF";
        ram_buffer(69199) := X"00602821";
        ram_buffer(69200) := X"02202021";
        ram_buffer(69201) := X"1000FF68";
        ram_buffer(69202) := X"241000FF";
        ram_buffer(69203) := X"14400044";
        ram_buffer(69204) := X"26040001";
        ram_buffer(69205) := X"308200FF";
        ram_buffer(69206) := X"28420002";
        ram_buffer(69207) := X"1440002F";
        ram_buffer(69208) := X"240200FF";
        ram_buffer(69209) := X"1082FFCE";
        ram_buffer(69210) := X"00661821";
        ram_buffer(69211) := X"00031842";
        ram_buffer(69212) := X"30620007";
        ram_buffer(69213) := X"1440FF8C";
        ram_buffer(69214) := X"00808021";
        ram_buffer(69215) := X"1000FFB9";
        ram_buffer(69216) := X"000310C2";
        ram_buffer(69217) := X"1000FF70";
        ram_buffer(69218) := X"24060001";
        ram_buffer(69219) := X"12000015";
        ram_buffer(69220) := X"240400FF";
        ram_buffer(69221) := X"10E40054";
        ram_buffer(69222) := X"3C040400";
        ram_buffer(69223) := X"00021023";
        ram_buffer(69224) := X"00641825";
        ram_buffer(69225) := X"2844001C";
        ram_buffer(69226) := X"10800075";
        ram_buffer(69227) := X"00022023";
        ram_buffer(69228) := X"00832004";
        ram_buffer(69229) := X"00431006";
        ram_buffer(69230) := X"0004182B";
        ram_buffer(69231) := X"00431825";
        ram_buffer(69232) := X"00C31823";
        ram_buffer(69233) := X"00E08021";
        ram_buffer(69234) := X"1000FF60";
        ram_buffer(69235) := X"00A08821";
        ram_buffer(69236) := X"1640FF64";
        ram_buffer(69237) := X"00000000";
        ram_buffer(69238) := X"00008821";
        ram_buffer(69239) := X"1000FFA4";
        ram_buffer(69240) := X"00008021";
        ram_buffer(69241) := X"1460003C";
        ram_buffer(69242) := X"00021027";
        ram_buffer(69243) := X"240200FF";
        ram_buffer(69244) := X"10E2003D";
        ram_buffer(69245) := X"00C01821";
        ram_buffer(69246) := X"00E08021";
        ram_buffer(69247) := X"1000FF2D";
        ram_buffer(69248) := X"00A08821";
        ram_buffer(69249) := X"1604FF7F";
        ram_buffer(69250) := X"2844001C";
        ram_buffer(69251) := X"1060FFA5";
        ram_buffer(69252) := X"02202021";
        ram_buffer(69253) := X"1000FF28";
        ram_buffer(69254) := X"000310C2";
        ram_buffer(69255) := X"16000021";
        ram_buffer(69256) := X"00000000";
        ram_buffer(69257) := X"1460005A";
        ram_buffer(69258) := X"00000000";
        ram_buffer(69259) := X"1000FF21";
        ram_buffer(69260) := X"00C01821";
        ram_buffer(69261) := X"16000013";
        ram_buffer(69262) := X"00000000";
        ram_buffer(69263) := X"1460003D";
        ram_buffer(69264) := X"00000000";
        ram_buffer(69265) := X"10C00050";
        ram_buffer(69266) := X"00001021";
        ram_buffer(69267) := X"00C01821";
        ram_buffer(69268) := X"1000FF18";
        ram_buffer(69269) := X"00A08821";
        ram_buffer(69270) := X"1000FF70";
        ram_buffer(69271) := X"24020001";
        ram_buffer(69272) := X"16000026";
        ram_buffer(69273) := X"240400FF";
        ram_buffer(69274) := X"1460003C";
        ram_buffer(69275) := X"00021027";
        ram_buffer(69276) := X"240200FF";
        ram_buffer(69277) := X"10E2003D";
        ram_buffer(69278) := X"00C01821";
        ram_buffer(69279) := X"1000FF0D";
        ram_buffer(69280) := X"00E08021";
        ram_buffer(69281) := X"14600009";
        ram_buffer(69282) := X"00000000";
        ram_buffer(69283) := X"10C0FFA9";
        ram_buffer(69284) := X"3C02003F";
        ram_buffer(69285) := X"00C01821";
        ram_buffer(69286) := X"00A08821";
        ram_buffer(69287) := X"1000FF05";
        ram_buffer(69288) := X"241000FF";
        ram_buffer(69289) := X"10600033";
        ram_buffer(69290) := X"00000000";
        ram_buffer(69291) := X"10C0FF01";
        ram_buffer(69292) := X"241000FF";
        ram_buffer(69293) := X"000318C2";
        ram_buffer(69294) := X"000610C2";
        ram_buffer(69295) := X"00431025";
        ram_buffer(69296) := X"3C040040";
        ram_buffer(69297) := X"00441024";
        ram_buffer(69298) := X"1440003F";
        ram_buffer(69299) := X"00000000";
        ram_buffer(69300) := X"1000FEF8";
        ram_buffer(69301) := X"000318C0";
        ram_buffer(69302) := X"1040FFB9";
        ram_buffer(69303) := X"240400FF";
        ram_buffer(69304) := X"14E4FFB1";
        ram_buffer(69305) := X"2844001C";
        ram_buffer(69306) := X"10C0003B";
        ram_buffer(69307) := X"00C01821";
        ram_buffer(69308) := X"241000FF";
        ram_buffer(69309) := X"1000FEEF";
        ram_buffer(69310) := X"00A08821";
        ram_buffer(69311) := X"10E4001B";
        ram_buffer(69312) := X"3C040400";
        ram_buffer(69313) := X"00021023";
        ram_buffer(69314) := X"00641825";
        ram_buffer(69315) := X"2844001C";
        ram_buffer(69316) := X"10800033";
        ram_buffer(69317) := X"00022023";
        ram_buffer(69318) := X"00832004";
        ram_buffer(69319) := X"00431006";
        ram_buffer(69320) := X"0004182B";
        ram_buffer(69321) := X"00431825";
        ram_buffer(69322) := X"00661821";
        ram_buffer(69323) := X"1000FF3C";
        ram_buffer(69324) := X"00E08021";
        ram_buffer(69325) := X"10C0FEE0";
        ram_buffer(69326) := X"000310C2";
        ram_buffer(69327) := X"00662023";
        ram_buffer(69328) := X"3C020400";
        ram_buffer(69329) := X"00821024";
        ram_buffer(69330) := X"1040FF5F";
        ram_buffer(69331) := X"00C31823";
        ram_buffer(69332) := X"30720007";
        ram_buffer(69333) := X"1000FF12";
        ram_buffer(69334) := X"00A08821";
        ram_buffer(69335) := X"1040FFF2";
        ram_buffer(69336) := X"240400FF";
        ram_buffer(69337) := X"14E4FFEA";
        ram_buffer(69338) := X"2844001C";
        ram_buffer(69339) := X"10C0FF4D";
        ram_buffer(69340) := X"02202021";
        ram_buffer(69341) := X"00C01821";
        ram_buffer(69342) := X"1000FECE";
        ram_buffer(69343) := X"241000FF";
        ram_buffer(69344) := X"1000FF8F";
        ram_buffer(69345) := X"24030001";
        ram_buffer(69346) := X"1000FF39";
        ram_buffer(69347) := X"00008821";
        ram_buffer(69348) := X"10C0FEC9";
        ram_buffer(69349) := X"000310C2";
        ram_buffer(69350) := X"00661821";
        ram_buffer(69351) := X"3C020400";
        ram_buffer(69352) := X"00621024";
        ram_buffer(69353) := X"1040FF4B";
        ram_buffer(69354) := X"30620007";
        ram_buffer(69355) := X"3C04FBFF";
        ram_buffer(69356) := X"3484FFFF";
        ram_buffer(69357) := X"24100001";
        ram_buffer(69358) := X"1440FEFB";
        ram_buffer(69359) := X"00641824";
        ram_buffer(69360) := X"1000FF28";
        ram_buffer(69361) := X"000310C2";
        ram_buffer(69362) := X"3C0301FF";
        ram_buffer(69363) := X"00008821";
        ram_buffer(69364) := X"1000FEB8";
        ram_buffer(69365) := X"3463FFF8";
        ram_buffer(69366) := X"1000FF31";
        ram_buffer(69367) := X"00A08821";
        ram_buffer(69368) := X"24030001";
        ram_buffer(69369) := X"00661821";
        ram_buffer(69370) := X"1000FF0D";
        ram_buffer(69371) := X"00E08021";
        ram_buffer(69372) := X"1000FF1F";
        ram_buffer(69373) := X"00008821";
        ram_buffer(69374) := X"27BDFFC0";
        ram_buffer(69375) := X"000415C2";
        ram_buffer(69376) := X"3C03007F";
        ram_buffer(69377) := X"3463FFFF";
        ram_buffer(69378) := X"AFB50030";
        ram_buffer(69379) := X"AFB10020";
        ram_buffer(69380) := X"0004AFC2";
        ram_buffer(69381) := X"305100FF";
        ram_buffer(69382) := X"AFB60034";
        ram_buffer(69383) := X"AFB4002C";
        ram_buffer(69384) := X"AFBF003C";
        ram_buffer(69385) := X"AFB70038";
        ram_buffer(69386) := X"AFB30028";
        ram_buffer(69387) := X"AFB20024";
        ram_buffer(69388) := X"AFB0001C";
        ram_buffer(69389) := X"0064A024";
        ram_buffer(69390) := X"12200053";
        ram_buffer(69391) := X"02A0B021";
        ram_buffer(69392) := X"240200FF";
        ram_buffer(69393) := X"12220023";
        ram_buffer(69394) := X"3C040080";
        ram_buffer(69395) := X"02842025";
        ram_buffer(69396) := X"0004A0C0";
        ram_buffer(69397) := X"2631FF81";
        ram_buffer(69398) := X"00009021";
        ram_buffer(69399) := X"0000B821";
        ram_buffer(69400) := X"000515C2";
        ram_buffer(69401) := X"3C10007F";
        ram_buffer(69402) := X"3610FFFF";
        ram_buffer(69403) := X"304200FF";
        ram_buffer(69404) := X"02058024";
        ram_buffer(69405) := X"10400022";
        ram_buffer(69406) := X"00059FC2";
        ram_buffer(69407) := X"240300FF";
        ram_buffer(69408) := X"10430046";
        ram_buffer(69409) := X"2E050001";
        ram_buffer(69410) := X"3C030080";
        ram_buffer(69411) := X"02038025";
        ram_buffer(69412) := X"001080C0";
        ram_buffer(69413) := X"2442FF81";
        ram_buffer(69414) := X"00002821";
        ram_buffer(69415) := X"00B23025";
        ram_buffer(69416) := X"02221021";
        ram_buffer(69417) := X"2CC30010";
        ram_buffer(69418) := X"02B34026";
        ram_buffer(69419) := X"10600066";
        ram_buffer(69420) := X"24490001";
        ram_buffer(69421) := X"3C07100D";
        ram_buffer(69422) := X"00063080";
        ram_buffer(69423) := X"24E7B5A0";
        ram_buffer(69424) := X"00E63021";
        ram_buffer(69425) := X"8CC30000";
        ram_buffer(69426) := X"00000000";
        ram_buffer(69427) := X"00600008";
        ram_buffer(69428) := X"00000000";
        ram_buffer(69429) := X"16800042";
        ram_buffer(69430) := X"2412000C";
        ram_buffer(69431) := X"000515C2";
        ram_buffer(69432) := X"3C10007F";
        ram_buffer(69433) := X"3610FFFF";
        ram_buffer(69434) := X"304200FF";
        ram_buffer(69435) := X"24120008";
        ram_buffer(69436) := X"24170002";
        ram_buffer(69437) := X"02058024";
        ram_buffer(69438) := X"1440FFE0";
        ram_buffer(69439) := X"00059FC2";
        ram_buffer(69440) := X"16000039";
        ram_buffer(69441) := X"00000000";
        ram_buffer(69442) := X"1000FFE4";
        ram_buffer(69443) := X"24050001";
        ram_buffer(69444) := X"02604021";
        ram_buffer(69445) := X"24020002";
        ram_buffer(69446) := X"10A20024";
        ram_buffer(69447) := X"01002021";
        ram_buffer(69448) := X"24020003";
        ram_buffer(69449) := X"10A200A3";
        ram_buffer(69450) := X"24020001";
        ram_buffer(69451) := X"14A20057";
        ram_buffer(69452) := X"01201021";
        ram_buffer(69453) := X"01002021";
        ram_buffer(69454) := X"00008021";
        ram_buffer(69455) := X"00001821";
        ram_buffer(69456) := X"001015C0";
        ram_buffer(69457) := X"3C10007F";
        ram_buffer(69458) := X"3610FFFF";
        ram_buffer(69459) := X"00708024";
        ram_buffer(69460) := X"8FBF003C";
        ram_buffer(69461) := X"02028025";
        ram_buffer(69462) := X"00041FC0";
        ram_buffer(69463) := X"02031025";
        ram_buffer(69464) := X"8FB70038";
        ram_buffer(69465) := X"8FB60034";
        ram_buffer(69466) := X"8FB50030";
        ram_buffer(69467) := X"8FB4002C";
        ram_buffer(69468) := X"8FB30028";
        ram_buffer(69469) := X"8FB20024";
        ram_buffer(69470) := X"8FB10020";
        ram_buffer(69471) := X"8FB0001C";
        ram_buffer(69472) := X"03E00008";
        ram_buffer(69473) := X"27BD0040";
        ram_buffer(69474) := X"1680000B";
        ram_buffer(69475) := X"02802021";
        ram_buffer(69476) := X"24120004";
        ram_buffer(69477) := X"1000FFB2";
        ram_buffer(69478) := X"24170001";
        ram_buffer(69479) := X"24030003";
        ram_buffer(69480) := X"1000FFBE";
        ram_buffer(69481) := X"00652823";
        ram_buffer(69482) := X"01002021";
        ram_buffer(69483) := X"241000FF";
        ram_buffer(69484) := X"1000FFE3";
        ram_buffer(69485) := X"00001821";
        ram_buffer(69486) := X"0C031D29";
        ram_buffer(69487) := X"AFA50010";
        ram_buffer(69488) := X"2443FFFB";
        ram_buffer(69489) := X"2411FF8A";
        ram_buffer(69490) := X"0074A004";
        ram_buffer(69491) := X"02228823";
        ram_buffer(69492) := X"00009021";
        ram_buffer(69493) := X"8FA50010";
        ram_buffer(69494) := X"1000FFA1";
        ram_buffer(69495) := X"0000B821";
        ram_buffer(69496) := X"1000FF9F";
        ram_buffer(69497) := X"24170003";
        ram_buffer(69498) := X"0C031D29";
        ram_buffer(69499) := X"02002021";
        ram_buffer(69500) := X"2443FFFB";
        ram_buffer(69501) := X"2406FF8A";
        ram_buffer(69502) := X"00708004";
        ram_buffer(69503) := X"00C21023";
        ram_buffer(69504) := X"1000FFA6";
        ram_buffer(69505) := X"00002821";
        ram_buffer(69506) := X"3C10003F";
        ram_buffer(69507) := X"3604FFFF";
        ram_buffer(69508) := X"0000B021";
        ram_buffer(69509) := X"3C10007F";
        ram_buffer(69510) := X"3610FFFF";
        ram_buffer(69511) := X"00901824";
        ram_buffer(69512) := X"32C40001";
        ram_buffer(69513) := X"1000FFC6";
        ram_buffer(69514) := X"241000FF";
        ram_buffer(69515) := X"02808021";
        ram_buffer(69516) := X"1000FFB8";
        ram_buffer(69517) := X"02E02821";
        ram_buffer(69518) := X"02808021";
        ram_buffer(69519) := X"02A04021";
        ram_buffer(69520) := X"1000FFB4";
        ram_buffer(69521) := X"02E02821";
        ram_buffer(69522) := X"02900019";
        ram_buffer(69523) := X"0000A812";
        ram_buffer(69524) := X"00158682";
        ram_buffer(69525) := X"00151980";
        ram_buffer(69526) := X"0000A010";
        ram_buffer(69527) := X"00142980";
        ram_buffer(69528) := X"0003182B";
        ram_buffer(69529) := X"00B08025";
        ram_buffer(69530) := X"02038025";
        ram_buffer(69531) := X"3C030800";
        ram_buffer(69532) := X"02031824";
        ram_buffer(69533) := X"10600006";
        ram_buffer(69534) := X"2445007F";
        ram_buffer(69535) := X"00101042";
        ram_buffer(69536) := X"32100001";
        ram_buffer(69537) := X"00508025";
        ram_buffer(69538) := X"01201021";
        ram_buffer(69539) := X"2445007F";
        ram_buffer(69540) := X"18A00026";
        ram_buffer(69541) := X"32030007";
        ram_buffer(69542) := X"10600006";
        ram_buffer(69543) := X"3C030800";
        ram_buffer(69544) := X"3203000F";
        ram_buffer(69545) := X"24040004";
        ram_buffer(69546) := X"10640002";
        ram_buffer(69547) := X"3C030800";
        ram_buffer(69548) := X"26100004";
        ram_buffer(69549) := X"02031824";
        ram_buffer(69550) := X"10600004";
        ram_buffer(69551) := X"3C03F7FF";
        ram_buffer(69552) := X"3463FFFF";
        ram_buffer(69553) := X"02038024";
        ram_buffer(69554) := X"24450080";
        ram_buffer(69555) := X"28A200FF";
        ram_buffer(69556) := X"1040FFB5";
        ram_buffer(69557) := X"00000000";
        ram_buffer(69558) := X"00108180";
        ram_buffer(69559) := X"00101A42";
        ram_buffer(69560) := X"01002021";
        ram_buffer(69561) := X"1000FF96";
        ram_buffer(69562) := X"30B000FF";
        ram_buffer(69563) := X"02908025";
        ram_buffer(69564) := X"3C030040";
        ram_buffer(69565) := X"02038024";
        ram_buffer(69566) := X"1600000A";
        ram_buffer(69567) := X"2464FFFF";
        ram_buffer(69568) := X"2463FFFF";
        ram_buffer(69569) := X"02832024";
        ram_buffer(69570) := X"1480FFC2";
        ram_buffer(69571) := X"00000000";
        ram_buffer(69572) := X"3C03003F";
        ram_buffer(69573) := X"00002021";
        ram_buffer(69574) := X"241000FF";
        ram_buffer(69575) := X"1000FF88";
        ram_buffer(69576) := X"3463FFFF";
        ram_buffer(69577) := X"1000FFBB";
        ram_buffer(69578) := X"0000B021";
        ram_buffer(69579) := X"14A00017";
        ram_buffer(69580) := X"24020001";
        ram_buffer(69581) := X"00102042";
        ram_buffer(69582) := X"24050001";
        ram_buffer(69583) := X"00051823";
        ram_buffer(69584) := X"00701804";
        ram_buffer(69585) := X"0003182B";
        ram_buffer(69586) := X"00831825";
        ram_buffer(69587) := X"30620007";
        ram_buffer(69588) := X"10400006";
        ram_buffer(69589) := X"3C020400";
        ram_buffer(69590) := X"3062000F";
        ram_buffer(69591) := X"24040004";
        ram_buffer(69592) := X"10440002";
        ram_buffer(69593) := X"3C020400";
        ram_buffer(69594) := X"24630004";
        ram_buffer(69595) := X"00621024";
        ram_buffer(69596) := X"1440000C";
        ram_buffer(69597) := X"00000000";
        ram_buffer(69598) := X"00031980";
        ram_buffer(69599) := X"00031A42";
        ram_buffer(69600) := X"00008021";
        ram_buffer(69601) := X"1000FF6E";
        ram_buffer(69602) := X"01002021";
        ram_buffer(69603) := X"00452823";
        ram_buffer(69604) := X"28A2001C";
        ram_buffer(69605) := X"1040FF67";
        ram_buffer(69606) := X"00B02006";
        ram_buffer(69607) := X"1000FFE8";
        ram_buffer(69608) := X"00051823";
        ram_buffer(69609) := X"24100001";
        ram_buffer(69610) := X"00001821";
        ram_buffer(69611) := X"1000FF64";
        ram_buffer(69612) := X"01002021";
        ram_buffer(69613) := X"3C03003F";
        ram_buffer(69614) := X"3463FFFF";
        ram_buffer(69615) := X"02032024";
        ram_buffer(69616) := X"1000FFD1";
        ram_buffer(69617) := X"0100B021";
        ram_buffer(69618) := X"3C06007F";
        ram_buffer(69619) := X"27BDFFE0";
        ram_buffer(69620) := X"34C6FFFF";
        ram_buffer(69621) := X"00053DC2";
        ram_buffer(69622) := X"00C41824";
        ram_buffer(69623) := X"AFB00010";
        ram_buffer(69624) := X"00C53024";
        ram_buffer(69625) := X"000485C2";
        ram_buffer(69626) := X"30E700FF";
        ram_buffer(69627) := X"240200FF";
        ram_buffer(69628) := X"AFB10014";
        ram_buffer(69629) := X"AFBF001C";
        ram_buffer(69630) := X"AFB20018";
        ram_buffer(69631) := X"321000FF";
        ram_buffer(69632) := X"00048FC2";
        ram_buffer(69633) := X"000318C0";
        ram_buffer(69634) := X"00052FC2";
        ram_buffer(69635) := X"10E20027";
        ram_buffer(69636) := X"000630C0";
        ram_buffer(69637) := X"38A50001";
        ram_buffer(69638) := X"10B10028";
        ram_buffer(69639) := X"02071023";
        ram_buffer(69640) := X"1840009B";
        ram_buffer(69641) := X"00000000";
        ram_buffer(69642) := X"14E0004D";
        ram_buffer(69643) := X"240400FF";
        ram_buffer(69644) := X"14C0007C";
        ram_buffer(69645) := X"2442FFFF";
        ram_buffer(69646) := X"240200FF";
        ram_buffer(69647) := X"1202007D";
        ram_buffer(69648) := X"00000000";
        ram_buffer(69649) := X"000310C2";
        ram_buffer(69650) := X"240300FF";
        ram_buffer(69651) := X"1603003E";
        ram_buffer(69652) := X"00000000";
        ram_buffer(69653) := X"1040007A";
        ram_buffer(69654) := X"02202821";
        ram_buffer(69655) := X"3C05003F";
        ram_buffer(69656) := X"34A5FFFF";
        ram_buffer(69657) := X"00451824";
        ram_buffer(69658) := X"146000A3";
        ram_buffer(69659) := X"00000000";
        ram_buffer(69660) := X"00001021";
        ram_buffer(69661) := X"241000FF";
        ram_buffer(69662) := X"3C03007F";
        ram_buffer(69663) := X"3463FFFF";
        ram_buffer(69664) := X"001085C0";
        ram_buffer(69665) := X"8FBF001C";
        ram_buffer(69666) := X"00A31824";
        ram_buffer(69667) := X"00701825";
        ram_buffer(69668) := X"000217C0";
        ram_buffer(69669) := X"8FB20018";
        ram_buffer(69670) := X"8FB10014";
        ram_buffer(69671) := X"8FB00010";
        ram_buffer(69672) := X"00621025";
        ram_buffer(69673) := X"03E00008";
        ram_buffer(69674) := X"27BD0020";
        ram_buffer(69675) := X"10C0FFD9";
        ram_buffer(69676) := X"00000000";
        ram_buffer(69677) := X"14B1FFDA";
        ram_buffer(69678) := X"02071023";
        ram_buffer(69679) := X"18400092";
        ram_buffer(69680) := X"00000000";
        ram_buffer(69681) := X"10E00062";
        ram_buffer(69682) := X"240400FF";
        ram_buffer(69683) := X"12040065";
        ram_buffer(69684) := X"3C040400";
        ram_buffer(69685) := X"00C43025";
        ram_buffer(69686) := X"2844001C";
        ram_buffer(69687) := X"108000D2";
        ram_buffer(69688) := X"00022023";
        ram_buffer(69689) := X"00862004";
        ram_buffer(69690) := X"00463006";
        ram_buffer(69691) := X"0004102B";
        ram_buffer(69692) := X"00C23025";
        ram_buffer(69693) := X"00661821";
        ram_buffer(69694) := X"3C020400";
        ram_buffer(69695) := X"00621024";
        ram_buffer(69696) := X"10400090";
        ram_buffer(69697) := X"240200FF";
        ram_buffer(69698) := X"26100001";
        ram_buffer(69699) := X"1202004D";
        ram_buffer(69700) := X"30A20001";
        ram_buffer(69701) := X"3C02FBFF";
        ram_buffer(69702) := X"3442FFFF";
        ram_buffer(69703) := X"00621024";
        ram_buffer(69704) := X"00021042";
        ram_buffer(69705) := X"30630001";
        ram_buffer(69706) := X"00431825";
        ram_buffer(69707) := X"30620007";
        ram_buffer(69708) := X"1440002D";
        ram_buffer(69709) := X"00A08821";
        ram_buffer(69710) := X"000310C2";
        ram_buffer(69711) := X"240300FF";
        ram_buffer(69712) := X"1203FFC4";
        ram_buffer(69713) := X"00000000";
        ram_buffer(69714) := X"3C06007F";
        ram_buffer(69715) := X"34C6FFFF";
        ram_buffer(69716) := X"00462824";
        ram_buffer(69717) := X"321000FF";
        ram_buffer(69718) := X"1000FFC7";
        ram_buffer(69719) := X"32220001";
        ram_buffer(69720) := X"12040034";
        ram_buffer(69721) := X"3C040400";
        ram_buffer(69722) := X"00C43025";
        ram_buffer(69723) := X"2844001C";
        ram_buffer(69724) := X"10800076";
        ram_buffer(69725) := X"00022023";
        ram_buffer(69726) := X"00862004";
        ram_buffer(69727) := X"00463006";
        ram_buffer(69728) := X"0004102B";
        ram_buffer(69729) := X"00C23025";
        ram_buffer(69730) := X"00661823";
        ram_buffer(69731) := X"3C120400";
        ram_buffer(69732) := X"00721024";
        ram_buffer(69733) := X"1040003A";
        ram_buffer(69734) := X"30620007";
        ram_buffer(69735) := X"2652FFFF";
        ram_buffer(69736) := X"00729024";
        ram_buffer(69737) := X"0C031D29";
        ram_buffer(69738) := X"02402021";
        ram_buffer(69739) := X"2442FFFB";
        ram_buffer(69740) := X"0050182A";
        ram_buffer(69741) := X"14600048";
        ram_buffer(69742) := X"00529004";
        ram_buffer(69743) := X"00501023";
        ram_buffer(69744) := X"24430001";
        ram_buffer(69745) := X"00031023";
        ram_buffer(69746) := X"00521004";
        ram_buffer(69747) := X"00729006";
        ram_buffer(69748) := X"0002182B";
        ram_buffer(69749) := X"02431825";
        ram_buffer(69750) := X"30720007";
        ram_buffer(69751) := X"00008021";
        ram_buffer(69752) := X"12400006";
        ram_buffer(69753) := X"3C020400";
        ram_buffer(69754) := X"3062000F";
        ram_buffer(69755) := X"24040004";
        ram_buffer(69756) := X"10440002";
        ram_buffer(69757) := X"3C020400";
        ram_buffer(69758) := X"24630004";
        ram_buffer(69759) := X"00621024";
        ram_buffer(69760) := X"1040FF90";
        ram_buffer(69761) := X"240200FF";
        ram_buffer(69762) := X"26100001";
        ram_buffer(69763) := X"1202002E";
        ram_buffer(69764) := X"00031980";
        ram_buffer(69765) := X"00032A42";
        ram_buffer(69766) := X"321000FF";
        ram_buffer(69767) := X"1000FF96";
        ram_buffer(69768) := X"32220001";
        ram_buffer(69769) := X"1040FFD8";
        ram_buffer(69770) := X"240400FF";
        ram_buffer(69771) := X"1604FFD0";
        ram_buffer(69772) := X"2844001C";
        ram_buffer(69773) := X"1460FF83";
        ram_buffer(69774) := X"00000000";
        ram_buffer(69775) := X"02202821";
        ram_buffer(69776) := X"30A20001";
        ram_buffer(69777) := X"241000FF";
        ram_buffer(69778) := X"1000FF8B";
        ram_buffer(69779) := X"00002821";
        ram_buffer(69780) := X"14C00056";
        ram_buffer(69781) := X"2442FFFF";
        ram_buffer(69782) := X"240200FF";
        ram_buffer(69783) := X"1602FF7A";
        ram_buffer(69784) := X"000310C2";
        ram_buffer(69785) := X"1060FFF6";
        ram_buffer(69786) := X"00000000";
        ram_buffer(69787) := X"1000FF76";
        ram_buffer(69788) := X"000310C2";
        ram_buffer(69789) := X"108000D1";
        ram_buffer(69790) := X"00801821";
        ram_buffer(69791) := X"30620007";
        ram_buffer(69792) := X"1440FFD9";
        ram_buffer(69793) := X"000310C2";
        ram_buffer(69794) := X"1000FF70";
        ram_buffer(69795) := X"240300FF";
        ram_buffer(69796) := X"14400030";
        ram_buffer(69797) := X"00000000";
        ram_buffer(69798) := X"26020001";
        ram_buffer(69799) := X"304200FF";
        ram_buffer(69800) := X"28420002";
        ram_buffer(69801) := X"14400057";
        ram_buffer(69802) := X"00669023";
        ram_buffer(69803) := X"3C020400";
        ram_buffer(69804) := X"02421024";
        ram_buffer(69805) := X"10400038";
        ram_buffer(69806) := X"00000000";
        ram_buffer(69807) := X"00C39023";
        ram_buffer(69808) := X"1000FFB8";
        ram_buffer(69809) := X"00A08821";
        ram_buffer(69810) := X"32220001";
        ram_buffer(69811) := X"241000FF";
        ram_buffer(69812) := X"1000FF69";
        ram_buffer(69813) := X"00002821";
        ram_buffer(69814) := X"3C03FBFF";
        ram_buffer(69815) := X"3463FFFF";
        ram_buffer(69816) := X"02431824";
        ram_buffer(69817) := X"02028023";
        ram_buffer(69818) := X"1000FFBD";
        ram_buffer(69819) := X"32520007";
        ram_buffer(69820) := X"00008821";
        ram_buffer(69821) := X"3443FFFF";
        ram_buffer(69822) := X"00602821";
        ram_buffer(69823) := X"32220001";
        ram_buffer(69824) := X"1000FF5D";
        ram_buffer(69825) := X"241000FF";
        ram_buffer(69826) := X"14400049";
        ram_buffer(69827) := X"26040001";
        ram_buffer(69828) := X"308200FF";
        ram_buffer(69829) := X"28420002";
        ram_buffer(69830) := X"14400034";
        ram_buffer(69831) := X"240200FF";
        ram_buffer(69832) := X"1082FFC8";
        ram_buffer(69833) := X"30A20001";
        ram_buffer(69834) := X"00663021";
        ram_buffer(69835) := X"00061842";
        ram_buffer(69836) := X"30620007";
        ram_buffer(69837) := X"1440FFAC";
        ram_buffer(69838) := X"00808021";
        ram_buffer(69839) := X"1000FF7F";
        ram_buffer(69840) := X"000310C2";
        ram_buffer(69841) := X"1000FFCD";
        ram_buffer(69842) := X"00A08821";
        ram_buffer(69843) := X"1000FF8E";
        ram_buffer(69844) := X"24060001";
        ram_buffer(69845) := X"1200001D";
        ram_buffer(69846) := X"240400FF";
        ram_buffer(69847) := X"10E40056";
        ram_buffer(69848) := X"3C040400";
        ram_buffer(69849) := X"00021023";
        ram_buffer(69850) := X"00641825";
        ram_buffer(69851) := X"2844001C";
        ram_buffer(69852) := X"10800078";
        ram_buffer(69853) := X"00022023";
        ram_buffer(69854) := X"00832004";
        ram_buffer(69855) := X"00431006";
        ram_buffer(69856) := X"0004182B";
        ram_buffer(69857) := X"00431825";
        ram_buffer(69858) := X"00C31823";
        ram_buffer(69859) := X"00E08021";
        ram_buffer(69860) := X"1000FF7E";
        ram_buffer(69861) := X"00A08821";
        ram_buffer(69862) := X"1640FF82";
        ram_buffer(69863) := X"00000000";
        ram_buffer(69864) := X"00008821";
        ram_buffer(69865) := X"1000FF68";
        ram_buffer(69866) := X"00008021";
        ram_buffer(69867) := X"1040FF51";
        ram_buffer(69868) := X"240400FF";
        ram_buffer(69869) := X"1604FF48";
        ram_buffer(69870) := X"00000000";
        ram_buffer(69871) := X"1060FFA0";
        ram_buffer(69872) := X"00000000";
        ram_buffer(69873) := X"1000FF20";
        ram_buffer(69874) := X"000310C2";
        ram_buffer(69875) := X"14600036";
        ram_buffer(69876) := X"00021027";
        ram_buffer(69877) := X"240200FF";
        ram_buffer(69878) := X"10E20037";
        ram_buffer(69879) := X"00C01821";
        ram_buffer(69880) := X"00E08021";
        ram_buffer(69881) := X"1000FF17";
        ram_buffer(69882) := X"00A08821";
        ram_buffer(69883) := X"16000021";
        ram_buffer(69884) := X"00000000";
        ram_buffer(69885) := X"1460005B";
        ram_buffer(69886) := X"00000000";
        ram_buffer(69887) := X"1000FF11";
        ram_buffer(69888) := X"00C01821";
        ram_buffer(69889) := X"16000013";
        ram_buffer(69890) := X"00000000";
        ram_buffer(69891) := X"1460003E";
        ram_buffer(69892) := X"00000000";
        ram_buffer(69893) := X"10C00051";
        ram_buffer(69894) := X"00001021";
        ram_buffer(69895) := X"00C01821";
        ram_buffer(69896) := X"1000FF08";
        ram_buffer(69897) := X"00A08821";
        ram_buffer(69898) := X"1000FF32";
        ram_buffer(69899) := X"24060001";
        ram_buffer(69900) := X"16000027";
        ram_buffer(69901) := X"240400FF";
        ram_buffer(69902) := X"1460003D";
        ram_buffer(69903) := X"00021027";
        ram_buffer(69904) := X"240200FF";
        ram_buffer(69905) := X"10E2003E";
        ram_buffer(69906) := X"00C01821";
        ram_buffer(69907) := X"1000FEFD";
        ram_buffer(69908) := X"00E08021";
        ram_buffer(69909) := X"14600009";
        ram_buffer(69910) := X"00000000";
        ram_buffer(69911) := X"10C0FFA4";
        ram_buffer(69912) := X"3C02003F";
        ram_buffer(69913) := X"00C01821";
        ram_buffer(69914) := X"00A08821";
        ram_buffer(69915) := X"1000FEF5";
        ram_buffer(69916) := X"241000FF";
        ram_buffer(69917) := X"10600034";
        ram_buffer(69918) := X"00000000";
        ram_buffer(69919) := X"10C0FEF1";
        ram_buffer(69920) := X"241000FF";
        ram_buffer(69921) := X"000318C2";
        ram_buffer(69922) := X"000610C2";
        ram_buffer(69923) := X"00431025";
        ram_buffer(69924) := X"3C040040";
        ram_buffer(69925) := X"00441024";
        ram_buffer(69926) := X"14400040";
        ram_buffer(69927) := X"00000000";
        ram_buffer(69928) := X"1000FEE8";
        ram_buffer(69929) := X"000318C0";
        ram_buffer(69930) := X"1040FFB7";
        ram_buffer(69931) := X"240400FF";
        ram_buffer(69932) := X"14E4FFAF";
        ram_buffer(69933) := X"2844001C";
        ram_buffer(69934) := X"10C0FF62";
        ram_buffer(69935) := X"30A20001";
        ram_buffer(69936) := X"00C01821";
        ram_buffer(69937) := X"241000FF";
        ram_buffer(69938) := X"1000FEDE";
        ram_buffer(69939) := X"00A08821";
        ram_buffer(69940) := X"10E4001B";
        ram_buffer(69941) := X"3C040400";
        ram_buffer(69942) := X"00021023";
        ram_buffer(69943) := X"00641825";
        ram_buffer(69944) := X"2844001C";
        ram_buffer(69945) := X"10800031";
        ram_buffer(69946) := X"00022023";
        ram_buffer(69947) := X"00832004";
        ram_buffer(69948) := X"00431006";
        ram_buffer(69949) := X"0004182B";
        ram_buffer(69950) := X"00431825";
        ram_buffer(69951) := X"00661821";
        ram_buffer(69952) := X"1000FEFD";
        ram_buffer(69953) := X"00E08021";
        ram_buffer(69954) := X"10C0FECF";
        ram_buffer(69955) := X"000310C2";
        ram_buffer(69956) := X"00662023";
        ram_buffer(69957) := X"3C020400";
        ram_buffer(69958) := X"00821024";
        ram_buffer(69959) := X"1040FF55";
        ram_buffer(69960) := X"00C31823";
        ram_buffer(69961) := X"30720007";
        ram_buffer(69962) := X"1000FF2D";
        ram_buffer(69963) := X"00A08821";
        ram_buffer(69964) := X"1040FFF2";
        ram_buffer(69965) := X"240400FF";
        ram_buffer(69966) := X"14E4FFEA";
        ram_buffer(69967) := X"2844001C";
        ram_buffer(69968) := X"10C0FF40";
        ram_buffer(69969) := X"30A20001";
        ram_buffer(69970) := X"00C01821";
        ram_buffer(69971) := X"1000FEBD";
        ram_buffer(69972) := X"241000FF";
        ram_buffer(69973) := X"1000FF8C";
        ram_buffer(69974) := X"24030001";
        ram_buffer(69975) := X"1000FEFA";
        ram_buffer(69976) := X"00008821";
        ram_buffer(69977) := X"10C0FEB8";
        ram_buffer(69978) := X"000310C2";
        ram_buffer(69979) := X"00661821";
        ram_buffer(69980) := X"3C020400";
        ram_buffer(69981) := X"00621024";
        ram_buffer(69982) := X"1040FF41";
        ram_buffer(69983) := X"30620007";
        ram_buffer(69984) := X"3C04FBFF";
        ram_buffer(69985) := X"3484FFFF";
        ram_buffer(69986) := X"24100001";
        ram_buffer(69987) := X"1440FF16";
        ram_buffer(69988) := X"00641824";
        ram_buffer(69989) := X"1000FEE9";
        ram_buffer(69990) := X"000310C2";
        ram_buffer(69991) := X"3C0301FF";
        ram_buffer(69992) := X"00008821";
        ram_buffer(69993) := X"1000FEA7";
        ram_buffer(69994) := X"3463FFF8";
        ram_buffer(69995) := X"24030001";
        ram_buffer(69996) := X"00661821";
        ram_buffer(69997) := X"1000FED0";
        ram_buffer(69998) := X"00E08021";
        ram_buffer(69999) := X"1000FEE2";
        ram_buffer(70000) := X"00008821";
        ram_buffer(70001) := X"00042DC2";
        ram_buffer(70002) := X"30A500FF";
        ram_buffer(70003) := X"3C03007F";
        ram_buffer(70004) := X"3463FFFF";
        ram_buffer(70005) := X"28A2007F";
        ram_buffer(70006) := X"00641824";
        ram_buffer(70007) := X"14400011";
        ram_buffer(70008) := X"000427C2";
        ram_buffer(70009) := X"28A2009E";
        ram_buffer(70010) := X"1040000A";
        ram_buffer(70011) := X"3C060080";
        ram_buffer(70012) := X"28A20096";
        ram_buffer(70013) := X"1440000E";
        ram_buffer(70014) := X"00661825";
        ram_buffer(70015) := X"24A2FF6A";
        ram_buffer(70016) := X"00431004";
        ram_buffer(70017) := X"10800008";
        ram_buffer(70018) := X"00000000";
        ram_buffer(70019) := X"03E00008";
        ram_buffer(70020) := X"00021023";
        ram_buffer(70021) := X"3C027FFF";
        ram_buffer(70022) := X"3442FFFF";
        ram_buffer(70023) := X"03E00008";
        ram_buffer(70024) := X"00821021";
        ram_buffer(70025) := X"00001021";
        ram_buffer(70026) := X"03E00008";
        ram_buffer(70027) := X"00000000";
        ram_buffer(70028) := X"24020096";
        ram_buffer(70029) := X"00451023";
        ram_buffer(70030) := X"1000FFF2";
        ram_buffer(70031) := X"00431006";
        ram_buffer(70032) := X"27BDFFE0";
        ram_buffer(70033) := X"AFBF001C";
        ram_buffer(70034) := X"AFB10018";
        ram_buffer(70035) := X"10800047";
        ram_buffer(70036) := X"AFB00014";
        ram_buffer(70037) := X"00808021";
        ram_buffer(70038) := X"04800053";
        ram_buffer(70039) := X"00048FC2";
        ram_buffer(70040) := X"0C031D29";
        ram_buffer(70041) := X"02002021";
        ram_buffer(70042) := X"2404009E";
        ram_buffer(70043) := X"00822023";
        ram_buffer(70044) := X"28830097";
        ram_buffer(70045) := X"10600015";
        ram_buffer(70046) := X"2883009A";
        ram_buffer(70047) := X"24020096";
        ram_buffer(70048) := X"00441023";
        ram_buffer(70049) := X"00508004";
        ram_buffer(70050) := X"3C02007F";
        ram_buffer(70051) := X"3442FFFF";
        ram_buffer(70052) := X"02028024";
        ram_buffer(70053) := X"308200FF";
        ram_buffer(70054) := X"3C04007F";
        ram_buffer(70055) := X"3484FFFF";
        ram_buffer(70056) := X"02201821";
        ram_buffer(70057) := X"000215C0";
        ram_buffer(70058) := X"8FBF001C";
        ram_buffer(70059) := X"02048024";
        ram_buffer(70060) := X"02028025";
        ram_buffer(70061) := X"00031FC0";
        ram_buffer(70062) := X"02031025";
        ram_buffer(70063) := X"8FB10018";
        ram_buffer(70064) := X"8FB00014";
        ram_buffer(70065) := X"03E00008";
        ram_buffer(70066) := X"27BD0020";
        ram_buffer(70067) := X"10600040";
        ram_buffer(70068) := X"24050005";
        ram_buffer(70069) := X"24030099";
        ram_buffer(70070) := X"00641823";
        ram_buffer(70071) := X"00708004";
        ram_buffer(70072) := X"3C03FBFF";
        ram_buffer(70073) := X"3463FFFF";
        ram_buffer(70074) := X"32050007";
        ram_buffer(70075) := X"10A00006";
        ram_buffer(70076) := X"02031824";
        ram_buffer(70077) := X"3210000F";
        ram_buffer(70078) := X"24050004";
        ram_buffer(70079) := X"12050003";
        ram_buffer(70080) := X"3C050400";
        ram_buffer(70081) := X"24630004";
        ram_buffer(70082) := X"3C050400";
        ram_buffer(70083) := X"00652824";
        ram_buffer(70084) := X"10A00007";
        ram_buffer(70085) := X"00038180";
        ram_buffer(70086) := X"3C04FBFF";
        ram_buffer(70087) := X"3484FFFF";
        ram_buffer(70088) := X"00641824";
        ram_buffer(70089) := X"2404009F";
        ram_buffer(70090) := X"00822023";
        ram_buffer(70091) := X"00038180";
        ram_buffer(70092) := X"308200FF";
        ram_buffer(70093) := X"3C04007F";
        ram_buffer(70094) := X"00108242";
        ram_buffer(70095) := X"3484FFFF";
        ram_buffer(70096) := X"02201821";
        ram_buffer(70097) := X"000215C0";
        ram_buffer(70098) := X"8FBF001C";
        ram_buffer(70099) := X"02048024";
        ram_buffer(70100) := X"02028025";
        ram_buffer(70101) := X"00031FC0";
        ram_buffer(70102) := X"02031025";
        ram_buffer(70103) := X"8FB10018";
        ram_buffer(70104) := X"8FB00014";
        ram_buffer(70105) := X"03E00008";
        ram_buffer(70106) := X"27BD0020";
        ram_buffer(70107) := X"3C04007F";
        ram_buffer(70108) := X"00001021";
        ram_buffer(70109) := X"00008021";
        ram_buffer(70110) := X"3484FFFF";
        ram_buffer(70111) := X"000215C0";
        ram_buffer(70112) := X"8FBF001C";
        ram_buffer(70113) := X"00001821";
        ram_buffer(70114) := X"02048024";
        ram_buffer(70115) := X"02028025";
        ram_buffer(70116) := X"00031FC0";
        ram_buffer(70117) := X"02031025";
        ram_buffer(70118) := X"8FB10018";
        ram_buffer(70119) := X"8FB00014";
        ram_buffer(70120) := X"03E00008";
        ram_buffer(70121) := X"27BD0020";
        ram_buffer(70122) := X"00048023";
        ram_buffer(70123) := X"0C031D29";
        ram_buffer(70124) := X"02002021";
        ram_buffer(70125) := X"2404009E";
        ram_buffer(70126) := X"00822023";
        ram_buffer(70127) := X"28830097";
        ram_buffer(70128) := X"1060FFC2";
        ram_buffer(70129) := X"2883009A";
        ram_buffer(70130) := X"1000FFAD";
        ram_buffer(70131) := X"24020096";
        ram_buffer(70132) := X"240300B9";
        ram_buffer(70133) := X"00641823";
        ram_buffer(70134) := X"00701804";
        ram_buffer(70135) := X"00A22823";
        ram_buffer(70136) := X"00B08006";
        ram_buffer(70137) := X"0003182B";
        ram_buffer(70138) := X"1000FFBD";
        ram_buffer(70139) := X"02038025";
        ram_buffer(70140) := X"3C08000F";
        ram_buffer(70141) := X"3508FFFF";
        ram_buffer(70142) := X"27BDFFD8";
        ram_buffer(70143) := X"01044824";
        ram_buffer(70144) := X"01064024";
        ram_buffer(70145) := X"00041502";
        ram_buffer(70146) := X"00056742";
        ram_buffer(70147) := X"00075742";
        ram_buffer(70148) := X"AFB10018";
        ram_buffer(70149) := X"000948C0";
        ram_buffer(70150) := X"00065D02";
        ram_buffer(70151) := X"000840C0";
        ram_buffer(70152) := X"00048FC2";
        ram_buffer(70153) := X"000627C2";
        ram_buffer(70154) := X"AFB00014";
        ram_buffer(70155) := X"AFBF0024";
        ram_buffer(70156) := X"305007FF";
        ram_buffer(70157) := X"AFB30020";
        ram_buffer(70158) := X"AFB2001C";
        ram_buffer(70159) := X"012C1025";
        ram_buffer(70160) := X"000528C0";
        ram_buffer(70161) := X"316607FF";
        ram_buffer(70162) := X"010A4025";
        ram_buffer(70163) := X"12240061";
        ram_buffer(70164) := X"000738C0";
        ram_buffer(70165) := X"02064823";
        ram_buffer(70166) := X"192000CE";
        ram_buffer(70167) := X"00000000";
        ram_buffer(70168) := X"14C0000B";
        ram_buffer(70169) := X"240307FF";
        ram_buffer(70170) := X"01071825";
        ram_buffer(70171) := X"1060007F";
        ram_buffer(70172) := X"240307FF";
        ram_buffer(70173) := X"2529FFFF";
        ram_buffer(70174) := X"1520010A";
        ram_buffer(70175) := X"00A79023";
        ram_buffer(70176) := X"00481023";
        ram_buffer(70177) := X"00B2282B";
        ram_buffer(70178) := X"10000015";
        ram_buffer(70179) := X"00451023";
        ram_buffer(70180) := X"120300A6";
        ram_buffer(70181) := X"3C030080";
        ram_buffer(70182) := X"01034025";
        ram_buffer(70183) := X"29230039";
        ram_buffer(70184) := X"106000E5";
        ram_buffer(70185) := X"29230020";
        ram_buffer(70186) := X"1060010D";
        ram_buffer(70187) := X"24040020";
        ram_buffer(70188) := X"00892023";
        ram_buffer(70189) := X"00881804";
        ram_buffer(70190) := X"01279006";
        ram_buffer(70191) := X"00873804";
        ram_buffer(70192) := X"00721825";
        ram_buffer(70193) := X"0007382B";
        ram_buffer(70194) := X"00673825";
        ram_buffer(70195) := X"01284006";
        ram_buffer(70196) := X"00A79023";
        ram_buffer(70197) := X"00484023";
        ram_buffer(70198) := X"00B2282B";
        ram_buffer(70199) := X"01051023";
        ram_buffer(70200) := X"3C130080";
        ram_buffer(70201) := X"00531824";
        ram_buffer(70202) := X"106000A6";
        ram_buffer(70203) := X"32430007";
        ram_buffer(70204) := X"2673FFFF";
        ram_buffer(70205) := X"00539824";
        ram_buffer(70206) := X"126000B9";
        ram_buffer(70207) := X"00000000";
        ram_buffer(70208) := X"0C031D29";
        ram_buffer(70209) := X"02602021";
        ram_buffer(70210) := X"2446FFF8";
        ram_buffer(70211) := X"28C30020";
        ram_buffer(70212) := X"106000BB";
        ram_buffer(70213) := X"2442FFD8";
        ram_buffer(70214) := X"00061823";
        ram_buffer(70215) := X"00721806";
        ram_buffer(70216) := X"00D31004";
        ram_buffer(70217) := X"00629825";
        ram_buffer(70218) := X"00D0102A";
        ram_buffer(70219) := X"144000B8";
        ram_buffer(70220) := X"00D29004";
        ram_buffer(70221) := X"00D03023";
        ram_buffer(70222) := X"24C20001";
        ram_buffer(70223) := X"28430020";
        ram_buffer(70224) := X"106000DC";
        ram_buffer(70225) := X"24030020";
        ram_buffer(70226) := X"24040020";
        ram_buffer(70227) := X"00822023";
        ram_buffer(70228) := X"00521806";
        ram_buffer(70229) := X"00923804";
        ram_buffer(70230) := X"00932004";
        ram_buffer(70231) := X"00832025";
        ram_buffer(70232) := X"0007382B";
        ram_buffer(70233) := X"00879025";
        ram_buffer(70234) := X"00531006";
        ram_buffer(70235) := X"32430007";
        ram_buffer(70236) := X"00008021";
        ram_buffer(70237) := X"10600041";
        ram_buffer(70238) := X"3C030080";
        ram_buffer(70239) := X"3243000F";
        ram_buffer(70240) := X"24040004";
        ram_buffer(70241) := X"1064003C";
        ram_buffer(70242) := X"26440004";
        ram_buffer(70243) := X"0092382B";
        ram_buffer(70244) := X"00471021";
        ram_buffer(70245) := X"3C030080";
        ram_buffer(70246) := X"00431824";
        ram_buffer(70247) := X"1460003A";
        ram_buffer(70248) := X"00809021";
        ram_buffer(70249) := X"00021F40";
        ram_buffer(70250) := X"001238C2";
        ram_buffer(70251) := X"00E33825";
        ram_buffer(70252) := X"000218C2";
        ram_buffer(70253) := X"240207FF";
        ram_buffer(70254) := X"12020060";
        ram_buffer(70255) := X"00000000";
        ram_buffer(70256) := X"3C06000F";
        ram_buffer(70257) := X"34C6FFFF";
        ram_buffer(70258) := X"00662824";
        ram_buffer(70259) := X"1000003B";
        ram_buffer(70260) := X"320207FF";
        ram_buffer(70261) := X"02062023";
        ram_buffer(70262) := X"1880009E";
        ram_buffer(70263) := X"00000000";
        ram_buffer(70264) := X"10C00047";
        ram_buffer(70265) := X"01071825";
        ram_buffer(70266) := X"240307FF";
        ram_buffer(70267) := X"1203004F";
        ram_buffer(70268) := X"3C030080";
        ram_buffer(70269) := X"01034025";
        ram_buffer(70270) := X"28830039";
        ram_buffer(70271) := X"146000E2";
        ram_buffer(70272) := X"28830020";
        ram_buffer(70273) := X"01073825";
        ram_buffer(70274) := X"0007382B";
        ram_buffer(70275) := X"00004021";
        ram_buffer(70276) := X"00E59021";
        ram_buffer(70277) := X"01024021";
        ram_buffer(70278) := X"0245282B";
        ram_buffer(70279) := X"00A81021";
        ram_buffer(70280) := X"3C030080";
        ram_buffer(70281) := X"00431824";
        ram_buffer(70282) := X"10600056";
        ram_buffer(70283) := X"32430007";
        ram_buffer(70284) := X"26100001";
        ram_buffer(70285) := X"240307FF";
        ram_buffer(70286) := X"120300FB";
        ram_buffer(70287) := X"00000000";
        ram_buffer(70288) := X"3C03FF7F";
        ram_buffer(70289) := X"3463FFFF";
        ram_buffer(70290) := X"00431024";
        ram_buffer(70291) := X"32470001";
        ram_buffer(70292) := X"00122042";
        ram_buffer(70293) := X"00879025";
        ram_buffer(70294) := X"00023FC0";
        ram_buffer(70295) := X"00F29025";
        ram_buffer(70296) := X"00021042";
        ram_buffer(70297) := X"1000FFC3";
        ram_buffer(70298) := X"32430007";
        ram_buffer(70299) := X"12030030";
        ram_buffer(70300) := X"00451825";
        ram_buffer(70301) := X"00A09021";
        ram_buffer(70302) := X"3C030080";
        ram_buffer(70303) := X"00431824";
        ram_buffer(70304) := X"1060FFC9";
        ram_buffer(70305) := X"00021F40";
        ram_buffer(70306) := X"26060001";
        ram_buffer(70307) := X"240307FF";
        ram_buffer(70308) := X"10C30065";
        ram_buffer(70309) := X"00000000";
        ram_buffer(70310) := X"3C05FF7F";
        ram_buffer(70311) := X"34A5FFFF";
        ram_buffer(70312) := X"00451024";
        ram_buffer(70313) := X"00022F40";
        ram_buffer(70314) := X"001238C2";
        ram_buffer(70315) := X"00021240";
        ram_buffer(70316) := X"00A73825";
        ram_buffer(70317) := X"00022B02";
        ram_buffer(70318) := X"30C207FF";
        ram_buffer(70319) := X"00023500";
        ram_buffer(70320) := X"3C02000F";
        ram_buffer(70321) := X"3442FFFF";
        ram_buffer(70322) := X"00A21024";
        ram_buffer(70323) := X"00111FC0";
        ram_buffer(70324) := X"00461025";
        ram_buffer(70325) := X"00431825";
        ram_buffer(70326) := X"8FBF0024";
        ram_buffer(70327) := X"00602021";
        ram_buffer(70328) := X"8FB30020";
        ram_buffer(70329) := X"8FB2001C";
        ram_buffer(70330) := X"8FB10018";
        ram_buffer(70331) := X"8FB00014";
        ram_buffer(70332) := X"00E01821";
        ram_buffer(70333) := X"00801021";
        ram_buffer(70334) := X"03E00008";
        ram_buffer(70335) := X"27BD0028";
        ram_buffer(70336) := X"1060FFDA";
        ram_buffer(70337) := X"240307FF";
        ram_buffer(70338) := X"2484FFFF";
        ram_buffer(70339) := X"14800005";
        ram_buffer(70340) := X"00A79021";
        ram_buffer(70341) := X"00481021";
        ram_buffer(70342) := X"0245282B";
        ram_buffer(70343) := X"1000FFC0";
        ram_buffer(70344) := X"00A21021";
        ram_buffer(70345) := X"1603FFB5";
        ram_buffer(70346) := X"28830039";
        ram_buffer(70347) := X"00451825";
        ram_buffer(70348) := X"1460FFD1";
        ram_buffer(70349) := X"00A09021";
        ram_buffer(70350) := X"00003821";
        ram_buffer(70351) := X"00671025";
        ram_buffer(70352) := X"1040003A";
        ram_buffer(70353) := X"240207FF";
        ram_buffer(70354) := X"3C050007";
        ram_buffer(70355) := X"34A5FFFF";
        ram_buffer(70356) := X"00651024";
        ram_buffer(70357) := X"00471825";
        ram_buffer(70358) := X"1460003B";
        ram_buffer(70359) := X"00000000";
        ram_buffer(70360) := X"00008821";
        ram_buffer(70361) := X"240207FF";
        ram_buffer(70362) := X"1000FFD4";
        ram_buffer(70363) := X"2407FFFF";
        ram_buffer(70364) := X"02461825";
        ram_buffer(70365) := X"10600129";
        ram_buffer(70366) := X"00003821";
        ram_buffer(70367) := X"00C01021";
        ram_buffer(70368) := X"32430007";
        ram_buffer(70369) := X"1460FF7D";
        ram_buffer(70370) := X"00021F40";
        ram_buffer(70371) := X"1000FF87";
        ram_buffer(70372) := X"001238C2";
        ram_buffer(70373) := X"1520005B";
        ram_buffer(70374) := X"26030001";
        ram_buffer(70375) := X"306307FF";
        ram_buffer(70376) := X"28630002";
        ram_buffer(70377) := X"14600097";
        ram_buffer(70378) := X"00A79023";
        ram_buffer(70379) := X"00B2182B";
        ram_buffer(70380) := X"00489823";
        ram_buffer(70381) := X"02639823";
        ram_buffer(70382) := X"3C030080";
        ram_buffer(70383) := X"02631824";
        ram_buffer(70384) := X"1060006C";
        ram_buffer(70385) := X"02531825";
        ram_buffer(70386) := X"00E59023";
        ram_buffer(70387) := X"01021023";
        ram_buffer(70388) := X"00F2382B";
        ram_buffer(70389) := X"00479823";
        ram_buffer(70390) := X"1660FF49";
        ram_buffer(70391) := X"00808821";
        ram_buffer(70392) := X"0C031D29";
        ram_buffer(70393) := X"02402021";
        ram_buffer(70394) := X"24420020";
        ram_buffer(70395) := X"2446FFF8";
        ram_buffer(70396) := X"28C30020";
        ram_buffer(70397) := X"1460FF49";
        ram_buffer(70398) := X"00061823";
        ram_buffer(70399) := X"2442FFD8";
        ram_buffer(70400) := X"00529804";
        ram_buffer(70401) := X"00D0102A";
        ram_buffer(70402) := X"1040FF4A";
        ram_buffer(70403) := X"00009021";
        ram_buffer(70404) := X"3C02FF7F";
        ram_buffer(70405) := X"3442FFFF";
        ram_buffer(70406) := X"02068023";
        ram_buffer(70407) := X"02621024";
        ram_buffer(70408) := X"1000FF54";
        ram_buffer(70409) := X"32430007";
        ram_buffer(70410) := X"240207FF";
        ram_buffer(70411) := X"00002821";
        ram_buffer(70412) := X"1000FFA2";
        ram_buffer(70413) := X"00003821";
        ram_buffer(70414) := X"01073825";
        ram_buffer(70415) := X"0007382B";
        ram_buffer(70416) := X"1000FF23";
        ram_buffer(70417) := X"00004021";
        ram_buffer(70418) := X"00402821";
        ram_buffer(70419) := X"1000FF9B";
        ram_buffer(70420) := X"240207FF";
        ram_buffer(70421) := X"14800080";
        ram_buffer(70422) := X"00000000";
        ram_buffer(70423) := X"26040001";
        ram_buffer(70424) := X"308307FF";
        ram_buffer(70425) := X"28630002";
        ram_buffer(70426) := X"1460005F";
        ram_buffer(70427) := X"00000000";
        ram_buffer(70428) := X"240307FF";
        ram_buffer(70429) := X"1083006C";
        ram_buffer(70430) := X"00481021";
        ram_buffer(70431) := X"00A73821";
        ram_buffer(70432) := X"00E5282B";
        ram_buffer(70433) := X"00A21021";
        ram_buffer(70434) := X"000297C0";
        ram_buffer(70435) := X"00073842";
        ram_buffer(70436) := X"02479025";
        ram_buffer(70437) := X"00021042";
        ram_buffer(70438) := X"32430007";
        ram_buffer(70439) := X"1000FF35";
        ram_buffer(70440) := X"00808021";
        ram_buffer(70441) := X"1603FEFD";
        ram_buffer(70442) := X"00451825";
        ram_buffer(70443) := X"1000FFA0";
        ram_buffer(70444) := X"00000000";
        ram_buffer(70445) := X"24C6FFE1";
        ram_buffer(70446) := X"10430047";
        ram_buffer(70447) := X"00D33006";
        ram_buffer(70448) := X"00023823";
        ram_buffer(70449) := X"00F33804";
        ram_buffer(70450) := X"02473825";
        ram_buffer(70451) := X"0007382B";
        ram_buffer(70452) := X"00C79025";
        ram_buffer(70453) := X"00001021";
        ram_buffer(70454) := X"1000FFA9";
        ram_buffer(70455) := X"00008021";
        ram_buffer(70456) := X"1124003F";
        ram_buffer(70457) := X"01281806";
        ram_buffer(70458) := X"00094823";
        ram_buffer(70459) := X"01284004";
        ram_buffer(70460) := X"01073825";
        ram_buffer(70461) := X"0007382B";
        ram_buffer(70462) := X"00673825";
        ram_buffer(70463) := X"1000FEF4";
        ram_buffer(70464) := X"00004021";
        ram_buffer(70465) := X"1200002B";
        ram_buffer(70466) := X"00451825";
        ram_buffer(70467) := X"240307FF";
        ram_buffer(70468) := X"10C300B8";
        ram_buffer(70469) := X"3C030080";
        ram_buffer(70470) := X"00094823";
        ram_buffer(70471) := X"00431025";
        ram_buffer(70472) := X"29230039";
        ram_buffer(70473) := X"10600071";
        ram_buffer(70474) := X"29230020";
        ram_buffer(70475) := X"106000BD";
        ram_buffer(70476) := X"24030020";
        ram_buffer(70477) := X"240A0020";
        ram_buffer(70478) := X"01495023";
        ram_buffer(70479) := X"01259006";
        ram_buffer(70480) := X"01421804";
        ram_buffer(70481) := X"01452804";
        ram_buffer(70482) := X"00721825";
        ram_buffer(70483) := X"0005902B";
        ram_buffer(70484) := X"00729025";
        ram_buffer(70485) := X"01224806";
        ram_buffer(70486) := X"00F29023";
        ram_buffer(70487) := X"01094823";
        ram_buffer(70488) := X"00F2382B";
        ram_buffer(70489) := X"01271023";
        ram_buffer(70490) := X"00C08021";
        ram_buffer(70491) := X"1000FEDC";
        ram_buffer(70492) := X"00808821";
        ram_buffer(70493) := X"1460FEE0";
        ram_buffer(70494) := X"00003821";
        ram_buffer(70495) := X"00008821";
        ram_buffer(70496) := X"1000FF0F";
        ram_buffer(70497) := X"00008021";
        ram_buffer(70498) := X"1060002A";
        ram_buffer(70499) := X"24060020";
        ram_buffer(70500) := X"00C43023";
        ram_buffer(70501) := X"00C81804";
        ram_buffer(70502) := X"00879006";
        ram_buffer(70503) := X"00C73804";
        ram_buffer(70504) := X"00721825";
        ram_buffer(70505) := X"0007382B";
        ram_buffer(70506) := X"00673825";
        ram_buffer(70507) := X"1000FF18";
        ram_buffer(70508) := X"00884006";
        ram_buffer(70509) := X"14600043";
        ram_buffer(70510) := X"00000000";
        ram_buffer(70511) := X"240207FF";
        ram_buffer(70512) := X"10C2008C";
        ram_buffer(70513) := X"01001021";
        ram_buffer(70514) := X"00E09021";
        ram_buffer(70515) := X"00C08021";
        ram_buffer(70516) := X"1000FF29";
        ram_buffer(70517) := X"00808821";
        ram_buffer(70518) := X"1000FFBB";
        ram_buffer(70519) := X"00003821";
        ram_buffer(70520) := X"1000FFC3";
        ram_buffer(70521) := X"00004021";
        ram_buffer(70522) := X"1600006C";
        ram_buffer(70523) := X"00451825";
        ram_buffer(70524) := X"146000A6";
        ram_buffer(70525) := X"01071825";
        ram_buffer(70526) := X"01001021";
        ram_buffer(70527) := X"1000FF1E";
        ram_buffer(70528) := X"00E09021";
        ram_buffer(70529) := X"1600001F";
        ram_buffer(70530) := X"00451825";
        ram_buffer(70531) := X"14600053";
        ram_buffer(70532) := X"01071825";
        ram_buffer(70533) := X"10600080";
        ram_buffer(70534) := X"00E09021";
        ram_buffer(70535) := X"01001021";
        ram_buffer(70536) := X"1000FF15";
        ram_buffer(70537) := X"00808821";
        ram_buffer(70538) := X"00001821";
        ram_buffer(70539) := X"1000FF43";
        ram_buffer(70540) := X"00003821";
        ram_buffer(70541) := X"10860076";
        ram_buffer(70542) := X"00881806";
        ram_buffer(70543) := X"00042023";
        ram_buffer(70544) := X"00884004";
        ram_buffer(70545) := X"01073825";
        ram_buffer(70546) := X"0007382B";
        ram_buffer(70547) := X"00673825";
        ram_buffer(70548) := X"1000FEEF";
        ram_buffer(70549) := X"00004021";
        ram_buffer(70550) := X"16000028";
        ram_buffer(70551) := X"240307FF";
        ram_buffer(70552) := X"00451825";
        ram_buffer(70553) := X"14600078";
        ram_buffer(70554) := X"00000000";
        ram_buffer(70555) := X"240207FF";
        ram_buffer(70556) := X"10C200A0";
        ram_buffer(70557) := X"01001021";
        ram_buffer(70558) := X"00E09021";
        ram_buffer(70559) := X"1000FEFE";
        ram_buffer(70560) := X"00C08021";
        ram_buffer(70561) := X"14600009";
        ram_buffer(70562) := X"00000000";
        ram_buffer(70563) := X"01071025";
        ram_buffer(70564) := X"10400076";
        ram_buffer(70565) := X"3C030007";
        ram_buffer(70566) := X"01001021";
        ram_buffer(70567) := X"00E09021";
        ram_buffer(70568) := X"00808821";
        ram_buffer(70569) := X"1000FEF4";
        ram_buffer(70570) := X"241007FF";
        ram_buffer(70571) := X"01073825";
        ram_buffer(70572) := X"14E00040";
        ram_buffer(70573) := X"000220C2";
        ram_buffer(70574) := X"00A09021";
        ram_buffer(70575) := X"1000FEEE";
        ram_buffer(70576) := X"241007FF";
        ram_buffer(70577) := X"00094827";
        ram_buffer(70578) := X"15200048";
        ram_buffer(70579) := X"240307FF";
        ram_buffer(70580) := X"00E59023";
        ram_buffer(70581) := X"01021023";
        ram_buffer(70582) := X"00F2382B";
        ram_buffer(70583) := X"00471023";
        ram_buffer(70584) := X"00C08021";
        ram_buffer(70585) := X"1000FE7E";
        ram_buffer(70586) := X"00808821";
        ram_buffer(70587) := X"00452825";
        ram_buffer(70588) := X"0005902B";
        ram_buffer(70589) := X"1000FF98";
        ram_buffer(70590) := X"00004821";
        ram_buffer(70591) := X"10C3007D";
        ram_buffer(70592) := X"3C030080";
        ram_buffer(70593) := X"00042023";
        ram_buffer(70594) := X"00431025";
        ram_buffer(70595) := X"28830039";
        ram_buffer(70596) := X"1060005A";
        ram_buffer(70597) := X"28830020";
        ram_buffer(70598) := X"1060007B";
        ram_buffer(70599) := X"24030020";
        ram_buffer(70600) := X"24090020";
        ram_buffer(70601) := X"01244823";
        ram_buffer(70602) := X"00859006";
        ram_buffer(70603) := X"01221804";
        ram_buffer(70604) := X"01252804";
        ram_buffer(70605) := X"00721825";
        ram_buffer(70606) := X"0005902B";
        ram_buffer(70607) := X"00729025";
        ram_buffer(70608) := X"00821006";
        ram_buffer(70609) := X"02479021";
        ram_buffer(70610) := X"00484021";
        ram_buffer(70611) := X"0247382B";
        ram_buffer(70612) := X"00E81021";
        ram_buffer(70613) := X"1000FEB2";
        ram_buffer(70614) := X"00C08021";
        ram_buffer(70615) := X"1060FEC6";
        ram_buffer(70616) := X"00A09021";
        ram_buffer(70617) := X"00A79023";
        ram_buffer(70618) := X"00481823";
        ram_buffer(70619) := X"00B2302B";
        ram_buffer(70620) := X"00663023";
        ram_buffer(70621) := X"3C030080";
        ram_buffer(70622) := X"00C31824";
        ram_buffer(70623) := X"1060FEFC";
        ram_buffer(70624) := X"01021023";
        ram_buffer(70625) := X"00E59023";
        ram_buffer(70626) := X"00F2382B";
        ram_buffer(70627) := X"00471023";
        ram_buffer(70628) := X"32430007";
        ram_buffer(70629) := X"1000FE77";
        ram_buffer(70630) := X"00808821";
        ram_buffer(70631) := X"1460FFC3";
        ram_buffer(70632) := X"00000000";
        ram_buffer(70633) := X"01001021";
        ram_buffer(70634) := X"00E09021";
        ram_buffer(70635) := X"1000FEB2";
        ram_buffer(70636) := X"241007FF";
        ram_buffer(70637) := X"000818C2";
        ram_buffer(70638) := X"00641825";
        ram_buffer(70639) := X"3C060008";
        ram_buffer(70640) := X"00661824";
        ram_buffer(70641) := X"14600040";
        ram_buffer(70642) := X"000528C2";
        ram_buffer(70643) := X"00021740";
        ram_buffer(70644) := X"00453825";
        ram_buffer(70645) := X"000420C0";
        ram_buffer(70646) := X"00071742";
        ram_buffer(70647) := X"00441025";
        ram_buffer(70648) := X"000790C0";
        ram_buffer(70649) := X"1000FEA4";
        ram_buffer(70650) := X"241007FF";
        ram_buffer(70651) := X"14C3FF4D";
        ram_buffer(70652) := X"29230039";
        ram_buffer(70653) := X"01071825";
        ram_buffer(70654) := X"10600039";
        ram_buffer(70655) := X"01001021";
        ram_buffer(70656) := X"00E09021";
        ram_buffer(70657) := X"241007FF";
        ram_buffer(70658) := X"1000FE9B";
        ram_buffer(70659) := X"00808821";
        ram_buffer(70660) := X"1000FF8C";
        ram_buffer(70661) := X"00004021";
        ram_buffer(70662) := X"00003821";
        ram_buffer(70663) := X"1000FE68";
        ram_buffer(70664) := X"00008821";
        ram_buffer(70665) := X"11230041";
        ram_buffer(70666) := X"01229006";
        ram_buffer(70667) := X"00094823";
        ram_buffer(70668) := X"01221804";
        ram_buffer(70669) := X"00652825";
        ram_buffer(70670) := X"0005182B";
        ram_buffer(70671) := X"02439025";
        ram_buffer(70672) := X"1000FF45";
        ram_buffer(70673) := X"00004821";
        ram_buffer(70674) := X"00042027";
        ram_buffer(70675) := X"14800027";
        ram_buffer(70676) := X"240307FF";
        ram_buffer(70677) := X"00A79021";
        ram_buffer(70678) := X"00481021";
        ram_buffer(70679) := X"0247382B";
        ram_buffer(70680) := X"00E21021";
        ram_buffer(70681) := X"1000FE6E";
        ram_buffer(70682) := X"00C08021";
        ram_buffer(70683) := X"3463FFFF";
        ram_buffer(70684) := X"2407FFFF";
        ram_buffer(70685) := X"1000FEB1";
        ram_buffer(70686) := X"00008821";
        ram_buffer(70687) := X"00451025";
        ram_buffer(70688) := X"0002902B";
        ram_buffer(70689) := X"1000FFAF";
        ram_buffer(70690) := X"00001021";
        ram_buffer(70691) := X"1060FE7A";
        ram_buffer(70692) := X"00A09021";
        ram_buffer(70693) := X"00A79021";
        ram_buffer(70694) := X"00481021";
        ram_buffer(70695) := X"0245282B";
        ram_buffer(70696) := X"00A21021";
        ram_buffer(70697) := X"3C030080";
        ram_buffer(70698) := X"00431824";
        ram_buffer(70699) := X"1060FEB4";
        ram_buffer(70700) := X"3C03FF7F";
        ram_buffer(70701) := X"3463FFFF";
        ram_buffer(70702) := X"00431024";
        ram_buffer(70703) := X"24100001";
        ram_buffer(70704) := X"1000FE2C";
        ram_buffer(70705) := X"32430007";
        ram_buffer(70706) := X"3C02003F";
        ram_buffer(70707) := X"00008821";
        ram_buffer(70708) := X"241007FF";
        ram_buffer(70709) := X"3442FFFF";
        ram_buffer(70710) := X"1000FE32";
        ram_buffer(70711) := X"2412FFF8";
        ram_buffer(70712) := X"00003821";
        ram_buffer(70713) := X"1000FE95";
        ram_buffer(70714) := X"00808821";
        ram_buffer(70715) := X"14C3FF88";
        ram_buffer(70716) := X"28830039";
        ram_buffer(70717) := X"01071825";
        ram_buffer(70718) := X"1460FFAB";
        ram_buffer(70719) := X"01001021";
        ram_buffer(70720) := X"1000FE8E";
        ram_buffer(70721) := X"00003821";
        ram_buffer(70722) := X"1083000A";
        ram_buffer(70723) := X"00829006";
        ram_buffer(70724) := X"00042023";
        ram_buffer(70725) := X"00821004";
        ram_buffer(70726) := X"00452825";
        ram_buffer(70727) := X"0005102B";
        ram_buffer(70728) := X"02429025";
        ram_buffer(70729) := X"1000FF87";
        ram_buffer(70730) := X"00001021";
        ram_buffer(70731) := X"1000FFC1";
        ram_buffer(70732) := X"00001821";
        ram_buffer(70733) := X"1000FFF8";
        ram_buffer(70734) := X"00001021";
        ram_buffer(70735) := X"27BDFFB8";
        ram_buffer(70736) := X"AFB50034";
        ram_buffer(70737) := X"AFB00020";
        ram_buffer(70738) := X"0004AD02";
        ram_buffer(70739) := X"3C10000F";
        ram_buffer(70740) := X"AFB40030";
        ram_buffer(70741) := X"3610FFFF";
        ram_buffer(70742) := X"0004A7C2";
        ram_buffer(70743) := X"32B507FF";
        ram_buffer(70744) := X"AFB7003C";
        ram_buffer(70745) := X"AFBF0044";
        ram_buffer(70746) := X"AFBE0040";
        ram_buffer(70747) := X"AFB60038";
        ram_buffer(70748) := X"AFB3002C";
        ram_buffer(70749) := X"AFB20028";
        ram_buffer(70750) := X"AFB10024";
        ram_buffer(70751) := X"02048024";
        ram_buffer(70752) := X"12A00079";
        ram_buffer(70753) := X"0280B821";
        ram_buffer(70754) := X"240207FF";
        ram_buffer(70755) := X"12A20026";
        ram_buffer(70756) := X"02051025";
        ram_buffer(70757) := X"3C040010";
        ram_buffer(70758) := X"02048025";
        ram_buffer(70759) := X"001080C0";
        ram_buffer(70760) := X"00052742";
        ram_buffer(70761) := X"00908025";
        ram_buffer(70762) := X"000590C0";
        ram_buffer(70763) := X"26B5FC01";
        ram_buffer(70764) := X"00009821";
        ram_buffer(70765) := X"0000F021";
        ram_buffer(70766) := X"00062502";
        ram_buffer(70767) := X"3C11000F";
        ram_buffer(70768) := X"3631FFFF";
        ram_buffer(70769) := X"308407FF";
        ram_buffer(70770) := X"00E01821";
        ram_buffer(70771) := X"02268824";
        ram_buffer(70772) := X"10800023";
        ram_buffer(70773) := X"0006B7C2";
        ram_buffer(70774) := X"240207FF";
        ram_buffer(70775) := X"1082007D";
        ram_buffer(70776) := X"3C020010";
        ram_buffer(70777) := X"02228825";
        ram_buffer(70778) := X"001188C0";
        ram_buffer(70779) := X"00071742";
        ram_buffer(70780) := X"00518825";
        ram_buffer(70781) := X"000718C0";
        ram_buffer(70782) := X"2484FC01";
        ram_buffer(70783) := X"00001021";
        ram_buffer(70784) := X"00533825";
        ram_buffer(70785) := X"00074080";
        ram_buffer(70786) := X"3C07100D";
        ram_buffer(70787) := X"24E7B5E0";
        ram_buffer(70788) := X"00E83821";
        ram_buffer(70789) := X"8CE60000";
        ram_buffer(70790) := X"02962826";
        ram_buffer(70791) := X"00A03821";
        ram_buffer(70792) := X"00C00008";
        ram_buffer(70793) := X"02A4A823";
        ram_buffer(70794) := X"1440007A";
        ram_buffer(70795) := X"00A09021";
        ram_buffer(70796) := X"00062502";
        ram_buffer(70797) := X"3C11000F";
        ram_buffer(70798) := X"3631FFFF";
        ram_buffer(70799) := X"308407FF";
        ram_buffer(70800) := X"24130008";
        ram_buffer(70801) := X"00008021";
        ram_buffer(70802) := X"00009021";
        ram_buffer(70803) := X"241E0002";
        ram_buffer(70804) := X"00E01821";
        ram_buffer(70805) := X"02268824";
        ram_buffer(70806) := X"1480FFDF";
        ram_buffer(70807) := X"0006B7C2";
        ram_buffer(70808) := X"02271025";
        ram_buffer(70809) := X"10400062";
        ram_buffer(70810) := X"00001821";
        ram_buffer(70811) := X"12200093";
        ram_buffer(70812) := X"00E02021";
        ram_buffer(70813) := X"02202021";
        ram_buffer(70814) := X"0C031D29";
        ram_buffer(70815) := X"AFA70010";
        ram_buffer(70816) := X"8FA70010";
        ram_buffer(70817) := X"2444FFF5";
        ram_buffer(70818) := X"2883001D";
        ram_buffer(70819) := X"10600087";
        ram_buffer(70820) := X"2405001D";
        ram_buffer(70821) := X"2443FFF8";
        ram_buffer(70822) := X"00A42823";
        ram_buffer(70823) := X"00718804";
        ram_buffer(70824) := X"00A72806";
        ram_buffer(70825) := X"00B18825";
        ram_buffer(70826) := X"00671804";
        ram_buffer(70827) := X"2402FC02";
        ram_buffer(70828) := X"00442023";
        ram_buffer(70829) := X"1000FFD2";
        ram_buffer(70830) := X"00001021";
        ram_buffer(70831) := X"02E03821";
        ram_buffer(70832) := X"30E50001";
        ram_buffer(70833) := X"240307FF";
        ram_buffer(70834) := X"00002021";
        ram_buffer(70835) := X"00009021";
        ram_buffer(70836) := X"3C10000F";
        ram_buffer(70837) := X"3610FFFF";
        ram_buffer(70838) := X"00031D00";
        ram_buffer(70839) := X"00908024";
        ram_buffer(70840) := X"02038025";
        ram_buffer(70841) := X"00052FC0";
        ram_buffer(70842) := X"02051825";
        ram_buffer(70843) := X"8FBF0044";
        ram_buffer(70844) := X"00602021";
        ram_buffer(70845) := X"8FBE0040";
        ram_buffer(70846) := X"02401821";
        ram_buffer(70847) := X"8FB7003C";
        ram_buffer(70848) := X"8FB60038";
        ram_buffer(70849) := X"8FB50034";
        ram_buffer(70850) := X"8FB40030";
        ram_buffer(70851) := X"8FB3002C";
        ram_buffer(70852) := X"8FB20028";
        ram_buffer(70853) := X"8FB10024";
        ram_buffer(70854) := X"8FB00020";
        ram_buffer(70855) := X"00801021";
        ram_buffer(70856) := X"03E00008";
        ram_buffer(70857) := X"27BD0048";
        ram_buffer(70858) := X"02C0B821";
        ram_buffer(70859) := X"02208021";
        ram_buffer(70860) := X"00609021";
        ram_buffer(70861) := X"0040F021";
        ram_buffer(70862) := X"24020002";
        ram_buffer(70863) := X"13C2FFDF";
        ram_buffer(70864) := X"24020003";
        ram_buffer(70865) := X"13C201A9";
        ram_buffer(70866) := X"3C040007";
        ram_buffer(70867) := X"24020001";
        ram_buffer(70868) := X"17C20108";
        ram_buffer(70869) := X"02E02821";
        ram_buffer(70870) := X"00001821";
        ram_buffer(70871) := X"00002021";
        ram_buffer(70872) := X"1000FFDB";
        ram_buffer(70873) := X"00009021";
        ram_buffer(70874) := X"02051025";
        ram_buffer(70875) := X"10400025";
        ram_buffer(70876) := X"24130004";
        ram_buffer(70877) := X"AFA70018";
        ram_buffer(70878) := X"12000059";
        ram_buffer(70879) := X"AFA60014";
        ram_buffer(70880) := X"02002021";
        ram_buffer(70881) := X"0C031D29";
        ram_buffer(70882) := X"AFA50010";
        ram_buffer(70883) := X"8FA50010";
        ram_buffer(70884) := X"8FA60014";
        ram_buffer(70885) := X"8FA70018";
        ram_buffer(70886) := X"2443FFF5";
        ram_buffer(70887) := X"2864001D";
        ram_buffer(70888) := X"1080004B";
        ram_buffer(70889) := X"2408001D";
        ram_buffer(70890) := X"2452FFF8";
        ram_buffer(70891) := X"01034023";
        ram_buffer(70892) := X"02508004";
        ram_buffer(70893) := X"01054006";
        ram_buffer(70894) := X"01108025";
        ram_buffer(70895) := X"02459004";
        ram_buffer(70896) := X"2415FC02";
        ram_buffer(70897) := X"02A3A823";
        ram_buffer(70898) := X"00009821";
        ram_buffer(70899) := X"1000FF7A";
        ram_buffer(70900) := X"0000F021";
        ram_buffer(70901) := X"02273825";
        ram_buffer(70902) := X"14E00008";
        ram_buffer(70903) := X"00000000";
        ram_buffer(70904) := X"00008821";
        ram_buffer(70905) := X"00001821";
        ram_buffer(70906) := X"1000FF85";
        ram_buffer(70907) := X"24020002";
        ram_buffer(70908) := X"00008821";
        ram_buffer(70909) := X"1000FF82";
        ram_buffer(70910) := X"24020001";
        ram_buffer(70911) := X"1000FF80";
        ram_buffer(70912) := X"24020003";
        ram_buffer(70913) := X"00008021";
        ram_buffer(70914) := X"00009021";
        ram_buffer(70915) := X"1000FF6A";
        ram_buffer(70916) := X"241E0001";
        ram_buffer(70917) := X"2413000C";
        ram_buffer(70918) := X"1000FF67";
        ram_buffer(70919) := X"241E0003";
        ram_buffer(70920) := X"3C100007";
        ram_buffer(70921) := X"3610FFFF";
        ram_buffer(70922) := X"2412FFFF";
        ram_buffer(70923) := X"0000B821";
        ram_buffer(70924) := X"3C04000F";
        ram_buffer(70925) := X"3484FFFF";
        ram_buffer(70926) := X"02042024";
        ram_buffer(70927) := X"02E02821";
        ram_buffer(70928) := X"1000FFA3";
        ram_buffer(70929) := X"240307FF";
        ram_buffer(70930) := X"0230102B";
        ram_buffer(70931) := X"1440002F";
        ram_buffer(70932) := X"00121042";
        ram_buffer(70933) := X"1211002A";
        ram_buffer(70934) := X"0243102B";
        ram_buffer(70935) := X"02403021";
        ram_buffer(70936) := X"26B5FFFF";
        ram_buffer(70937) := X"1000002D";
        ram_buffer(70938) := X"00009021";
        ram_buffer(70939) := X"02118825";
        ram_buffer(70940) := X"3C040008";
        ram_buffer(70941) := X"02248824";
        ram_buffer(70942) := X"162000BA";
        ram_buffer(70943) := X"00000000";
        ram_buffer(70944) := X"2484FFFF";
        ram_buffer(70945) := X"02048024";
        ram_buffer(70946) := X"02501025";
        ram_buffer(70947) := X"1440FFE8";
        ram_buffer(70948) := X"00000000";
        ram_buffer(70949) := X"3C040007";
        ram_buffer(70950) := X"00002821";
        ram_buffer(70951) := X"240307FF";
        ram_buffer(70952) := X"3484FFFF";
        ram_buffer(70953) := X"1000FF8A";
        ram_buffer(70954) := X"2412FFFF";
        ram_buffer(70955) := X"2442FFD8";
        ram_buffer(70956) := X"00478804";
        ram_buffer(70957) := X"1000FF7D";
        ram_buffer(70958) := X"00001821";
        ram_buffer(70959) := X"0C031D29";
        ram_buffer(70960) := X"AFA70010";
        ram_buffer(70961) := X"8FA70010";
        ram_buffer(70962) := X"1000FF6E";
        ram_buffer(70963) := X"24420020";
        ram_buffer(70964) := X"2442FFD8";
        ram_buffer(70965) := X"00458004";
        ram_buffer(70966) := X"1000FFB9";
        ram_buffer(70967) := X"00009021";
        ram_buffer(70968) := X"00A02021";
        ram_buffer(70969) := X"0C031D29";
        ram_buffer(70970) := X"AFA50010";
        ram_buffer(70971) := X"8FA70018";
        ram_buffer(70972) := X"8FA60014";
        ram_buffer(70973) := X"8FA50010";
        ram_buffer(70974) := X"1000FFA7";
        ram_buffer(70975) := X"24420020";
        ram_buffer(70976) := X"1440FFD7";
        ram_buffer(70977) := X"02403021";
        ram_buffer(70978) := X"00121042";
        ram_buffer(70979) := X"001037C0";
        ram_buffer(70980) := X"00C23025";
        ram_buffer(70981) := X"00108042";
        ram_buffer(70982) := X"001297C0";
        ram_buffer(70983) := X"00032602";
        ram_buffer(70984) := X"00118A00";
        ram_buffer(70985) := X"02248825";
        ram_buffer(70986) := X"00115402";
        ram_buffer(70987) := X"15400002";
        ram_buffer(70988) := X"020A001B";
        ram_buffer(70989) := X"0007000D";
        ram_buffer(70990) := X"322BFFFF";
        ram_buffer(70991) := X"00064C02";
        ram_buffer(70992) := X"00002012";
        ram_buffer(70993) := X"00006010";
        ram_buffer(70994) := X"000C6400";
        ram_buffer(70995) := X"012C4025";
        ram_buffer(70996) := X"01640018";
        ram_buffer(70997) := X"00008012";
        ram_buffer(70998) := X"0110102B";
        ram_buffer(70999) := X"1040000A";
        ram_buffer(71000) := X"00031A00";
        ram_buffer(71001) := X"01114021";
        ram_buffer(71002) := X"0111102B";
        ram_buffer(71003) := X"144000B0";
        ram_buffer(71004) := X"2485FFFF";
        ram_buffer(71005) := X"0110102B";
        ram_buffer(71006) := X"104000AD";
        ram_buffer(71007) := X"00000000";
        ram_buffer(71008) := X"2484FFFE";
        ram_buffer(71009) := X"01114021";
        ram_buffer(71010) := X"01104023";
        ram_buffer(71011) := X"15400002";
        ram_buffer(71012) := X"010A001B";
        ram_buffer(71013) := X"0007000D";
        ram_buffer(71014) := X"30C6FFFF";
        ram_buffer(71015) := X"00008012";
        ram_buffer(71016) := X"00004010";
        ram_buffer(71017) := X"00084400";
        ram_buffer(71018) := X"00C82825";
        ram_buffer(71019) := X"01700018";
        ram_buffer(71020) := X"00001012";
        ram_buffer(71021) := X"00A2302B";
        ram_buffer(71022) := X"10C0000A";
        ram_buffer(71023) := X"00000000";
        ram_buffer(71024) := X"00B12821";
        ram_buffer(71025) := X"00B1302B";
        ram_buffer(71026) := X"14C00097";
        ram_buffer(71027) := X"2608FFFF";
        ram_buffer(71028) := X"00A2302B";
        ram_buffer(71029) := X"10C00094";
        ram_buffer(71030) := X"00000000";
        ram_buffer(71031) := X"2610FFFE";
        ram_buffer(71032) := X"00B12821";
        ram_buffer(71033) := X"00042400";
        ram_buffer(71034) := X"00908025";
        ram_buffer(71035) := X"02030019";
        ram_buffer(71036) := X"00A22823";
        ram_buffer(71037) := X"00004010";
        ram_buffer(71038) := X"00A8102B";
        ram_buffer(71039) := X"00004812";
        ram_buffer(71040) := X"14400049";
        ram_buffer(71041) := X"01003021";
        ram_buffer(71042) := X"10A80045";
        ram_buffer(71043) := X"0249102B";
        ram_buffer(71044) := X"00A82823";
        ram_buffer(71045) := X"02494023";
        ram_buffer(71046) := X"0248902B";
        ram_buffer(71047) := X"00B22823";
        ram_buffer(71048) := X"122500AE";
        ram_buffer(71049) := X"00081402";
        ram_buffer(71050) := X"15400002";
        ram_buffer(71051) := X"00AA001B";
        ram_buffer(71052) := X"0007000D";
        ram_buffer(71053) := X"00002812";
        ram_buffer(71054) := X"00003010";
        ram_buffer(71055) := X"00063400";
        ram_buffer(71056) := X"00463025";
        ram_buffer(71057) := X"01650018";
        ram_buffer(71058) := X"00009012";
        ram_buffer(71059) := X"00D2102B";
        ram_buffer(71060) := X"1040000A";
        ram_buffer(71061) := X"00000000";
        ram_buffer(71062) := X"00D13021";
        ram_buffer(71063) := X"00D1102B";
        ram_buffer(71064) := X"144000A0";
        ram_buffer(71065) := X"24A4FFFF";
        ram_buffer(71066) := X"00D2102B";
        ram_buffer(71067) := X"1040009D";
        ram_buffer(71068) := X"00000000";
        ram_buffer(71069) := X"24A5FFFE";
        ram_buffer(71070) := X"00D13021";
        ram_buffer(71071) := X"00D23023";
        ram_buffer(71072) := X"15400002";
        ram_buffer(71073) := X"00CA001B";
        ram_buffer(71074) := X"0007000D";
        ram_buffer(71075) := X"3108FFFF";
        ram_buffer(71076) := X"00005012";
        ram_buffer(71077) := X"00003010";
        ram_buffer(71078) := X"00063400";
        ram_buffer(71079) := X"01062025";
        ram_buffer(71080) := X"016A0018";
        ram_buffer(71081) := X"00005812";
        ram_buffer(71082) := X"008B102B";
        ram_buffer(71083) := X"1040000A";
        ram_buffer(71084) := X"00000000";
        ram_buffer(71085) := X"00912021";
        ram_buffer(71086) := X"0091102B";
        ram_buffer(71087) := X"1440008B";
        ram_buffer(71088) := X"2546FFFF";
        ram_buffer(71089) := X"008B102B";
        ram_buffer(71090) := X"10400088";
        ram_buffer(71091) := X"00000000";
        ram_buffer(71092) := X"254AFFFE";
        ram_buffer(71093) := X"00912021";
        ram_buffer(71094) := X"00052C00";
        ram_buffer(71095) := X"00AA9025";
        ram_buffer(71096) := X"00720019";
        ram_buffer(71097) := X"008B2023";
        ram_buffer(71098) := X"00004010";
        ram_buffer(71099) := X"0088282B";
        ram_buffer(71100) := X"00004812";
        ram_buffer(71101) := X"00003012";
        ram_buffer(71102) := X"10A0003E";
        ram_buffer(71103) := X"01001021";
        ram_buffer(71104) := X"02242021";
        ram_buffer(71105) := X"0091502B";
        ram_buffer(71106) := X"1140007A";
        ram_buffer(71107) := X"2645FFFF";
        ram_buffer(71108) := X"1082004C";
        ram_buffer(71109) := X"00A09021";
        ram_buffer(71110) := X"10000017";
        ram_buffer(71111) := X"36520001";
        ram_buffer(71112) := X"1040004F";
        ram_buffer(71113) := X"00000000";
        ram_buffer(71114) := X"02439021";
        ram_buffer(71115) := X"0243202B";
        ram_buffer(71116) := X"00911021";
        ram_buffer(71117) := X"00452821";
        ram_buffer(71118) := X"0225102B";
        ram_buffer(71119) := X"10400033";
        ram_buffer(71120) := X"260CFFFF";
        ram_buffer(71121) := X"00A8102B";
        ram_buffer(71122) := X"1440007A";
        ram_buffer(71123) := X"00000000";
        ram_buffer(71124) := X"10C50040";
        ram_buffer(71125) := X"0249102B";
        ram_buffer(71126) := X"00A82823";
        ram_buffer(71127) := X"1000FFAD";
        ram_buffer(71128) := X"01808021";
        ram_buffer(71129) := X"2490FFFF";
        ram_buffer(71130) := X"2412FFFF";
        ram_buffer(71131) := X"1000FF30";
        ram_buffer(71132) := X"0000B821";
        ram_buffer(71133) := X"02E03821";
        ram_buffer(71134) := X"26A303FF";
        ram_buffer(71135) := X"1860003A";
        ram_buffer(71136) := X"00000000";
        ram_buffer(71137) := X"32420007";
        ram_buffer(71138) := X"10400009";
        ram_buffer(71139) := X"3C020100";
        ram_buffer(71140) := X"3242000F";
        ram_buffer(71141) := X"24040004";
        ram_buffer(71142) := X"10440004";
        ram_buffer(71143) := X"26420004";
        ram_buffer(71144) := X"0052902B";
        ram_buffer(71145) := X"02128021";
        ram_buffer(71146) := X"00409021";
        ram_buffer(71147) := X"3C020100";
        ram_buffer(71148) := X"02021024";
        ram_buffer(71149) := X"10400006";
        ram_buffer(71150) := X"286207FF";
        ram_buffer(71151) := X"3C02FEFF";
        ram_buffer(71152) := X"3442FFFF";
        ram_buffer(71153) := X"02028024";
        ram_buffer(71154) := X"26A30400";
        ram_buffer(71155) := X"286207FF";
        ram_buffer(71156) := X"1040FEBB";
        ram_buffer(71157) := X"00101740";
        ram_buffer(71158) := X"001290C2";
        ram_buffer(71159) := X"00108240";
        ram_buffer(71160) := X"00529025";
        ram_buffer(71161) := X"00102302";
        ram_buffer(71162) := X"306307FF";
        ram_buffer(71163) := X"1000FEB8";
        ram_buffer(71164) := X"30E50001";
        ram_buffer(71165) := X"1488FFC8";
        ram_buffer(71166) := X"00000000";
        ram_buffer(71167) := X"1120FFDE";
        ram_buffer(71168) := X"02242021";
        ram_buffer(71169) := X"1000FFC0";
        ram_buffer(71170) := X"0091502B";
        ram_buffer(71171) := X"1625FFD2";
        ram_buffer(71172) := X"00000000";
        ram_buffer(71173) := X"1080FFCC";
        ram_buffer(71174) := X"00A8102B";
        ram_buffer(71175) := X"02282823";
        ram_buffer(71176) := X"1000FF7C";
        ram_buffer(71177) := X"01808021";
        ram_buffer(71178) := X"1000FF6E";
        ram_buffer(71179) := X"01008021";
        ram_buffer(71180) := X"1000FF55";
        ram_buffer(71181) := X"00A02021";
        ram_buffer(71182) := X"15000045";
        ram_buffer(71183) := X"00034040";
        ram_buffer(71184) := X"00A09021";
        ram_buffer(71185) := X"1066FFCD";
        ram_buffer(71186) := X"26A303FF";
        ram_buffer(71187) := X"1000FFCB";
        ram_buffer(71188) := X"36520001";
        ram_buffer(71189) := X"14400037";
        ram_buffer(71190) := X"00000000";
        ram_buffer(71191) := X"01808021";
        ram_buffer(71192) := X"1000FF6C";
        ram_buffer(71193) := X"00002821";
        ram_buffer(71194) := X"1460002A";
        ram_buffer(71195) := X"24020001";
        ram_buffer(71196) := X"24030020";
        ram_buffer(71197) := X"00621823";
        ram_buffer(71198) := X"00702004";
        ram_buffer(71199) := X"00522806";
        ram_buffer(71200) := X"00721804";
        ram_buffer(71201) := X"0003182B";
        ram_buffer(71202) := X"00852825";
        ram_buffer(71203) := X"00A32825";
        ram_buffer(71204) := X"30A30007";
        ram_buffer(71205) := X"10600008";
        ram_buffer(71206) := X"00501006";
        ram_buffer(71207) := X"30A3000F";
        ram_buffer(71208) := X"24040004";
        ram_buffer(71209) := X"10640004";
        ram_buffer(71210) := X"00A01821";
        ram_buffer(71211) := X"24650004";
        ram_buffer(71212) := X"00A3182B";
        ram_buffer(71213) := X"00431021";
        ram_buffer(71214) := X"3C030080";
        ram_buffer(71215) := X"00431824";
        ram_buffer(71216) := X"1060002A";
        ram_buffer(71217) := X"00000000";
        ram_buffer(71218) := X"24030001";
        ram_buffer(71219) := X"00002021";
        ram_buffer(71220) := X"00009021";
        ram_buffer(71221) := X"1000FE7E";
        ram_buffer(71222) := X"30E50001";
        ram_buffer(71223) := X"1000FFA6";
        ram_buffer(71224) := X"2412FFFF";
        ram_buffer(71225) := X"1000FF65";
        ram_buffer(71226) := X"00802821";
        ram_buffer(71227) := X"1000FF7A";
        ram_buffer(71228) := X"00C05021";
        ram_buffer(71229) := X"0088502B";
        ram_buffer(71230) := X"15400014";
        ram_buffer(71231) := X"00000000";
        ram_buffer(71232) := X"1044FFCD";
        ram_buffer(71233) := X"0069402B";
        ram_buffer(71234) := X"00A09021";
        ram_buffer(71235) := X"1000FF9A";
        ram_buffer(71236) := X"36520001";
        ram_buffer(71237) := X"00431023";
        ram_buffer(71238) := X"28440039";
        ram_buffer(71239) := X"1480001C";
        ram_buffer(71240) := X"30E50001";
        ram_buffer(71241) := X"00001821";
        ram_buffer(71242) := X"00002021";
        ram_buffer(71243) := X"1000FE68";
        ram_buffer(71244) := X"00009021";
        ram_buffer(71245) := X"02439021";
        ram_buffer(71246) := X"0243302B";
        ram_buffer(71247) := X"00D13021";
        ram_buffer(71248) := X"00C52821";
        ram_buffer(71249) := X"1000FF32";
        ram_buffer(71250) := X"2610FFFE";
        ram_buffer(71251) := X"00034040";
        ram_buffer(71252) := X"0103182B";
        ram_buffer(71253) := X"00718821";
        ram_buffer(71254) := X"2645FFFE";
        ram_buffer(71255) := X"00912021";
        ram_buffer(71256) := X"1000FF6B";
        ram_buffer(71257) := X"01001821";
        ram_buffer(71258) := X"00602821";
        ram_buffer(71259) := X"00022240";
        ram_buffer(71260) := X"00042302";
        ram_buffer(71261) := X"00021740";
        ram_buffer(71262) := X"00A01821";
        ram_buffer(71263) := X"000318C2";
        ram_buffer(71264) := X"00629025";
        ram_buffer(71265) := X"30E50001";
        ram_buffer(71266) := X"1000FE51";
        ram_buffer(71267) := X"00001821";
        ram_buffer(71268) := X"28440020";
        ram_buffer(71269) := X"1480FFB6";
        ram_buffer(71270) := X"2404FFE1";
        ram_buffer(71271) := X"00831823";
        ram_buffer(71272) := X"24040020";
        ram_buffer(71273) := X"1044000F";
        ram_buffer(71274) := X"00701806";
        ram_buffer(71275) := X"00021023";
        ram_buffer(71276) := X"00501004";
        ram_buffer(71277) := X"00521025";
        ram_buffer(71278) := X"0002102B";
        ram_buffer(71279) := X"00621825";
        ram_buffer(71280) := X"30620007";
        ram_buffer(71281) := X"1040FFED";
        ram_buffer(71282) := X"00002021";
        ram_buffer(71283) := X"3062000F";
        ram_buffer(71284) := X"24040004";
        ram_buffer(71285) := X"1044FFE4";
        ram_buffer(71286) := X"00001021";
        ram_buffer(71287) := X"1000FFB4";
        ram_buffer(71288) := X"24650004";
        ram_buffer(71289) := X"1000FFF3";
        ram_buffer(71290) := X"00001021";
        ram_buffer(71291) := X"3484FFFF";
        ram_buffer(71292) := X"02048024";
        ram_buffer(71293) := X"1000FEA5";
        ram_buffer(71294) := X"02501025";
        ram_buffer(71295) := X"00041D02";
        ram_buffer(71296) := X"3C02000F";
        ram_buffer(71297) := X"3442FFFF";
        ram_buffer(71298) := X"00064502";
        ram_buffer(71299) := X"306307FF";
        ram_buffer(71300) := X"240A07FF";
        ram_buffer(71301) := X"00444824";
        ram_buffer(71302) := X"00A06021";
        ram_buffer(71303) := X"00461024";
        ram_buffer(71304) := X"000427C2";
        ram_buffer(71305) := X"00E05821";
        ram_buffer(71306) := X"310807FF";
        ram_buffer(71307) := X"106A0018";
        ram_buffer(71308) := X"000637C2";
        ram_buffer(71309) := X"240A07FF";
        ram_buffer(71310) := X"110A0010";
        ram_buffer(71311) := X"00000000";
        ram_buffer(71312) := X"10680003";
        ram_buffer(71313) := X"00000000";
        ram_buffer(71314) := X"03E00008";
        ram_buffer(71315) := X"24020001";
        ram_buffer(71316) := X"1522FFFD";
        ram_buffer(71317) := X"00000000";
        ram_buffer(71318) := X"158BFFFB";
        ram_buffer(71319) := X"00000000";
        ram_buffer(71320) := X"10860010";
        ram_buffer(71321) := X"00000000";
        ram_buffer(71322) := X"1460FFF7";
        ram_buffer(71323) := X"00000000";
        ram_buffer(71324) := X"01251025";
        ram_buffer(71325) := X"03E00008";
        ram_buffer(71326) := X"0002102B";
        ram_buffer(71327) := X"00473825";
        ram_buffer(71328) := X"10E0FFEF";
        ram_buffer(71329) := X"00000000";
        ram_buffer(71330) := X"03E00008";
        ram_buffer(71331) := X"24020001";
        ram_buffer(71332) := X"01255025";
        ram_buffer(71333) := X"1140FFE8";
        ram_buffer(71334) := X"240A07FF";
        ram_buffer(71335) := X"03E00008";
        ram_buffer(71336) := X"24020001";
        ram_buffer(71337) := X"03E00008";
        ram_buffer(71338) := X"00001021";
        ram_buffer(71339) := X"00041D02";
        ram_buffer(71340) := X"3C02000F";
        ram_buffer(71341) := X"3442FFFF";
        ram_buffer(71342) := X"00064502";
        ram_buffer(71343) := X"306307FF";
        ram_buffer(71344) := X"240907FF";
        ram_buffer(71345) := X"00445024";
        ram_buffer(71346) := X"310807FF";
        ram_buffer(71347) := X"00461024";
        ram_buffer(71348) := X"000427C2";
        ram_buffer(71349) := X"10690023";
        ram_buffer(71350) := X"000637C2";
        ram_buffer(71351) := X"240907FF";
        ram_buffer(71352) := X"11090016";
        ram_buffer(71353) := X"00474825";
        ram_buffer(71354) := X"1460000A";
        ram_buffer(71355) := X"01454825";
        ram_buffer(71356) := X"15000016";
        ram_buffer(71357) := X"2D2B0001";
        ram_buffer(71358) := X"00476025";
        ram_buffer(71359) := X"15800013";
        ram_buffer(71360) := X"00000000";
        ram_buffer(71361) := X"15200009";
        ram_buffer(71362) := X"00001021";
        ram_buffer(71363) := X"03E00008";
        ram_buffer(71364) := X"00000000";
        ram_buffer(71365) := X"15000003";
        ram_buffer(71366) := X"00474825";
        ram_buffer(71367) := X"11200003";
        ram_buffer(71368) := X"00000000";
        ram_buffer(71369) := X"10860014";
        ram_buffer(71370) := X"0103302A";
        ram_buffer(71371) := X"1080FFF7";
        ram_buffer(71372) := X"24020001";
        ram_buffer(71373) := X"03E00008";
        ram_buffer(71374) := X"2402FFFF";
        ram_buffer(71375) := X"1120FFEA";
        ram_buffer(71376) := X"00000000";
        ram_buffer(71377) := X"03E00008";
        ram_buffer(71378) := X"2402FFFE";
        ram_buffer(71379) := X"1160FFF5";
        ram_buffer(71380) := X"00000000";
        ram_buffer(71381) := X"10C0FFF7";
        ram_buffer(71382) := X"00000000";
        ram_buffer(71383) := X"03E00008";
        ram_buffer(71384) := X"24020001";
        ram_buffer(71385) := X"01454825";
        ram_buffer(71386) := X"1120FFDD";
        ram_buffer(71387) := X"240907FF";
        ram_buffer(71388) := X"1000FFF4";
        ram_buffer(71389) := X"00000000";
        ram_buffer(71390) := X"14C0FFEC";
        ram_buffer(71391) := X"00000000";
        ram_buffer(71392) := X"0068182A";
        ram_buffer(71393) := X"14600007";
        ram_buffer(71394) := X"004A182B";
        ram_buffer(71395) := X"1460FFE7";
        ram_buffer(71396) := X"00000000";
        ram_buffer(71397) := X"11420009";
        ram_buffer(71398) := X"0142102B";
        ram_buffer(71399) := X"10400005";
        ram_buffer(71400) := X"00000000";
        ram_buffer(71401) := X"1480FFED";
        ram_buffer(71402) := X"00000000";
        ram_buffer(71403) := X"1000FFE1";
        ram_buffer(71404) := X"00000000";
        ram_buffer(71405) := X"03E00008";
        ram_buffer(71406) := X"00000000";
        ram_buffer(71407) := X"00E5102B";
        ram_buffer(71408) := X"1440FFDA";
        ram_buffer(71409) := X"00000000";
        ram_buffer(71410) := X"00A7282B";
        ram_buffer(71411) := X"14A0FFF5";
        ram_buffer(71412) := X"00000000";
        ram_buffer(71413) := X"03E00008";
        ram_buffer(71414) := X"00001021";
        ram_buffer(71415) := X"00041D02";
        ram_buffer(71416) := X"3C02000F";
        ram_buffer(71417) := X"3442FFFF";
        ram_buffer(71418) := X"00064502";
        ram_buffer(71419) := X"306307FF";
        ram_buffer(71420) := X"240907FF";
        ram_buffer(71421) := X"00445024";
        ram_buffer(71422) := X"310807FF";
        ram_buffer(71423) := X"00461024";
        ram_buffer(71424) := X"000427C2";
        ram_buffer(71425) := X"10690021";
        ram_buffer(71426) := X"000637C2";
        ram_buffer(71427) := X"240907FF";
        ram_buffer(71428) := X"11090014";
        ram_buffer(71429) := X"00474825";
        ram_buffer(71430) := X"1460000A";
        ram_buffer(71431) := X"01454825";
        ram_buffer(71432) := X"15000014";
        ram_buffer(71433) := X"2D2B0001";
        ram_buffer(71434) := X"00476025";
        ram_buffer(71435) := X"15800011";
        ram_buffer(71436) := X"00000000";
        ram_buffer(71437) := X"15200007";
        ram_buffer(71438) := X"00001021";
        ram_buffer(71439) := X"03E00008";
        ram_buffer(71440) := X"00000000";
        ram_buffer(71441) := X"11000016";
        ram_buffer(71442) := X"00474825";
        ram_buffer(71443) := X"10C40018";
        ram_buffer(71444) := X"0103482A";
        ram_buffer(71445) := X"1080FFF9";
        ram_buffer(71446) := X"24020001";
        ram_buffer(71447) := X"03E00008";
        ram_buffer(71448) := X"2402FFFF";
        ram_buffer(71449) := X"1120FFEC";
        ram_buffer(71450) := X"00000000";
        ram_buffer(71451) := X"03E00008";
        ram_buffer(71452) := X"24020002";
        ram_buffer(71453) := X"1160FFF5";
        ram_buffer(71454) := X"00000000";
        ram_buffer(71455) := X"10C0FFF7";
        ram_buffer(71456) := X"00000000";
        ram_buffer(71457) := X"03E00008";
        ram_buffer(71458) := X"24020001";
        ram_buffer(71459) := X"01454825";
        ram_buffer(71460) := X"1120FFDF";
        ram_buffer(71461) := X"240907FF";
        ram_buffer(71462) := X"03E00008";
        ram_buffer(71463) := X"24020002";
        ram_buffer(71464) := X"1520FFEA";
        ram_buffer(71465) := X"00000000";
        ram_buffer(71466) := X"1000FFEA";
        ram_buffer(71467) := X"00000000";
        ram_buffer(71468) := X"11200005";
        ram_buffer(71469) := X"00000000";
        ram_buffer(71470) := X"14C0FFE8";
        ram_buffer(71471) := X"24020001";
        ram_buffer(71472) := X"03E00008";
        ram_buffer(71473) := X"00000000";
        ram_buffer(71474) := X"0068182A";
        ram_buffer(71475) := X"1460FFEB";
        ram_buffer(71476) := X"00000000";
        ram_buffer(71477) := X"004A182B";
        ram_buffer(71478) := X"1460FFDE";
        ram_buffer(71479) := X"00000000";
        ram_buffer(71480) := X"11420009";
        ram_buffer(71481) := X"0142102B";
        ram_buffer(71482) := X"10400005";
        ram_buffer(71483) := X"00000000";
        ram_buffer(71484) := X"1480FFE4";
        ram_buffer(71485) := X"00000000";
        ram_buffer(71486) := X"1000FFD8";
        ram_buffer(71487) := X"00000000";
        ram_buffer(71488) := X"03E00008";
        ram_buffer(71489) := X"00000000";
        ram_buffer(71490) := X"00E5102B";
        ram_buffer(71491) := X"1440FFD1";
        ram_buffer(71492) := X"00000000";
        ram_buffer(71493) := X"00A7282B";
        ram_buffer(71494) := X"14A0FFF5";
        ram_buffer(71495) := X"00000000";
        ram_buffer(71496) := X"03E00008";
        ram_buffer(71497) := X"00001021";
        ram_buffer(71498) := X"27BDFFB8";
        ram_buffer(71499) := X"00044502";
        ram_buffer(71500) := X"AFB00020";
        ram_buffer(71501) := X"3C10000F";
        ram_buffer(71502) := X"AFB60038";
        ram_buffer(71503) := X"AFB3002C";
        ram_buffer(71504) := X"3610FFFF";
        ram_buffer(71505) := X"00049FC2";
        ram_buffer(71506) := X"311607FF";
        ram_buffer(71507) := X"AFB50034";
        ram_buffer(71508) := X"AFB40030";
        ram_buffer(71509) := X"AFBF0044";
        ram_buffer(71510) := X"AFBE0040";
        ram_buffer(71511) := X"AFB7003C";
        ram_buffer(71512) := X"AFB20028";
        ram_buffer(71513) := X"AFB10024";
        ram_buffer(71514) := X"0204A824";
        ram_buffer(71515) := X"12C00075";
        ram_buffer(71516) := X"0260A021";
        ram_buffer(71517) := X"240207FF";
        ram_buffer(71518) := X"12C2002A";
        ram_buffer(71519) := X"00A08821";
        ram_buffer(71520) := X"3C100010";
        ram_buffer(71521) := X"02B08025";
        ram_buffer(71522) := X"001080C0";
        ram_buffer(71523) := X"00052742";
        ram_buffer(71524) := X"0090A825";
        ram_buffer(71525) := X"000588C0";
        ram_buffer(71526) := X"26D6FC01";
        ram_buffer(71527) := X"00009021";
        ram_buffer(71528) := X"0000B821";
        ram_buffer(71529) := X"00064D02";
        ram_buffer(71530) := X"3C02000F";
        ram_buffer(71531) := X"3442FFFF";
        ram_buffer(71532) := X"312807FF";
        ram_buffer(71533) := X"00E02021";
        ram_buffer(71534) := X"00468024";
        ram_buffer(71535) := X"11000028";
        ram_buffer(71536) := X"0006F7C2";
        ram_buffer(71537) := X"240207FF";
        ram_buffer(71538) := X"1102007A";
        ram_buffer(71539) := X"3C020010";
        ram_buffer(71540) := X"02028025";
        ram_buffer(71541) := X"001080C0";
        ram_buffer(71542) := X"00071742";
        ram_buffer(71543) := X"00508025";
        ram_buffer(71544) := X"000720C0";
        ram_buffer(71545) := X"2508FC01";
        ram_buffer(71546) := X"00001021";
        ram_buffer(71547) := X"00523825";
        ram_buffer(71548) := X"02C84021";
        ram_buffer(71549) := X"2CE50010";
        ram_buffer(71550) := X"027E1826";
        ram_buffer(71551) := X"10A00096";
        ram_buffer(71552) := X"250A0001";
        ram_buffer(71553) := X"3C09100D";
        ram_buffer(71554) := X"00073880";
        ram_buffer(71555) := X"2529B620";
        ram_buffer(71556) := X"01273821";
        ram_buffer(71557) := X"8CE50000";
        ram_buffer(71558) := X"00000000";
        ram_buffer(71559) := X"00A00008";
        ram_buffer(71560) := X"00000000";
        ram_buffer(71561) := X"02A52825";
        ram_buffer(71562) := X"14A00076";
        ram_buffer(71563) := X"2412000C";
        ram_buffer(71564) := X"00064D02";
        ram_buffer(71565) := X"3C02000F";
        ram_buffer(71566) := X"3442FFFF";
        ram_buffer(71567) := X"312807FF";
        ram_buffer(71568) := X"24120008";
        ram_buffer(71569) := X"0000A821";
        ram_buffer(71570) := X"00008821";
        ram_buffer(71571) := X"24170002";
        ram_buffer(71572) := X"00E02021";
        ram_buffer(71573) := X"00468024";
        ram_buffer(71574) := X"1500FFDA";
        ram_buffer(71575) := X"0006F7C2";
        ram_buffer(71576) := X"02071025";
        ram_buffer(71577) := X"1040005E";
        ram_buffer(71578) := X"00002021";
        ram_buffer(71579) := X"120000DF";
        ram_buffer(71580) := X"00E02021";
        ram_buffer(71581) := X"02002021";
        ram_buffer(71582) := X"0C031D29";
        ram_buffer(71583) := X"AFA70010";
        ram_buffer(71584) := X"8FA70010";
        ram_buffer(71585) := X"2448FFF5";
        ram_buffer(71586) := X"2903001D";
        ram_buffer(71587) := X"106000D3";
        ram_buffer(71588) := X"2403001D";
        ram_buffer(71589) := X"2444FFF8";
        ram_buffer(71590) := X"00681823";
        ram_buffer(71591) := X"00908004";
        ram_buffer(71592) := X"00671806";
        ram_buffer(71593) := X"00708025";
        ram_buffer(71594) := X"00872004";
        ram_buffer(71595) := X"2407FC02";
        ram_buffer(71596) := X"00E84023";
        ram_buffer(71597) := X"1000FFCD";
        ram_buffer(71598) := X"00001021";
        ram_buffer(71599) := X"03C01821";
        ram_buffer(71600) := X"24050002";
        ram_buffer(71601) := X"10450042";
        ram_buffer(71602) := X"24050003";
        ram_buffer(71603) := X"10450119";
        ram_buffer(71604) := X"3C050007";
        ram_buffer(71605) := X"24050001";
        ram_buffer(71606) := X"14450092";
        ram_buffer(71607) := X"01404021";
        ram_buffer(71608) := X"00008021";
        ram_buffer(71609) := X"00002021";
        ram_buffer(71610) := X"00008821";
        ram_buffer(71611) := X"00101500";
        ram_buffer(71612) := X"3C10000F";
        ram_buffer(71613) := X"3610FFFF";
        ram_buffer(71614) := X"00908024";
        ram_buffer(71615) := X"02028025";
        ram_buffer(71616) := X"00031FC0";
        ram_buffer(71617) := X"02031825";
        ram_buffer(71618) := X"8FBF0044";
        ram_buffer(71619) := X"00602021";
        ram_buffer(71620) := X"8FBE0040";
        ram_buffer(71621) := X"02201821";
        ram_buffer(71622) := X"8FB7003C";
        ram_buffer(71623) := X"8FB60038";
        ram_buffer(71624) := X"8FB50034";
        ram_buffer(71625) := X"8FB40030";
        ram_buffer(71626) := X"8FB3002C";
        ram_buffer(71627) := X"8FB20028";
        ram_buffer(71628) := X"8FB10024";
        ram_buffer(71629) := X"8FB00020";
        ram_buffer(71630) := X"00801021";
        ram_buffer(71631) := X"03E00008";
        ram_buffer(71632) := X"27BD0048";
        ram_buffer(71633) := X"02A51025";
        ram_buffer(71634) := X"1040002A";
        ram_buffer(71635) := X"24120004";
        ram_buffer(71636) := X"AFA70018";
        ram_buffer(71637) := X"12A000AD";
        ram_buffer(71638) := X"AFA60014";
        ram_buffer(71639) := X"02A02021";
        ram_buffer(71640) := X"0C031D29";
        ram_buffer(71641) := X"AFA50010";
        ram_buffer(71642) := X"8FA50010";
        ram_buffer(71643) := X"8FA60014";
        ram_buffer(71644) := X"8FA70018";
        ram_buffer(71645) := X"2443FFF5";
        ram_buffer(71646) := X"2864001D";
        ram_buffer(71647) := X"108000A0";
        ram_buffer(71648) := X"2444FFD8";
        ram_buffer(71649) := X"2408001D";
        ram_buffer(71650) := X"2451FFF8";
        ram_buffer(71651) := X"01034023";
        ram_buffer(71652) := X"02352004";
        ram_buffer(71653) := X"01054006";
        ram_buffer(71654) := X"0104A825";
        ram_buffer(71655) := X"02258804";
        ram_buffer(71656) := X"2408FC02";
        ram_buffer(71657) := X"0103B023";
        ram_buffer(71658) := X"00009021";
        ram_buffer(71659) := X"1000FF7D";
        ram_buffer(71660) := X"0000B821";
        ram_buffer(71661) := X"02073825";
        ram_buffer(71662) := X"14E0000C";
        ram_buffer(71663) := X"00000000";
        ram_buffer(71664) := X"00008021";
        ram_buffer(71665) := X"00002021";
        ram_buffer(71666) := X"1000FF88";
        ram_buffer(71667) := X"24020002";
        ram_buffer(71668) := X"241007FF";
        ram_buffer(71669) := X"00002021";
        ram_buffer(71670) := X"1000FFC4";
        ram_buffer(71671) := X"00008821";
        ram_buffer(71672) := X"00008021";
        ram_buffer(71673) := X"1000FF81";
        ram_buffer(71674) := X"24020001";
        ram_buffer(71675) := X"1000FF7F";
        ram_buffer(71676) := X"24020003";
        ram_buffer(71677) := X"0000A821";
        ram_buffer(71678) := X"00008821";
        ram_buffer(71679) := X"1000FF69";
        ram_buffer(71680) := X"24170001";
        ram_buffer(71681) := X"1000FF67";
        ram_buffer(71682) := X"24170003";
        ram_buffer(71683) := X"3C100007";
        ram_buffer(71684) := X"3605FFFF";
        ram_buffer(71685) := X"2411FFFF";
        ram_buffer(71686) := X"0000A021";
        ram_buffer(71687) := X"3C10000F";
        ram_buffer(71688) := X"3610FFFF";
        ram_buffer(71689) := X"00B02024";
        ram_buffer(71690) := X"32830001";
        ram_buffer(71691) := X"1000FFAF";
        ram_buffer(71692) := X"241007FF";
        ram_buffer(71693) := X"02A08021";
        ram_buffer(71694) := X"02202021";
        ram_buffer(71695) := X"1000FFA0";
        ram_buffer(71696) := X"02E01021";
        ram_buffer(71697) := X"02A08021";
        ram_buffer(71698) := X"02202021";
        ram_buffer(71699) := X"02601821";
        ram_buffer(71700) := X"1000FF9B";
        ram_buffer(71701) := X"02E01021";
        ram_buffer(71702) := X"02300019";
        ram_buffer(71703) := X"00003812";
        ram_buffer(71704) := X"00003010";
        ram_buffer(71705) := X"00000000";
        ram_buffer(71706) := X"00000000";
        ram_buffer(71707) := X"02240019";
        ram_buffer(71708) := X"00006812";
        ram_buffer(71709) := X"00006010";
        ram_buffer(71710) := X"01874821";
        ram_buffer(71711) := X"0127102B";
        ram_buffer(71712) := X"02150019";
        ram_buffer(71713) := X"00008010";
        ram_buffer(71714) := X"00008812";
        ram_buffer(71715) := X"00D13821";
        ram_buffer(71716) := X"00000000";
        ram_buffer(71717) := X"00950019";
        ram_buffer(71718) := X"0047A821";
        ram_buffer(71719) := X"00E6382B";
        ram_buffer(71720) := X"02A2302B";
        ram_buffer(71721) := X"00E63025";
        ram_buffer(71722) := X"00D03021";
        ram_buffer(71723) := X"3C020100";
        ram_buffer(71724) := X"00002812";
        ram_buffer(71725) := X"01253821";
        ram_buffer(71726) := X"00E5282B";
        ram_buffer(71727) := X"00002010";
        ram_buffer(71728) := X"02A48021";
        ram_buffer(71729) := X"00B04821";
        ram_buffer(71730) := X"0204202B";
        ram_buffer(71731) := X"0125802B";
        ram_buffer(71732) := X"00908025";
        ram_buffer(71733) := X"00D08021";
        ram_buffer(71734) := X"00072240";
        ram_buffer(71735) := X"00102A40";
        ram_buffer(71736) := X"008D2025";
        ram_buffer(71737) := X"000985C2";
        ram_buffer(71738) := X"0004202B";
        ram_buffer(71739) := X"00B08025";
        ram_buffer(71740) := X"00073DC2";
        ram_buffer(71741) := X"00873825";
        ram_buffer(71742) := X"02021024";
        ram_buffer(71743) := X"00092240";
        ram_buffer(71744) := X"10400008";
        ram_buffer(71745) := X"00E42025";
        ram_buffer(71746) := X"00041042";
        ram_buffer(71747) := X"30840001";
        ram_buffer(71748) := X"00102FC0";
        ram_buffer(71749) := X"00442025";
        ram_buffer(71750) := X"00A42025";
        ram_buffer(71751) := X"00108042";
        ram_buffer(71752) := X"01404021";
        ram_buffer(71753) := X"250203FF";
        ram_buffer(71754) := X"18400043";
        ram_buffer(71755) := X"00000000";
        ram_buffer(71756) := X"30850007";
        ram_buffer(71757) := X"10A00009";
        ram_buffer(71758) := X"3C050100";
        ram_buffer(71759) := X"3085000F";
        ram_buffer(71760) := X"24060004";
        ram_buffer(71761) := X"10A60004";
        ram_buffer(71762) := X"24850004";
        ram_buffer(71763) := X"00A4202B";
        ram_buffer(71764) := X"02048021";
        ram_buffer(71765) := X"00A02021";
        ram_buffer(71766) := X"3C050100";
        ram_buffer(71767) := X"02052824";
        ram_buffer(71768) := X"10A00006";
        ram_buffer(71769) := X"284507FF";
        ram_buffer(71770) := X"3C02FEFF";
        ram_buffer(71771) := X"3442FFFF";
        ram_buffer(71772) := X"02028024";
        ram_buffer(71773) := X"25020400";
        ram_buffer(71774) := X"284507FF";
        ram_buffer(71775) := X"10A0FF94";
        ram_buffer(71776) := X"00000000";
        ram_buffer(71777) := X"000420C2";
        ram_buffer(71778) := X"00108F40";
        ram_buffer(71779) := X"00108240";
        ram_buffer(71780) := X"02248825";
        ram_buffer(71781) := X"00102302";
        ram_buffer(71782) := X"1000FF54";
        ram_buffer(71783) := X"305007FF";
        ram_buffer(71784) := X"3C050008";
        ram_buffer(71785) := X"02B08025";
        ram_buffer(71786) := X"02058024";
        ram_buffer(71787) := X"1600001F";
        ram_buffer(71788) := X"24A5FFFF";
        ram_buffer(71789) := X"02A52824";
        ram_buffer(71790) := X"02251025";
        ram_buffer(71791) := X"1440FF97";
        ram_buffer(71792) := X"00000000";
        ram_buffer(71793) := X"3C040007";
        ram_buffer(71794) := X"00001821";
        ram_buffer(71795) := X"241007FF";
        ram_buffer(71796) := X"3484FFFF";
        ram_buffer(71797) := X"1000FF45";
        ram_buffer(71798) := X"2411FFFF";
        ram_buffer(71799) := X"2442FFD8";
        ram_buffer(71800) := X"00478004";
        ram_buffer(71801) := X"1000FF31";
        ram_buffer(71802) := X"00002021";
        ram_buffer(71803) := X"0C031D29";
        ram_buffer(71804) := X"AFA70010";
        ram_buffer(71805) := X"8FA70010";
        ram_buffer(71806) := X"1000FF22";
        ram_buffer(71807) := X"24420020";
        ram_buffer(71808) := X"0085A804";
        ram_buffer(71809) := X"1000FF66";
        ram_buffer(71810) := X"00008821";
        ram_buffer(71811) := X"00A02021";
        ram_buffer(71812) := X"0C031D29";
        ram_buffer(71813) := X"AFA50010";
        ram_buffer(71814) := X"8FA70018";
        ram_buffer(71815) := X"8FA60014";
        ram_buffer(71816) := X"8FA50010";
        ram_buffer(71817) := X"1000FF53";
        ram_buffer(71818) := X"24420020";
        ram_buffer(71819) := X"2411FFFF";
        ram_buffer(71820) := X"1000FF7A";
        ram_buffer(71821) := X"0000A021";
        ram_buffer(71822) := X"1440001B";
        ram_buffer(71823) := X"24050001";
        ram_buffer(71824) := X"24020020";
        ram_buffer(71825) := X"00451023";
        ram_buffer(71826) := X"00503004";
        ram_buffer(71827) := X"00A43806";
        ram_buffer(71828) := X"00441004";
        ram_buffer(71829) := X"0002102B";
        ram_buffer(71830) := X"00C73025";
        ram_buffer(71831) := X"00C23025";
        ram_buffer(71832) := X"30C20007";
        ram_buffer(71833) := X"10400008";
        ram_buffer(71834) := X"00B02806";
        ram_buffer(71835) := X"30C2000F";
        ram_buffer(71836) := X"24040004";
        ram_buffer(71837) := X"10440004";
        ram_buffer(71838) := X"00C01021";
        ram_buffer(71839) := X"24460004";
        ram_buffer(71840) := X"00C2102B";
        ram_buffer(71841) := X"00A22821";
        ram_buffer(71842) := X"3C020080";
        ram_buffer(71843) := X"00A21024";
        ram_buffer(71844) := X"1040001D";
        ram_buffer(71845) := X"00000000";
        ram_buffer(71846) := X"24100001";
        ram_buffer(71847) := X"00002021";
        ram_buffer(71848) := X"1000FF12";
        ram_buffer(71849) := X"00008821";
        ram_buffer(71850) := X"00A22823";
        ram_buffer(71851) := X"28A60039";
        ram_buffer(71852) := X"10C0FF0B";
        ram_buffer(71853) := X"28A60020";
        ram_buffer(71854) := X"14C0FFE1";
        ram_buffer(71855) := X"2406FFE1";
        ram_buffer(71856) := X"00C21023";
        ram_buffer(71857) := X"00503006";
        ram_buffer(71858) := X"24020020";
        ram_buffer(71859) := X"10A20003";
        ram_buffer(71860) := X"00001021";
        ram_buffer(71861) := X"00051023";
        ram_buffer(71862) := X"00501004";
        ram_buffer(71863) := X"00441025";
        ram_buffer(71864) := X"0002102B";
        ram_buffer(71865) := X"00C21025";
        ram_buffer(71866) := X"30450007";
        ram_buffer(71867) := X"14A0000B";
        ram_buffer(71868) := X"00002021";
        ram_buffer(71869) := X"000210C2";
        ram_buffer(71870) := X"00A28825";
        ram_buffer(71871) := X"1000FEFB";
        ram_buffer(71872) := X"00008021";
        ram_buffer(71873) := X"00002821";
        ram_buffer(71874) := X"00052240";
        ram_buffer(71875) := X"00042302";
        ram_buffer(71876) := X"00052F40";
        ram_buffer(71877) := X"1000FFF7";
        ram_buffer(71878) := X"00C01021";
        ram_buffer(71879) := X"3044000F";
        ram_buffer(71880) := X"24050004";
        ram_buffer(71881) := X"1085FFF7";
        ram_buffer(71882) := X"00403021";
        ram_buffer(71883) := X"1000FFD3";
        ram_buffer(71884) := X"00002821";
        ram_buffer(71885) := X"34A5FFFF";
        ram_buffer(71886) := X"02052824";
        ram_buffer(71887) := X"00851025";
        ram_buffer(71888) := X"00808821";
        ram_buffer(71889) := X"1000FF9D";
        ram_buffer(71890) := X"0060A021";
        ram_buffer(71891) := X"3C08000F";
        ram_buffer(71892) := X"3508FFFF";
        ram_buffer(71893) := X"01044824";
        ram_buffer(71894) := X"00065502";
        ram_buffer(71895) := X"01064024";
        ram_buffer(71896) := X"27BDFFD8";
        ram_buffer(71897) := X"00041502";
        ram_buffer(71898) := X"00056742";
        ram_buffer(71899) := X"00075F42";
        ram_buffer(71900) := X"000948C0";
        ram_buffer(71901) := X"000840C0";
        ram_buffer(71902) := X"314A07FF";
        ram_buffer(71903) := X"240307FF";
        ram_buffer(71904) := X"000528C0";
        ram_buffer(71905) := X"AFB10018";
        ram_buffer(71906) := X"AFB00014";
        ram_buffer(71907) := X"305107FF";
        ram_buffer(71908) := X"AFBF0024";
        ram_buffer(71909) := X"AFB30020";
        ram_buffer(71910) := X"AFB2001C";
        ram_buffer(71911) := X"000487C2";
        ram_buffer(71912) := X"012C1025";
        ram_buffer(71913) := X"000637C2";
        ram_buffer(71914) := X"010B4025";
        ram_buffer(71915) := X"11430012";
        ram_buffer(71916) := X"000738C0";
        ram_buffer(71917) := X"38C60001";
        ram_buffer(71918) := X"10D00066";
        ram_buffer(71919) := X"022A2023";
        ram_buffer(71920) := X"188000D5";
        ram_buffer(71921) := X"00000000";
        ram_buffer(71922) := X"15400010";
        ram_buffer(71923) := X"240307FF";
        ram_buffer(71924) := X"01071825";
        ram_buffer(71925) := X"10600085";
        ram_buffer(71926) := X"240307FF";
        ram_buffer(71927) := X"2484FFFF";
        ram_buffer(71928) := X"148000AF";
        ram_buffer(71929) := X"00A79023";
        ram_buffer(71930) := X"00481023";
        ram_buffer(71931) := X"00B2282B";
        ram_buffer(71932) := X"1000001A";
        ram_buffer(71933) := X"00451023";
        ram_buffer(71934) := X"01071825";
        ram_buffer(71935) := X"1460FFEE";
        ram_buffer(71936) := X"00000000";
        ram_buffer(71937) := X"1000FFEC";
        ram_buffer(71938) := X"38C60001";
        ram_buffer(71939) := X"122300A6";
        ram_buffer(71940) := X"3C030080";
        ram_buffer(71941) := X"01034025";
        ram_buffer(71942) := X"28830039";
        ram_buffer(71943) := X"106000E8";
        ram_buffer(71944) := X"28830020";
        ram_buffer(71945) := X"1060010C";
        ram_buffer(71946) := X"24060020";
        ram_buffer(71947) := X"00C43023";
        ram_buffer(71948) := X"00C81804";
        ram_buffer(71949) := X"00879006";
        ram_buffer(71950) := X"00C73804";
        ram_buffer(71951) := X"00721825";
        ram_buffer(71952) := X"0007382B";
        ram_buffer(71953) := X"00673825";
        ram_buffer(71954) := X"00884006";
        ram_buffer(71955) := X"00A79023";
        ram_buffer(71956) := X"00484023";
        ram_buffer(71957) := X"00B2282B";
        ram_buffer(71958) := X"01051023";
        ram_buffer(71959) := X"3C130080";
        ram_buffer(71960) := X"00531824";
        ram_buffer(71961) := X"106000A8";
        ram_buffer(71962) := X"32430007";
        ram_buffer(71963) := X"2673FFFF";
        ram_buffer(71964) := X"00539824";
        ram_buffer(71965) := X"126000BB";
        ram_buffer(71966) := X"00000000";
        ram_buffer(71967) := X"0C031D29";
        ram_buffer(71968) := X"02602021";
        ram_buffer(71969) := X"2446FFF8";
        ram_buffer(71970) := X"28C30020";
        ram_buffer(71971) := X"106000BD";
        ram_buffer(71972) := X"2442FFD8";
        ram_buffer(71973) := X"00061823";
        ram_buffer(71974) := X"00721806";
        ram_buffer(71975) := X"00D31004";
        ram_buffer(71976) := X"00629825";
        ram_buffer(71977) := X"00D1102A";
        ram_buffer(71978) := X"144000BA";
        ram_buffer(71979) := X"00D29004";
        ram_buffer(71980) := X"00D13023";
        ram_buffer(71981) := X"24C20001";
        ram_buffer(71982) := X"28430020";
        ram_buffer(71983) := X"106000DB";
        ram_buffer(71984) := X"24030020";
        ram_buffer(71985) := X"00621823";
        ram_buffer(71986) := X"00522006";
        ram_buffer(71987) := X"00723804";
        ram_buffer(71988) := X"00731804";
        ram_buffer(71989) := X"00641825";
        ram_buffer(71990) := X"0007382B";
        ram_buffer(71991) := X"00679025";
        ram_buffer(71992) := X"00531006";
        ram_buffer(71993) := X"32430007";
        ram_buffer(71994) := X"00008821";
        ram_buffer(71995) := X"10600043";
        ram_buffer(71996) := X"3C030080";
        ram_buffer(71997) := X"3243000F";
        ram_buffer(71998) := X"24040004";
        ram_buffer(71999) := X"1064003E";
        ram_buffer(72000) := X"26430004";
        ram_buffer(72001) := X"0072382B";
        ram_buffer(72002) := X"00471021";
        ram_buffer(72003) := X"00609021";
        ram_buffer(72004) := X"3C030080";
        ram_buffer(72005) := X"00431824";
        ram_buffer(72006) := X"1460003B";
        ram_buffer(72007) := X"00000000";
        ram_buffer(72008) := X"00021F40";
        ram_buffer(72009) := X"001238C2";
        ram_buffer(72010) := X"00E33825";
        ram_buffer(72011) := X"000218C2";
        ram_buffer(72012) := X"240207FF";
        ram_buffer(72013) := X"12220062";
        ram_buffer(72014) := X"00000000";
        ram_buffer(72015) := X"3C06000F";
        ram_buffer(72016) := X"34C6FFFF";
        ram_buffer(72017) := X"00662824";
        ram_buffer(72018) := X"322207FF";
        ram_buffer(72019) := X"1000003C";
        ram_buffer(72020) := X"32030001";
        ram_buffer(72021) := X"022A1823";
        ram_buffer(72022) := X"186000A1";
        ram_buffer(72023) := X"00000000";
        ram_buffer(72024) := X"11400048";
        ram_buffer(72025) := X"01072025";
        ram_buffer(72026) := X"240407FF";
        ram_buffer(72027) := X"122400E9";
        ram_buffer(72028) := X"3C040080";
        ram_buffer(72029) := X"01044025";
        ram_buffer(72030) := X"28640039";
        ram_buffer(72031) := X"148000EB";
        ram_buffer(72032) := X"28640020";
        ram_buffer(72033) := X"01073825";
        ram_buffer(72034) := X"0007382B";
        ram_buffer(72035) := X"00004021";
        ram_buffer(72036) := X"00E59021";
        ram_buffer(72037) := X"01024021";
        ram_buffer(72038) := X"0245282B";
        ram_buffer(72039) := X"00A81021";
        ram_buffer(72040) := X"3C030080";
        ram_buffer(72041) := X"00431824";
        ram_buffer(72042) := X"10600103";
        ram_buffer(72043) := X"240307FF";
        ram_buffer(72044) := X"26310001";
        ram_buffer(72045) := X"1223010B";
        ram_buffer(72046) := X"00000000";
        ram_buffer(72047) := X"3C03FF7F";
        ram_buffer(72048) := X"3463FFFF";
        ram_buffer(72049) := X"00431024";
        ram_buffer(72050) := X"32470001";
        ram_buffer(72051) := X"00121842";
        ram_buffer(72052) := X"00673825";
        ram_buffer(72053) := X"000297C0";
        ram_buffer(72054) := X"02479025";
        ram_buffer(72055) := X"00021042";
        ram_buffer(72056) := X"32430007";
        ram_buffer(72057) := X"1000FFC1";
        ram_buffer(72058) := X"00C08021";
        ram_buffer(72059) := X"1223002F";
        ram_buffer(72060) := X"00451825";
        ram_buffer(72061) := X"00A09021";
        ram_buffer(72062) := X"3C030080";
        ram_buffer(72063) := X"00431824";
        ram_buffer(72064) := X"1060FFC8";
        ram_buffer(72065) := X"00021F40";
        ram_buffer(72066) := X"26260001";
        ram_buffer(72067) := X"240307FF";
        ram_buffer(72068) := X"10C30067";
        ram_buffer(72069) := X"32030001";
        ram_buffer(72070) := X"3C05FF7F";
        ram_buffer(72071) := X"34A5FFFF";
        ram_buffer(72072) := X"00451024";
        ram_buffer(72073) := X"00021F40";
        ram_buffer(72074) := X"001238C2";
        ram_buffer(72075) := X"00021240";
        ram_buffer(72076) := X"00673825";
        ram_buffer(72077) := X"00022B02";
        ram_buffer(72078) := X"32030001";
        ram_buffer(72079) := X"30C207FF";
        ram_buffer(72080) := X"00023500";
        ram_buffer(72081) := X"3C02000F";
        ram_buffer(72082) := X"3442FFFF";
        ram_buffer(72083) := X"00A21024";
        ram_buffer(72084) := X"00461025";
        ram_buffer(72085) := X"00031FC0";
        ram_buffer(72086) := X"00431825";
        ram_buffer(72087) := X"8FBF0024";
        ram_buffer(72088) := X"00602021";
        ram_buffer(72089) := X"8FB30020";
        ram_buffer(72090) := X"8FB2001C";
        ram_buffer(72091) := X"8FB10018";
        ram_buffer(72092) := X"8FB00014";
        ram_buffer(72093) := X"00E01821";
        ram_buffer(72094) := X"00801021";
        ram_buffer(72095) := X"03E00008";
        ram_buffer(72096) := X"27BD0028";
        ram_buffer(72097) := X"1480009E";
        ram_buffer(72098) := X"2463FFFF";
        ram_buffer(72099) := X"240307FF";
        ram_buffer(72100) := X"1623FFD9";
        ram_buffer(72101) := X"00A09021";
        ram_buffer(72102) := X"1000009F";
        ram_buffer(72103) := X"00451825";
        ram_buffer(72104) := X"1623FF5E";
        ram_buffer(72105) := X"28830039";
        ram_buffer(72106) := X"00451825";
        ram_buffer(72107) := X"1460FFD2";
        ram_buffer(72108) := X"00A09021";
        ram_buffer(72109) := X"02003021";
        ram_buffer(72110) := X"00003821";
        ram_buffer(72111) := X"00C08021";
        ram_buffer(72112) := X"00671025";
        ram_buffer(72113) := X"10400039";
        ram_buffer(72114) := X"00000000";
        ram_buffer(72115) := X"3C050007";
        ram_buffer(72116) := X"34A5FFFF";
        ram_buffer(72117) := X"00651024";
        ram_buffer(72118) := X"00471825";
        ram_buffer(72119) := X"1460003C";
        ram_buffer(72120) := X"00000000";
        ram_buffer(72121) := X"00001821";
        ram_buffer(72122) := X"240207FF";
        ram_buffer(72123) := X"1000FFD4";
        ram_buffer(72124) := X"2407FFFF";
        ram_buffer(72125) := X"02441825";
        ram_buffer(72126) := X"10600133";
        ram_buffer(72127) := X"00003821";
        ram_buffer(72128) := X"00801021";
        ram_buffer(72129) := X"32430007";
        ram_buffer(72130) := X"1460FF7A";
        ram_buffer(72131) := X"00021F40";
        ram_buffer(72132) := X"1000FF85";
        ram_buffer(72133) := X"001238C2";
        ram_buffer(72134) := X"14800058";
        ram_buffer(72135) := X"26230001";
        ram_buffer(72136) := X"306307FF";
        ram_buffer(72137) := X"28630002";
        ram_buffer(72138) := X"146000A5";
        ram_buffer(72139) := X"00A79023";
        ram_buffer(72140) := X"00B2182B";
        ram_buffer(72141) := X"00489823";
        ram_buffer(72142) := X"02639823";
        ram_buffer(72143) := X"3C030080";
        ram_buffer(72144) := X"02631824";
        ram_buffer(72145) := X"10600069";
        ram_buffer(72146) := X"02531825";
        ram_buffer(72147) := X"00E59023";
        ram_buffer(72148) := X"01021023";
        ram_buffer(72149) := X"00F2382B";
        ram_buffer(72150) := X"00479823";
        ram_buffer(72151) := X"1660FF47";
        ram_buffer(72152) := X"00C08021";
        ram_buffer(72153) := X"0C031D29";
        ram_buffer(72154) := X"02402021";
        ram_buffer(72155) := X"24420020";
        ram_buffer(72156) := X"2446FFF8";
        ram_buffer(72157) := X"28C30020";
        ram_buffer(72158) := X"1460FF47";
        ram_buffer(72159) := X"00061823";
        ram_buffer(72160) := X"2442FFD8";
        ram_buffer(72161) := X"00529804";
        ram_buffer(72162) := X"00D1102A";
        ram_buffer(72163) := X"1040FF48";
        ram_buffer(72164) := X"00009021";
        ram_buffer(72165) := X"3C02FF7F";
        ram_buffer(72166) := X"3442FFFF";
        ram_buffer(72167) := X"02268823";
        ram_buffer(72168) := X"02621024";
        ram_buffer(72169) := X"1000FF51";
        ram_buffer(72170) := X"32430007";
        ram_buffer(72171) := X"32030001";
        ram_buffer(72172) := X"240207FF";
        ram_buffer(72173) := X"00002821";
        ram_buffer(72174) := X"1000FFA1";
        ram_buffer(72175) := X"00003821";
        ram_buffer(72176) := X"01073825";
        ram_buffer(72177) := X"0007382B";
        ram_buffer(72178) := X"1000FF20";
        ram_buffer(72179) := X"00004021";
        ram_buffer(72180) := X"00402821";
        ram_buffer(72181) := X"32030001";
        ram_buffer(72182) := X"1000FF99";
        ram_buffer(72183) := X"240207FF";
        ram_buffer(72184) := X"1460008D";
        ram_buffer(72185) := X"26240001";
        ram_buffer(72186) := X"308307FF";
        ram_buffer(72187) := X"28630002";
        ram_buffer(72188) := X"1460006A";
        ram_buffer(72189) := X"00000000";
        ram_buffer(72190) := X"240307FF";
        ram_buffer(72191) := X"10830079";
        ram_buffer(72192) := X"00481021";
        ram_buffer(72193) := X"00A73821";
        ram_buffer(72194) := X"00E5282B";
        ram_buffer(72195) := X"00A21021";
        ram_buffer(72196) := X"000297C0";
        ram_buffer(72197) := X"00073842";
        ram_buffer(72198) := X"02479025";
        ram_buffer(72199) := X"00021042";
        ram_buffer(72200) := X"32430007";
        ram_buffer(72201) := X"1000FF31";
        ram_buffer(72202) := X"00808821";
        ram_buffer(72203) := X"24C6FFE1";
        ram_buffer(72204) := X"10430056";
        ram_buffer(72205) := X"00D33006";
        ram_buffer(72206) := X"00023823";
        ram_buffer(72207) := X"00F33804";
        ram_buffer(72208) := X"02473825";
        ram_buffer(72209) := X"0007382B";
        ram_buffer(72210) := X"00C79025";
        ram_buffer(72211) := X"00001021";
        ram_buffer(72212) := X"1000FFAC";
        ram_buffer(72213) := X"00008821";
        ram_buffer(72214) := X"1086004E";
        ram_buffer(72215) := X"00881806";
        ram_buffer(72216) := X"00042023";
        ram_buffer(72217) := X"00884004";
        ram_buffer(72218) := X"01073825";
        ram_buffer(72219) := X"0007382B";
        ram_buffer(72220) := X"00673825";
        ram_buffer(72221) := X"1000FEF5";
        ram_buffer(72222) := X"00004021";
        ram_buffer(72223) := X"12200036";
        ram_buffer(72224) := X"00451825";
        ram_buffer(72225) := X"240307FF";
        ram_buffer(72226) := X"114300C5";
        ram_buffer(72227) := X"3C030080";
        ram_buffer(72228) := X"00042023";
        ram_buffer(72229) := X"00431025";
        ram_buffer(72230) := X"28830039";
        ram_buffer(72231) := X"1060007E";
        ram_buffer(72232) := X"28830020";
        ram_buffer(72233) := X"106000CA";
        ram_buffer(72234) := X"24030020";
        ram_buffer(72235) := X"24090020";
        ram_buffer(72236) := X"01244823";
        ram_buffer(72237) := X"00859006";
        ram_buffer(72238) := X"01221804";
        ram_buffer(72239) := X"01252804";
        ram_buffer(72240) := X"00721825";
        ram_buffer(72241) := X"0005902B";
        ram_buffer(72242) := X"00729025";
        ram_buffer(72243) := X"00821006";
        ram_buffer(72244) := X"00F29023";
        ram_buffer(72245) := X"01021023";
        ram_buffer(72246) := X"00F2382B";
        ram_buffer(72247) := X"00471023";
        ram_buffer(72248) := X"01408821";
        ram_buffer(72249) := X"1000FEDD";
        ram_buffer(72250) := X"00C08021";
        ram_buffer(72251) := X"1460FEE1";
        ram_buffer(72252) := X"00003821";
        ram_buffer(72253) := X"00008021";
        ram_buffer(72254) := X"1000FF10";
        ram_buffer(72255) := X"00008821";
        ram_buffer(72256) := X"1060001E";
        ram_buffer(72257) := X"00A79021";
        ram_buffer(72258) := X"240407FF";
        ram_buffer(72259) := X"1624FF1B";
        ram_buffer(72260) := X"28640039";
        ram_buffer(72261) := X"00451825";
        ram_buffer(72262) := X"1460FF37";
        ram_buffer(72263) := X"00A09021";
        ram_buffer(72264) := X"00003821";
        ram_buffer(72265) := X"1000FF66";
        ram_buffer(72266) := X"00C08021";
        ram_buffer(72267) := X"10800031";
        ram_buffer(72268) := X"24090020";
        ram_buffer(72269) := X"01234823";
        ram_buffer(72270) := X"01282004";
        ram_buffer(72271) := X"00679006";
        ram_buffer(72272) := X"01273804";
        ram_buffer(72273) := X"00922025";
        ram_buffer(72274) := X"0007382B";
        ram_buffer(72275) := X"00873825";
        ram_buffer(72276) := X"1000FF0F";
        ram_buffer(72277) := X"00684006";
        ram_buffer(72278) := X"1460004A";
        ram_buffer(72279) := X"00000000";
        ram_buffer(72280) := X"240207FF";
        ram_buffer(72281) := X"1142008E";
        ram_buffer(72282) := X"01001021";
        ram_buffer(72283) := X"00E09021";
        ram_buffer(72284) := X"01408821";
        ram_buffer(72285) := X"1000FF20";
        ram_buffer(72286) := X"00C08021";
        ram_buffer(72287) := X"00481021";
        ram_buffer(72288) := X"0245282B";
        ram_buffer(72289) := X"1000FF06";
        ram_buffer(72290) := X"00A21021";
        ram_buffer(72291) := X"1000FFAC";
        ram_buffer(72292) := X"00003821";
        ram_buffer(72293) := X"1000FFB4";
        ram_buffer(72294) := X"00004021";
        ram_buffer(72295) := X"1620006A";
        ram_buffer(72296) := X"00451825";
        ram_buffer(72297) := X"146000A4";
        ram_buffer(72298) := X"01071825";
        ram_buffer(72299) := X"01001021";
        ram_buffer(72300) := X"1000FF11";
        ram_buffer(72301) := X"00E09021";
        ram_buffer(72302) := X"1000FF52";
        ram_buffer(72303) := X"00C08021";
        ram_buffer(72304) := X"16200020";
        ram_buffer(72305) := X"00451825";
        ram_buffer(72306) := X"1460004F";
        ram_buffer(72307) := X"01071825";
        ram_buffer(72308) := X"1060007C";
        ram_buffer(72309) := X"00E09021";
        ram_buffer(72310) := X"01001021";
        ram_buffer(72311) := X"1000FF06";
        ram_buffer(72312) := X"00C08021";
        ram_buffer(72313) := X"00001821";
        ram_buffer(72314) := X"00003821";
        ram_buffer(72315) := X"1000FF34";
        ram_buffer(72316) := X"00C08021";
        ram_buffer(72317) := X"10690071";
        ram_buffer(72318) := X"00682006";
        ram_buffer(72319) := X"00031823";
        ram_buffer(72320) := X"00684004";
        ram_buffer(72321) := X"01073825";
        ram_buffer(72322) := X"0007382B";
        ram_buffer(72323) := X"00873825";
        ram_buffer(72324) := X"1000FEDF";
        ram_buffer(72325) := X"00004021";
        ram_buffer(72326) := X"16200023";
        ram_buffer(72327) := X"240407FF";
        ram_buffer(72328) := X"00452025";
        ram_buffer(72329) := X"14800073";
        ram_buffer(72330) := X"00031827";
        ram_buffer(72331) := X"240207FF";
        ram_buffer(72332) := X"11420098";
        ram_buffer(72333) := X"01001021";
        ram_buffer(72334) := X"00E09021";
        ram_buffer(72335) := X"1000FEEE";
        ram_buffer(72336) := X"01408821";
        ram_buffer(72337) := X"14600009";
        ram_buffer(72338) := X"00000000";
        ram_buffer(72339) := X"01071025";
        ram_buffer(72340) := X"10400070";
        ram_buffer(72341) := X"3C030007";
        ram_buffer(72342) := X"01001021";
        ram_buffer(72343) := X"00E09021";
        ram_buffer(72344) := X"00C08021";
        ram_buffer(72345) := X"1000FEE4";
        ram_buffer(72346) := X"241107FF";
        ram_buffer(72347) := X"01073825";
        ram_buffer(72348) := X"14E0003B";
        ram_buffer(72349) := X"000220C2";
        ram_buffer(72350) := X"00A09021";
        ram_buffer(72351) := X"1000FEDE";
        ram_buffer(72352) := X"241107FF";
        ram_buffer(72353) := X"00042027";
        ram_buffer(72354) := X"14800043";
        ram_buffer(72355) := X"240307FF";
        ram_buffer(72356) := X"1000FF90";
        ram_buffer(72357) := X"00E59023";
        ram_buffer(72358) := X"00451025";
        ram_buffer(72359) := X"0002902B";
        ram_buffer(72360) := X"1000FF8B";
        ram_buffer(72361) := X"00001021";
        ram_buffer(72362) := X"1144007A";
        ram_buffer(72363) := X"3C040080";
        ram_buffer(72364) := X"00031823";
        ram_buffer(72365) := X"00441025";
        ram_buffer(72366) := X"28640039";
        ram_buffer(72367) := X"1080005A";
        ram_buffer(72368) := X"28640020";
        ram_buffer(72369) := X"10800078";
        ram_buffer(72370) := X"24040020";
        ram_buffer(72371) := X"24090020";
        ram_buffer(72372) := X"01234823";
        ram_buffer(72373) := X"00659006";
        ram_buffer(72374) := X"01222004";
        ram_buffer(72375) := X"01252804";
        ram_buffer(72376) := X"00922025";
        ram_buffer(72377) := X"0005902B";
        ram_buffer(72378) := X"00929025";
        ram_buffer(72379) := X"00621006";
        ram_buffer(72380) := X"02479021";
        ram_buffer(72381) := X"00484021";
        ram_buffer(72382) := X"0247382B";
        ram_buffer(72383) := X"00E81021";
        ram_buffer(72384) := X"1000FEA7";
        ram_buffer(72385) := X"01408821";
        ram_buffer(72386) := X"1060FEBB";
        ram_buffer(72387) := X"00A09021";
        ram_buffer(72388) := X"00A79023";
        ram_buffer(72389) := X"00481823";
        ram_buffer(72390) := X"00B2202B";
        ram_buffer(72391) := X"00642023";
        ram_buffer(72392) := X"3C030080";
        ram_buffer(72393) := X"00831824";
        ram_buffer(72394) := X"1060FEF2";
        ram_buffer(72395) := X"01021023";
        ram_buffer(72396) := X"00E59023";
        ram_buffer(72397) := X"00F2382B";
        ram_buffer(72398) := X"00471023";
        ram_buffer(72399) := X"32430007";
        ram_buffer(72400) := X"1000FE6A";
        ram_buffer(72401) := X"00C08021";
        ram_buffer(72402) := X"1460FFC8";
        ram_buffer(72403) := X"00000000";
        ram_buffer(72404) := X"01001021";
        ram_buffer(72405) := X"00E09021";
        ram_buffer(72406) := X"1000FEA7";
        ram_buffer(72407) := X"241107FF";
        ram_buffer(72408) := X"000818C2";
        ram_buffer(72409) := X"00641825";
        ram_buffer(72410) := X"3C060008";
        ram_buffer(72411) := X"00661824";
        ram_buffer(72412) := X"14600040";
        ram_buffer(72413) := X"000528C2";
        ram_buffer(72414) := X"00021740";
        ram_buffer(72415) := X"00453825";
        ram_buffer(72416) := X"000420C0";
        ram_buffer(72417) := X"00071742";
        ram_buffer(72418) := X"00441025";
        ram_buffer(72419) := X"000790C0";
        ram_buffer(72420) := X"1000FE99";
        ram_buffer(72421) := X"241107FF";
        ram_buffer(72422) := X"1543FF40";
        ram_buffer(72423) := X"28830039";
        ram_buffer(72424) := X"01071825";
        ram_buffer(72425) := X"1060FF5E";
        ram_buffer(72426) := X"01001021";
        ram_buffer(72427) := X"00E09021";
        ram_buffer(72428) := X"241107FF";
        ram_buffer(72429) := X"1000FE90";
        ram_buffer(72430) := X"00C08021";
        ram_buffer(72431) := X"1000FF91";
        ram_buffer(72432) := X"00004021";
        ram_buffer(72433) := X"00003821";
        ram_buffer(72434) := X"1000FE5C";
        ram_buffer(72435) := X"00008021";
        ram_buffer(72436) := X"1083003E";
        ram_buffer(72437) := X"00829006";
        ram_buffer(72438) := X"00042023";
        ram_buffer(72439) := X"00821004";
        ram_buffer(72440) := X"00452825";
        ram_buffer(72441) := X"0005102B";
        ram_buffer(72442) := X"02429025";
        ram_buffer(72443) := X"1000FF38";
        ram_buffer(72444) := X"00001021";
        ram_buffer(72445) := X"14600025";
        ram_buffer(72446) := X"240407FF";
        ram_buffer(72447) := X"00A79021";
        ram_buffer(72448) := X"00481021";
        ram_buffer(72449) := X"0247382B";
        ram_buffer(72450) := X"00E21021";
        ram_buffer(72451) := X"1000FE64";
        ram_buffer(72452) := X"01408821";
        ram_buffer(72453) := X"00003021";
        ram_buffer(72454) := X"3463FFFF";
        ram_buffer(72455) := X"2407FFFF";
        ram_buffer(72456) := X"1000FEA7";
        ram_buffer(72457) := X"00C08021";
        ram_buffer(72458) := X"00451025";
        ram_buffer(72459) := X"0002902B";
        ram_buffer(72460) := X"1000FFAF";
        ram_buffer(72461) := X"00001021";
        ram_buffer(72462) := X"1060FE6F";
        ram_buffer(72463) := X"00A09021";
        ram_buffer(72464) := X"00A79021";
        ram_buffer(72465) := X"00481021";
        ram_buffer(72466) := X"0245282B";
        ram_buffer(72467) := X"00A21021";
        ram_buffer(72468) := X"3C030080";
        ram_buffer(72469) := X"00431824";
        ram_buffer(72470) := X"1060FEAA";
        ram_buffer(72471) := X"3C03FF7F";
        ram_buffer(72472) := X"3463FFFF";
        ram_buffer(72473) := X"00431024";
        ram_buffer(72474) := X"24110001";
        ram_buffer(72475) := X"1000FE1F";
        ram_buffer(72476) := X"32430007";
        ram_buffer(72477) := X"3C02003F";
        ram_buffer(72478) := X"00008021";
        ram_buffer(72479) := X"241107FF";
        ram_buffer(72480) := X"3442FFFF";
        ram_buffer(72481) := X"1000FE26";
        ram_buffer(72482) := X"2412FFF8";
        ram_buffer(72483) := X"1544FF8B";
        ram_buffer(72484) := X"28640039";
        ram_buffer(72485) := X"01071825";
        ram_buffer(72486) := X"1460FFAE";
        ram_buffer(72487) := X"01001021";
        ram_buffer(72488) := X"1000FF20";
        ram_buffer(72489) := X"00003821";
        ram_buffer(72490) := X"1064000A";
        ram_buffer(72491) := X"00629006";
        ram_buffer(72492) := X"00031823";
        ram_buffer(72493) := X"00621004";
        ram_buffer(72494) := X"00452825";
        ram_buffer(72495) := X"0005102B";
        ram_buffer(72496) := X"02429025";
        ram_buffer(72497) := X"1000FF8A";
        ram_buffer(72498) := X"00001021";
        ram_buffer(72499) := X"1000FFC4";
        ram_buffer(72500) := X"00001021";
        ram_buffer(72501) := X"1000FFF8";
        ram_buffer(72502) := X"00001021";
        ram_buffer(72503) := X"00043502";
        ram_buffer(72504) := X"30C607FF";
        ram_buffer(72505) := X"3C03000F";
        ram_buffer(72506) := X"3463FFFF";
        ram_buffer(72507) := X"28C703FF";
        ram_buffer(72508) := X"00641824";
        ram_buffer(72509) := X"14E00015";
        ram_buffer(72510) := X"000427C2";
        ram_buffer(72511) := X"28C2041E";
        ram_buffer(72512) := X"1040000E";
        ram_buffer(72513) := X"24070433";
        ram_buffer(72514) := X"00E63823";
        ram_buffer(72515) := X"3C020010";
        ram_buffer(72516) := X"28E80020";
        ram_buffer(72517) := X"11000010";
        ram_buffer(72518) := X"00621825";
        ram_buffer(72519) := X"24C6FBED";
        ram_buffer(72520) := X"00E51006";
        ram_buffer(72521) := X"00C31804";
        ram_buffer(72522) := X"00621025";
        ram_buffer(72523) := X"10800008";
        ram_buffer(72524) := X"00000000";
        ram_buffer(72525) := X"03E00008";
        ram_buffer(72526) := X"00021023";
        ram_buffer(72527) := X"3C027FFF";
        ram_buffer(72528) := X"3442FFFF";
        ram_buffer(72529) := X"03E00008";
        ram_buffer(72530) := X"00821021";
        ram_buffer(72531) := X"00001021";
        ram_buffer(72532) := X"03E00008";
        ram_buffer(72533) := X"00000000";
        ram_buffer(72534) := X"24020413";
        ram_buffer(72535) := X"00461023";
        ram_buffer(72536) := X"1000FFF2";
        ram_buffer(72537) := X"00431006";
        ram_buffer(72538) := X"00041D02";
        ram_buffer(72539) := X"306607FF";
        ram_buffer(72540) := X"3C02000F";
        ram_buffer(72541) := X"3442FFFF";
        ram_buffer(72542) := X"28C303FF";
        ram_buffer(72543) := X"00441024";
        ram_buffer(72544) := X"14600008";
        ram_buffer(72545) := X"000427C2";
        ram_buffer(72546) := X"10800008";
        ram_buffer(72547) := X"28C3041F";
        ram_buffer(72548) := X"28C3041E";
        ram_buffer(72549) := X"14600003";
        ram_buffer(72550) := X"38840001";
        ram_buffer(72551) := X"03E00008";
        ram_buffer(72552) := X"00041023";
        ram_buffer(72553) := X"03E00008";
        ram_buffer(72554) := X"00001021";
        ram_buffer(72555) := X"1060FFFB";
        ram_buffer(72556) := X"38840001";
        ram_buffer(72557) := X"24040433";
        ram_buffer(72558) := X"00862023";
        ram_buffer(72559) := X"3C030010";
        ram_buffer(72560) := X"28870020";
        ram_buffer(72561) := X"14E00005";
        ram_buffer(72562) := X"00431025";
        ram_buffer(72563) := X"24030413";
        ram_buffer(72564) := X"00661823";
        ram_buffer(72565) := X"03E00008";
        ram_buffer(72566) := X"00621006";
        ram_buffer(72567) := X"24C3FBED";
        ram_buffer(72568) := X"00852806";
        ram_buffer(72569) := X"00621004";
        ram_buffer(72570) := X"03E00008";
        ram_buffer(72571) := X"00451025";
        ram_buffer(72572) := X"27BDFFE0";
        ram_buffer(72573) := X"AFBF001C";
        ram_buffer(72574) := X"AFB10018";
        ram_buffer(72575) := X"1080002C";
        ram_buffer(72576) := X"AFB00014";
        ram_buffer(72577) := X"00808021";
        ram_buffer(72578) := X"0480002E";
        ram_buffer(72579) := X"00048FC2";
        ram_buffer(72580) := X"0C031D29";
        ram_buffer(72581) := X"02002021";
        ram_buffer(72582) := X"2403041E";
        ram_buffer(72583) := X"00621823";
        ram_buffer(72584) := X"24050433";
        ram_buffer(72585) := X"00A32823";
        ram_buffer(72586) := X"28A40020";
        ram_buffer(72587) := X"14800018";
        ram_buffer(72588) := X"2404000B";
        ram_buffer(72589) := X"24020413";
        ram_buffer(72590) := X"00431023";
        ram_buffer(72591) := X"3C04000F";
        ram_buffer(72592) := X"00501004";
        ram_buffer(72593) := X"3484FFFF";
        ram_buffer(72594) := X"00441024";
        ram_buffer(72595) := X"00008021";
        ram_buffer(72596) := X"306407FF";
        ram_buffer(72597) := X"3C03000F";
        ram_buffer(72598) := X"3463FFFF";
        ram_buffer(72599) := X"00042500";
        ram_buffer(72600) := X"00431024";
        ram_buffer(72601) := X"00441025";
        ram_buffer(72602) := X"00111FC0";
        ram_buffer(72603) := X"00431825";
        ram_buffer(72604) := X"8FBF001C";
        ram_buffer(72605) := X"00602021";
        ram_buffer(72606) := X"8FB10018";
        ram_buffer(72607) := X"02001821";
        ram_buffer(72608) := X"00801021";
        ram_buffer(72609) := X"8FB00014";
        ram_buffer(72610) := X"03E00008";
        ram_buffer(72611) := X"27BD0020";
        ram_buffer(72612) := X"00821023";
        ram_buffer(72613) := X"3C04000F";
        ram_buffer(72614) := X"00501006";
        ram_buffer(72615) := X"3484FFFF";
        ram_buffer(72616) := X"00441024";
        ram_buffer(72617) := X"00B08004";
        ram_buffer(72618) := X"1000FFEA";
        ram_buffer(72619) := X"306407FF";
        ram_buffer(72620) := X"00008821";
        ram_buffer(72621) := X"00002021";
        ram_buffer(72622) := X"00001021";
        ram_buffer(72623) := X"1000FFE5";
        ram_buffer(72624) := X"00008021";
        ram_buffer(72625) := X"00048023";
        ram_buffer(72626) := X"0C031D29";
        ram_buffer(72627) := X"02002021";
        ram_buffer(72628) := X"2403041E";
        ram_buffer(72629) := X"00621823";
        ram_buffer(72630) := X"24050433";
        ram_buffer(72631) := X"00A32823";
        ram_buffer(72632) := X"28A40020";
        ram_buffer(72633) := X"1080FFD3";
        ram_buffer(72634) := X"2404000B";
        ram_buffer(72635) := X"1000FFE9";
        ram_buffer(72636) := X"00821023";
        ram_buffer(72637) := X"27BDFFE8";
        ram_buffer(72638) := X"AFB00010";
        ram_buffer(72639) := X"AFBF0014";
        ram_buffer(72640) := X"10800031";
        ram_buffer(72641) := X"00808021";
        ram_buffer(72642) := X"0C031D29";
        ram_buffer(72643) := X"00000000";
        ram_buffer(72644) := X"2403041E";
        ram_buffer(72645) := X"00621823";
        ram_buffer(72646) := X"24050433";
        ram_buffer(72647) := X"00A32823";
        ram_buffer(72648) := X"28A40020";
        ram_buffer(72649) := X"14800015";
        ram_buffer(72650) := X"2404000B";
        ram_buffer(72651) := X"24020413";
        ram_buffer(72652) := X"00431023";
        ram_buffer(72653) := X"3C04000F";
        ram_buffer(72654) := X"00501004";
        ram_buffer(72655) := X"3484FFFF";
        ram_buffer(72656) := X"306307FF";
        ram_buffer(72657) := X"00441024";
        ram_buffer(72658) := X"00032500";
        ram_buffer(72659) := X"3C03000F";
        ram_buffer(72660) := X"3463FFFF";
        ram_buffer(72661) := X"00431024";
        ram_buffer(72662) := X"00441825";
        ram_buffer(72663) := X"8FBF0014";
        ram_buffer(72664) := X"00008021";
        ram_buffer(72665) := X"00602021";
        ram_buffer(72666) := X"00801021";
        ram_buffer(72667) := X"02001821";
        ram_buffer(72668) := X"8FB00010";
        ram_buffer(72669) := X"03E00008";
        ram_buffer(72670) := X"27BD0018";
        ram_buffer(72671) := X"00821023";
        ram_buffer(72672) := X"00502006";
        ram_buffer(72673) := X"3C02000F";
        ram_buffer(72674) := X"306307FF";
        ram_buffer(72675) := X"3442FFFF";
        ram_buffer(72676) := X"00821024";
        ram_buffer(72677) := X"00032500";
        ram_buffer(72678) := X"3C03000F";
        ram_buffer(72679) := X"3463FFFF";
        ram_buffer(72680) := X"00431024";
        ram_buffer(72681) := X"00441825";
        ram_buffer(72682) := X"8FBF0014";
        ram_buffer(72683) := X"00B08004";
        ram_buffer(72684) := X"00602021";
        ram_buffer(72685) := X"00801021";
        ram_buffer(72686) := X"02001821";
        ram_buffer(72687) := X"8FB00010";
        ram_buffer(72688) := X"03E00008";
        ram_buffer(72689) := X"27BD0018";
        ram_buffer(72690) := X"00001821";
        ram_buffer(72691) := X"00032500";
        ram_buffer(72692) := X"3C03000F";
        ram_buffer(72693) := X"3463FFFF";
        ram_buffer(72694) := X"00001021";
        ram_buffer(72695) := X"00431024";
        ram_buffer(72696) := X"00441825";
        ram_buffer(72697) := X"8FBF0014";
        ram_buffer(72698) := X"00602021";
        ram_buffer(72699) := X"00801021";
        ram_buffer(72700) := X"02001821";
        ram_buffer(72701) := X"8FB00010";
        ram_buffer(72702) := X"03E00008";
        ram_buffer(72703) := X"27BD0018";
        ram_buffer(72704) := X"00851825";
        ram_buffer(72705) := X"1060005D";
        ram_buffer(72706) := X"3C02000F";
        ram_buffer(72707) := X"27BDFFE0";
        ram_buffer(72708) := X"AFB20018";
        ram_buffer(72709) := X"AFB10014";
        ram_buffer(72710) := X"AFB00010";
        ram_buffer(72711) := X"AFBF001C";
        ram_buffer(72712) := X"00A08021";
        ram_buffer(72713) := X"00808821";
        ram_buffer(72714) := X"10800019";
        ram_buffer(72715) := X"00809021";
        ram_buffer(72716) := X"0C031D29";
        ram_buffer(72717) := X"00000000";
        ram_buffer(72718) := X"2407043E";
        ram_buffer(72719) := X"00E23823";
        ram_buffer(72720) := X"28E50434";
        ram_buffer(72721) := X"10A0001B";
        ram_buffer(72722) := X"28E30437";
        ram_buffer(72723) := X"24080433";
        ram_buffer(72724) := X"01074023";
        ram_buffer(72725) := X"1100007B";
        ram_buffer(72726) := X"02002821";
        ram_buffer(72727) := X"29030020";
        ram_buffer(72728) := X"10600063";
        ram_buffer(72729) := X"2406002B";
        ram_buffer(72730) := X"00C21023";
        ram_buffer(72731) := X"01112004";
        ram_buffer(72732) := X"00503006";
        ram_buffer(72733) := X"00C41025";
        ram_buffer(72734) := X"3C04000F";
        ram_buffer(72735) := X"3484FFFF";
        ram_buffer(72736) := X"01102804";
        ram_buffer(72737) := X"00442024";
        ram_buffer(72738) := X"1000002F";
        ram_buffer(72739) := X"30E707FF";
        ram_buffer(72740) := X"0C031D29";
        ram_buffer(72741) := X"00A02021";
        ram_buffer(72742) := X"24420020";
        ram_buffer(72743) := X"2407043E";
        ram_buffer(72744) := X"00E23823";
        ram_buffer(72745) := X"28E50434";
        ram_buffer(72746) := X"14A0FFE9";
        ram_buffer(72747) := X"24080433";
        ram_buffer(72748) := X"28E30437";
        ram_buffer(72749) := X"1060003B";
        ram_buffer(72750) := X"24060436";
        ram_buffer(72751) := X"00C73023";
        ram_buffer(72752) := X"10C00007";
        ram_buffer(72753) := X"02002821";
        ram_buffer(72754) := X"24120028";
        ram_buffer(72755) := X"02429023";
        ram_buffer(72756) := X"02454006";
        ram_buffer(72757) := X"00D11804";
        ram_buffer(72758) := X"01039025";
        ram_buffer(72759) := X"00C52804";
        ram_buffer(72760) := X"3C03FF7F";
        ram_buffer(72761) := X"3463FFFF";
        ram_buffer(72762) := X"30A40007";
        ram_buffer(72763) := X"10800008";
        ram_buffer(72764) := X"02431824";
        ram_buffer(72765) := X"30A4000F";
        ram_buffer(72766) := X"24060004";
        ram_buffer(72767) := X"10860004";
        ram_buffer(72768) := X"24A40004";
        ram_buffer(72769) := X"0085282B";
        ram_buffer(72770) := X"00651821";
        ram_buffer(72771) := X"00802821";
        ram_buffer(72772) := X"3C080080";
        ram_buffer(72773) := X"00684024";
        ram_buffer(72774) := X"11000005";
        ram_buffer(72775) := X"3C04FF7F";
        ram_buffer(72776) := X"3484FFFF";
        ram_buffer(72777) := X"2407043F";
        ram_buffer(72778) := X"00641824";
        ram_buffer(72779) := X"00E23823";
        ram_buffer(72780) := X"00031740";
        ram_buffer(72781) := X"000528C2";
        ram_buffer(72782) := X"00031A40";
        ram_buffer(72783) := X"00452825";
        ram_buffer(72784) := X"00032302";
        ram_buffer(72785) := X"30E707FF";
        ram_buffer(72786) := X"3C02000F";
        ram_buffer(72787) := X"3442FFFF";
        ram_buffer(72788) := X"00822024";
        ram_buffer(72789) := X"8FBF001C";
        ram_buffer(72790) := X"00073D00";
        ram_buffer(72791) := X"00872025";
        ram_buffer(72792) := X"8FB20018";
        ram_buffer(72793) := X"8FB10014";
        ram_buffer(72794) := X"8FB00010";
        ram_buffer(72795) := X"00801021";
        ram_buffer(72796) := X"00A01821";
        ram_buffer(72797) := X"03E00008";
        ram_buffer(72798) := X"27BD0020";
        ram_buffer(72799) := X"3442FFFF";
        ram_buffer(72800) := X"00003821";
        ram_buffer(72801) := X"00002021";
        ram_buffer(72802) := X"00073D00";
        ram_buffer(72803) := X"00822024";
        ram_buffer(72804) := X"00002821";
        ram_buffer(72805) := X"00872025";
        ram_buffer(72806) := X"00801021";
        ram_buffer(72807) := X"03E00008";
        ram_buffer(72808) := X"00A01821";
        ram_buffer(72809) := X"24030008";
        ram_buffer(72810) := X"00621823";
        ram_buffer(72811) := X"30640020";
        ram_buffer(72812) := X"1080001E";
        ram_buffer(72813) := X"00032827";
        ram_buffer(72814) := X"00712806";
        ram_buffer(72815) := X"00001821";
        ram_buffer(72816) := X"24080476";
        ram_buffer(72817) := X"01074023";
        ram_buffer(72818) := X"31040020";
        ram_buffer(72819) := X"10800011";
        ram_buffer(72820) := X"00102042";
        ram_buffer(72821) := X"01102004";
        ram_buffer(72822) := X"00008021";
        ram_buffer(72823) := X"00908025";
        ram_buffer(72824) := X"0010802B";
        ram_buffer(72825) := X"00B02825";
        ram_buffer(72826) := X"1000FFBD";
        ram_buffer(72827) := X"00609021";
        ram_buffer(72828) := X"24020413";
        ram_buffer(72829) := X"00471023";
        ram_buffer(72830) := X"00502004";
        ram_buffer(72831) := X"3C02000F";
        ram_buffer(72832) := X"3442FFFF";
        ram_buffer(72833) := X"00822024";
        ram_buffer(72834) := X"30E707FF";
        ram_buffer(72835) := X"1000FFCE";
        ram_buffer(72836) := X"00002821";
        ram_buffer(72837) := X"00083027";
        ram_buffer(72838) := X"00C43006";
        ram_buffer(72839) := X"01112004";
        ram_buffer(72840) := X"00C42025";
        ram_buffer(72841) := X"1000FFED";
        ram_buffer(72842) := X"01108004";
        ram_buffer(72843) := X"00112040";
        ram_buffer(72844) := X"00A42004";
        ram_buffer(72845) := X"00702806";
        ram_buffer(72846) := X"00852825";
        ram_buffer(72847) := X"1000FFE0";
        ram_buffer(72848) := X"00711806";
        ram_buffer(72849) := X"3C06000F";
        ram_buffer(72850) := X"34C6FFFF";
        ram_buffer(72851) := X"02262024";
        ram_buffer(72852) := X"1000FFBD";
        ram_buffer(72853) := X"30E707FF";
        ram_buffer(72854) := X"00043D02";
        ram_buffer(72855) := X"30E707FF";
        ram_buffer(72856) := X"3C02000F";
        ram_buffer(72857) := X"24E60001";
        ram_buffer(72858) := X"3442FFFF";
        ram_buffer(72859) := X"00441024";
        ram_buffer(72860) := X"30C607FF";
        ram_buffer(72861) := X"000427C2";
        ram_buffer(72862) := X"000210C0";
        ram_buffer(72863) := X"00051F42";
        ram_buffer(72864) := X"28C60002";
        ram_buffer(72865) := X"00804021";
        ram_buffer(72866) := X"00621825";
        ram_buffer(72867) := X"14C0003D";
        ram_buffer(72868) := X"000548C0";
        ram_buffer(72869) := X"24E2FC80";
        ram_buffer(72870) := X"284600FF";
        ram_buffer(72871) := X"10C00049";
        ram_buffer(72872) := X"00000000";
        ram_buffer(72873) := X"1840001E";
        ram_buffer(72874) := X"00053180";
        ram_buffer(72875) := X"0006302B";
        ram_buffer(72876) := X"000318C0";
        ram_buffer(72877) := X"00C31825";
        ram_buffer(72878) := X"00092F42";
        ram_buffer(72879) := X"00652825";
        ram_buffer(72880) := X"30A30007";
        ram_buffer(72881) := X"10600005";
        ram_buffer(72882) := X"30A3000F";
        ram_buffer(72883) := X"24060004";
        ram_buffer(72884) := X"10660003";
        ram_buffer(72885) := X"3C030400";
        ram_buffer(72886) := X"24A50004";
        ram_buffer(72887) := X"3C030400";
        ram_buffer(72888) := X"00A31824";
        ram_buffer(72889) := X"10600013";
        ram_buffer(72890) := X"240300FF";
        ram_buffer(72891) := X"24420001";
        ram_buffer(72892) := X"10430034";
        ram_buffer(72893) := X"00052980";
        ram_buffer(72894) := X"00052A42";
        ram_buffer(72895) := X"304200FF";
        ram_buffer(72896) := X"00021DC0";
        ram_buffer(72897) := X"3C02007F";
        ram_buffer(72898) := X"3442FFFF";
        ram_buffer(72899) := X"00A22824";
        ram_buffer(72900) := X"00A32825";
        ram_buffer(72901) := X"000417C0";
        ram_buffer(72902) := X"03E00008";
        ram_buffer(72903) := X"00A21025";
        ram_buffer(72904) := X"2845FFE9";
        ram_buffer(72905) := X"10A00041";
        ram_buffer(72906) := X"240A001E";
        ram_buffer(72907) := X"00001021";
        ram_buffer(72908) := X"24050005";
        ram_buffer(72909) := X"240300FF";
        ram_buffer(72910) := X"14430016";
        ram_buffer(72911) := X"000528C2";
        ram_buffer(72912) := X"10A00020";
        ram_buffer(72913) := X"3C03003F";
        ram_buffer(72914) := X"3463FFFF";
        ram_buffer(72915) := X"00A32824";
        ram_buffer(72916) := X"14A00034";
        ram_buffer(72917) := X"01002021";
        ram_buffer(72918) := X"240200FF";
        ram_buffer(72919) := X"00602821";
        ram_buffer(72920) := X"00021DC0";
        ram_buffer(72921) := X"3C02007F";
        ram_buffer(72922) := X"3442FFFF";
        ram_buffer(72923) := X"00002021";
        ram_buffer(72924) := X"00A22824";
        ram_buffer(72925) := X"00A32825";
        ram_buffer(72926) := X"000417C0";
        ram_buffer(72927) := X"03E00008";
        ram_buffer(72928) := X"00A21025";
        ram_buffer(72929) := X"14E00019";
        ram_buffer(72930) := X"00692825";
        ram_buffer(72931) := X"14A0FFE8";
        ram_buffer(72932) := X"00001021";
        ram_buffer(72933) := X"3C03007F";
        ram_buffer(72934) := X"3463FFFF";
        ram_buffer(72935) := X"304200FF";
        ram_buffer(72936) := X"00A32824";
        ram_buffer(72937) := X"00021DC0";
        ram_buffer(72938) := X"3C02007F";
        ram_buffer(72939) := X"3442FFFF";
        ram_buffer(72940) := X"00A22824";
        ram_buffer(72941) := X"00A32825";
        ram_buffer(72942) := X"000417C0";
        ram_buffer(72943) := X"03E00008";
        ram_buffer(72944) := X"00A21025";
        ram_buffer(72945) := X"240200FF";
        ram_buffer(72946) := X"00021DC0";
        ram_buffer(72947) := X"3C02007F";
        ram_buffer(72948) := X"3442FFFF";
        ram_buffer(72949) := X"00002821";
        ram_buffer(72950) := X"00A22824";
        ram_buffer(72951) := X"00A32825";
        ram_buffer(72952) := X"000417C0";
        ram_buffer(72953) := X"03E00008";
        ram_buffer(72954) := X"00A21025";
        ram_buffer(72955) := X"00691025";
        ram_buffer(72956) := X"1040FFF4";
        ram_buffer(72957) := X"000318C0";
        ram_buffer(72958) := X"00092F42";
        ram_buffer(72959) := X"00A32825";
        ram_buffer(72960) := X"3C0301FF";
        ram_buffer(72961) := X"3463FFF8";
        ram_buffer(72962) := X"00A32824";
        ram_buffer(72963) := X"14A00015";
        ram_buffer(72964) := X"00000000";
        ram_buffer(72965) := X"3C05003F";
        ram_buffer(72966) := X"00004021";
        ram_buffer(72967) := X"34A5FFFF";
        ram_buffer(72968) := X"01002021";
        ram_buffer(72969) := X"1000FFB6";
        ram_buffer(72970) := X"240200FF";
        ram_buffer(72971) := X"01425023";
        ram_buffer(72972) := X"3C050080";
        ram_buffer(72973) := X"294B0020";
        ram_buffer(72974) := X"1160000C";
        ram_buffer(72975) := X"00651825";
        ram_buffer(72976) := X"24E6FC82";
        ram_buffer(72977) := X"00C93804";
        ram_buffer(72978) := X"0007382B";
        ram_buffer(72979) := X"00C31804";
        ram_buffer(72980) := X"00E33025";
        ram_buffer(72981) := X"01492806";
        ram_buffer(72982) := X"00C52825";
        ram_buffer(72983) := X"1000FF98";
        ram_buffer(72984) := X"00001021";
        ram_buffer(72985) := X"1000FF96";
        ram_buffer(72986) := X"240200FF";
        ram_buffer(72987) := X"2405FFFE";
        ram_buffer(72988) := X"00A22823";
        ram_buffer(72989) := X"24020020";
        ram_buffer(72990) := X"11420008";
        ram_buffer(72991) := X"00A32806";
        ram_buffer(72992) := X"24E7FCA2";
        ram_buffer(72993) := X"00E31804";
        ram_buffer(72994) := X"00691825";
        ram_buffer(72995) := X"0003182B";
        ram_buffer(72996) := X"00652825";
        ram_buffer(72997) := X"1000FF8A";
        ram_buffer(72998) := X"00001021";
        ram_buffer(72999) := X"1000FFFA";
        ram_buffer(73000) := X"00001821";
        ram_buffer(73001) := X"3C020001";
        ram_buffer(73002) := X"0082102B";
        ram_buffer(73003) := X"1040000C";
        ram_buffer(73004) := X"3C020100";
        ram_buffer(73005) := X"2C820100";
        ram_buffer(73006) := X"10400014";
        ram_buffer(73007) := X"3C03100D";
        ram_buffer(73008) := X"00001021";
        ram_buffer(73009) := X"00442006";
        ram_buffer(73010) := X"2463B660";
        ram_buffer(73011) := X"00832021";
        ram_buffer(73012) := X"90820000";
        ram_buffer(73013) := X"24050020";
        ram_buffer(73014) := X"03E00008";
        ram_buffer(73015) := X"00A21023";
        ram_buffer(73016) := X"0082102B";
        ram_buffer(73017) := X"14400011";
        ram_buffer(73018) := X"3C03100D";
        ram_buffer(73019) := X"24020018";
        ram_buffer(73020) := X"00442006";
        ram_buffer(73021) := X"2463B660";
        ram_buffer(73022) := X"00832021";
        ram_buffer(73023) := X"90820000";
        ram_buffer(73024) := X"24050008";
        ram_buffer(73025) := X"03E00008";
        ram_buffer(73026) := X"00A21023";
        ram_buffer(73027) := X"24020008";
        ram_buffer(73028) := X"00442006";
        ram_buffer(73029) := X"2463B660";
        ram_buffer(73030) := X"00832021";
        ram_buffer(73031) := X"90820000";
        ram_buffer(73032) := X"24050018";
        ram_buffer(73033) := X"03E00008";
        ram_buffer(73034) := X"00A21023";
        ram_buffer(73035) := X"24020010";
        ram_buffer(73036) := X"00442006";
        ram_buffer(73037) := X"2463B660";
        ram_buffer(73038) := X"00832021";
        ram_buffer(73039) := X"90820000";
        ram_buffer(73040) := X"24050010";
        ram_buffer(73041) := X"03E00008";
        ram_buffer(73042) := X"00A21023";
        ram_buffer(73043) := X"3C02100D";
        ram_buffer(73044) := X"8C42C7A0";
        ram_buffer(73045) := X"2403FFFF";
        ram_buffer(73046) := X"10430012";
        ram_buffer(73047) := X"00000000";
        ram_buffer(73048) := X"27BDFFE0";
        ram_buffer(73049) := X"AFB00014";
        ram_buffer(73050) := X"3C10100D";
        ram_buffer(73051) := X"AFB10018";
        ram_buffer(73052) := X"AFBF001C";
        ram_buffer(73053) := X"2610C7A0";
        ram_buffer(73054) := X"2411FFFF";
        ram_buffer(73055) := X"0040F809";
        ram_buffer(73056) := X"2610FFFC";
        ram_buffer(73057) := X"8E020000";
        ram_buffer(73058) := X"00000000";
        ram_buffer(73059) := X"1451FFFB";
        ram_buffer(73060) := X"00000000";
        ram_buffer(73061) := X"8FBF001C";
        ram_buffer(73062) := X"8FB10018";
        ram_buffer(73063) := X"8FB00014";
        ram_buffer(73064) := X"27BD0020";
        ram_buffer(73065) := X"03E00008";
        ram_buffer(73066) := X"00000000";
        ram_buffer(73067) := X"27BDFFE0";
        ram_buffer(73068) := X"AFBF0014";
        ram_buffer(73069) := X"04110001";
        ram_buffer(73070) := X"00000000";
        ram_buffer(73071) := X"0C020148";
        ram_buffer(73072) := X"00000000";
        ram_buffer(73073) := X"8FBF0014";
        ram_buffer(73074) := X"27BD0020";
        ram_buffer(73075) := X"03E00008";
        ram_buffer(73076) := X"00000000";
        ram_buffer(73077) := X"00000000";
        ram_buffer(73078) := X"75736167";
        ram_buffer(73079) := X"653A2025";
        ram_buffer(73080) := X"73205B73";
        ram_buffer(73081) := X"77697463";
        ram_buffer(73082) := X"6865735D";
        ram_buffer(73083) := X"20000000";
        ram_buffer(73084) := X"5B696E70";
        ram_buffer(73085) := X"75746669";
        ram_buffer(73086) := X"6C655D0A";
        ram_buffer(73087) := X"00000000";
        ram_buffer(73088) := X"53776974";
        ram_buffer(73089) := X"63686573";
        ram_buffer(73090) := X"20286E61";
        ram_buffer(73091) := X"6D657320";
        ram_buffer(73092) := X"6D617920";
        ram_buffer(73093) := X"62652061";
        ram_buffer(73094) := X"62627265";
        ram_buffer(73095) := X"76696174";
        ram_buffer(73096) := X"6564293A";
        ram_buffer(73097) := X"0A000000";
        ram_buffer(73098) := X"20202D71";
        ram_buffer(73099) := X"75616C69";
        ram_buffer(73100) := X"7479204E";
        ram_buffer(73101) := X"20202020";
        ram_buffer(73102) := X"20436F6D";
        ram_buffer(73103) := X"70726573";
        ram_buffer(73104) := X"73696F6E";
        ram_buffer(73105) := X"20717561";
        ram_buffer(73106) := X"6C697479";
        ram_buffer(73107) := X"2028302E";
        ram_buffer(73108) := X"2E313030";
        ram_buffer(73109) := X"3B20352D";
        ram_buffer(73110) := X"39352069";
        ram_buffer(73111) := X"73207573";
        ram_buffer(73112) := X"6566756C";
        ram_buffer(73113) := X"2072616E";
        ram_buffer(73114) := X"6765290A";
        ram_buffer(73115) := X"00000000";
        ram_buffer(73116) := X"20202D67";
        ram_buffer(73117) := X"72617973";
        ram_buffer(73118) := X"63616C65";
        ram_buffer(73119) := X"20202020";
        ram_buffer(73120) := X"20437265";
        ram_buffer(73121) := X"61746520";
        ram_buffer(73122) := X"6D6F6E6F";
        ram_buffer(73123) := X"6368726F";
        ram_buffer(73124) := X"6D65204A";
        ram_buffer(73125) := X"50454720";
        ram_buffer(73126) := X"66696C65";
        ram_buffer(73127) := X"0A000000";
        ram_buffer(73128) := X"20202D6F";
        ram_buffer(73129) := X"7074696D";
        ram_buffer(73130) := X"697A6520";
        ram_buffer(73131) := X"20202020";
        ram_buffer(73132) := X"204F7074";
        ram_buffer(73133) := X"696D697A";
        ram_buffer(73134) := X"65204875";
        ram_buffer(73135) := X"66666D61";
        ram_buffer(73136) := X"6E207461";
        ram_buffer(73137) := X"626C6520";
        ram_buffer(73138) := X"28736D61";
        ram_buffer(73139) := X"6C6C6572";
        ram_buffer(73140) := X"2066696C";
        ram_buffer(73141) := X"652C2062";
        ram_buffer(73142) := X"75742073";
        ram_buffer(73143) := X"6C6F7720";
        ram_buffer(73144) := X"636F6D70";
        ram_buffer(73145) := X"72657373";
        ram_buffer(73146) := X"696F6E29";
        ram_buffer(73147) := X"0A000000";
        ram_buffer(73148) := X"20202D70";
        ram_buffer(73149) := X"726F6772";
        ram_buffer(73150) := X"65737369";
        ram_buffer(73151) := X"76652020";
        ram_buffer(73152) := X"20437265";
        ram_buffer(73153) := X"61746520";
        ram_buffer(73154) := X"70726F67";
        ram_buffer(73155) := X"72657373";
        ram_buffer(73156) := X"69766520";
        ram_buffer(73157) := X"4A504547";
        ram_buffer(73158) := X"2066696C";
        ram_buffer(73159) := X"650A0000";
        ram_buffer(73160) := X"20202D74";
        ram_buffer(73161) := X"61726761";
        ram_buffer(73162) := X"20202020";
        ram_buffer(73163) := X"20202020";
        ram_buffer(73164) := X"20496E70";
        ram_buffer(73165) := X"75742066";
        ram_buffer(73166) := X"696C6520";
        ram_buffer(73167) := X"69732054";
        ram_buffer(73168) := X"61726761";
        ram_buffer(73169) := X"20666F72";
        ram_buffer(73170) := X"6D617420";
        ram_buffer(73171) := X"28757375";
        ram_buffer(73172) := X"616C6C79";
        ram_buffer(73173) := X"206E6F74";
        ram_buffer(73174) := X"206E6565";
        ram_buffer(73175) := X"64656429";
        ram_buffer(73176) := X"0A000000";
        ram_buffer(73177) := X"53776974";
        ram_buffer(73178) := X"63686573";
        ram_buffer(73179) := X"20666F72";
        ram_buffer(73180) := X"20616476";
        ram_buffer(73181) := X"616E6365";
        ram_buffer(73182) := X"64207573";
        ram_buffer(73183) := X"6572733A";
        ram_buffer(73184) := X"0A000000";
        ram_buffer(73185) := X"20286465";
        ram_buffer(73186) := X"6661756C";
        ram_buffer(73187) := X"74290000";
        ram_buffer(73188) := X"20202D64";
        ram_buffer(73189) := X"63742069";
        ram_buffer(73190) := X"6E742020";
        ram_buffer(73191) := X"20202020";
        ram_buffer(73192) := X"20557365";
        ram_buffer(73193) := X"20696E74";
        ram_buffer(73194) := X"65676572";
        ram_buffer(73195) := X"20444354";
        ram_buffer(73196) := X"206D6574";
        ram_buffer(73197) := X"686F6425";
        ram_buffer(73198) := X"730A0000";
        ram_buffer(73199) := X"20202D64";
        ram_buffer(73200) := X"63742066";
        ram_buffer(73201) := X"61737420";
        ram_buffer(73202) := X"20202020";
        ram_buffer(73203) := X"20557365";
        ram_buffer(73204) := X"20666173";
        ram_buffer(73205) := X"7420696E";
        ram_buffer(73206) := X"74656765";
        ram_buffer(73207) := X"72204443";
        ram_buffer(73208) := X"5420286C";
        ram_buffer(73209) := X"65737320";
        ram_buffer(73210) := X"61636375";
        ram_buffer(73211) := X"72617465";
        ram_buffer(73212) := X"2925730A";
        ram_buffer(73213) := X"00000000";
        ram_buffer(73214) := X"20202D64";
        ram_buffer(73215) := X"63742066";
        ram_buffer(73216) := X"6C6F6174";
        ram_buffer(73217) := X"20202020";
        ram_buffer(73218) := X"20557365";
        ram_buffer(73219) := X"20666C6F";
        ram_buffer(73220) := X"6174696E";
        ram_buffer(73221) := X"672D706F";
        ram_buffer(73222) := X"696E7420";
        ram_buffer(73223) := X"44435420";
        ram_buffer(73224) := X"6D657468";
        ram_buffer(73225) := X"6F642573";
        ram_buffer(73226) := X"0A000000";
        ram_buffer(73227) := X"20202D72";
        ram_buffer(73228) := X"65737461";
        ram_buffer(73229) := X"7274204E";
        ram_buffer(73230) := X"20202020";
        ram_buffer(73231) := X"20536574";
        ram_buffer(73232) := X"20726573";
        ram_buffer(73233) := X"74617274";
        ram_buffer(73234) := X"20696E74";
        ram_buffer(73235) := X"65727661";
        ram_buffer(73236) := X"6C20696E";
        ram_buffer(73237) := X"20726F77";
        ram_buffer(73238) := X"732C206F";
        ram_buffer(73239) := X"7220696E";
        ram_buffer(73240) := X"20626C6F";
        ram_buffer(73241) := X"636B7320";
        ram_buffer(73242) := X"77697468";
        ram_buffer(73243) := X"20420A00";
        ram_buffer(73244) := X"20202D73";
        ram_buffer(73245) := X"6D6F6F74";
        ram_buffer(73246) := X"68204E20";
        ram_buffer(73247) := X"20202020";
        ram_buffer(73248) := X"20536D6F";
        ram_buffer(73249) := X"6F746820";
        ram_buffer(73250) := X"64697468";
        ram_buffer(73251) := X"65726564";
        ram_buffer(73252) := X"20696E70";
        ram_buffer(73253) := X"75742028";
        ram_buffer(73254) := X"4E3D312E";
        ram_buffer(73255) := X"2E313030";
        ram_buffer(73256) := X"20697320";
        ram_buffer(73257) := X"73747265";
        ram_buffer(73258) := X"6E677468";
        ram_buffer(73259) := X"290A0000";
        ram_buffer(73260) := X"20202D6D";
        ram_buffer(73261) := X"61786D65";
        ram_buffer(73262) := X"6D6F7279";
        ram_buffer(73263) := X"204E2020";
        ram_buffer(73264) := X"204D6178";
        ram_buffer(73265) := X"696D756D";
        ram_buffer(73266) := X"206D656D";
        ram_buffer(73267) := X"6F727920";
        ram_buffer(73268) := X"746F2075";
        ram_buffer(73269) := X"73652028";
        ram_buffer(73270) := X"696E206B";
        ram_buffer(73271) := X"62797465";
        ram_buffer(73272) := X"73290A00";
        ram_buffer(73273) := X"20202D6F";
        ram_buffer(73274) := X"75746669";
        ram_buffer(73275) := X"6C65206E";
        ram_buffer(73276) := X"616D6520";
        ram_buffer(73277) := X"20537065";
        ram_buffer(73278) := X"63696679";
        ram_buffer(73279) := X"206E616D";
        ram_buffer(73280) := X"6520666F";
        ram_buffer(73281) := X"72206F75";
        ram_buffer(73282) := X"74707574";
        ram_buffer(73283) := X"2066696C";
        ram_buffer(73284) := X"650A0000";
        ram_buffer(73285) := X"20202D76";
        ram_buffer(73286) := X"6572626F";
        ram_buffer(73287) := X"73652020";
        ram_buffer(73288) := X"6F722020";
        ram_buffer(73289) := X"2D646562";
        ram_buffer(73290) := X"75672020";
        ram_buffer(73291) := X"20456D69";
        ram_buffer(73292) := X"74206465";
        ram_buffer(73293) := X"62756720";
        ram_buffer(73294) := X"6F757470";
        ram_buffer(73295) := X"75740A00";
        ram_buffer(73296) := X"53776974";
        ram_buffer(73297) := X"63686573";
        ram_buffer(73298) := X"20666F72";
        ram_buffer(73299) := X"2077697A";
        ram_buffer(73300) := X"61726473";
        ram_buffer(73301) := X"3A0A0000";
        ram_buffer(73302) := X"20202D62";
        ram_buffer(73303) := X"6173656C";
        ram_buffer(73304) := X"696E6520";
        ram_buffer(73305) := X"20202020";
        ram_buffer(73306) := X"20466F72";
        ram_buffer(73307) := X"63652062";
        ram_buffer(73308) := X"6173656C";
        ram_buffer(73309) := X"696E6520";
        ram_buffer(73310) := X"6F757470";
        ram_buffer(73311) := X"75740A00";
        ram_buffer(73312) := X"20202D71";
        ram_buffer(73313) := X"7461626C";
        ram_buffer(73314) := X"65732066";
        ram_buffer(73315) := X"696C6520";
        ram_buffer(73316) := X"20557365";
        ram_buffer(73317) := X"20717561";
        ram_buffer(73318) := X"6E74697A";
        ram_buffer(73319) := X"6174696F";
        ram_buffer(73320) := X"6E207461";
        ram_buffer(73321) := X"626C6573";
        ram_buffer(73322) := X"20676976";
        ram_buffer(73323) := X"656E2069";
        ram_buffer(73324) := X"6E206669";
        ram_buffer(73325) := X"6C650A00";
        ram_buffer(73326) := X"20202D71";
        ram_buffer(73327) := X"736C6F74";
        ram_buffer(73328) := X"73204E5B";
        ram_buffer(73329) := X"2C2E2E2E";
        ram_buffer(73330) := X"5D202020";
        ram_buffer(73331) := X"20536574";
        ram_buffer(73332) := X"20636F6D";
        ram_buffer(73333) := X"706F6E65";
        ram_buffer(73334) := X"6E742071";
        ram_buffer(73335) := X"75616E74";
        ram_buffer(73336) := X"697A6174";
        ram_buffer(73337) := X"696F6E20";
        ram_buffer(73338) := X"7461626C";
        ram_buffer(73339) := X"65730A00";
        ram_buffer(73340) := X"20202D73";
        ram_buffer(73341) := X"616D706C";
        ram_buffer(73342) := X"65204878";
        ram_buffer(73343) := X"565B2C2E";
        ram_buffer(73344) := X"2E2E5D20";
        ram_buffer(73345) := X"20536574";
        ram_buffer(73346) := X"20636F6D";
        ram_buffer(73347) := X"706F6E65";
        ram_buffer(73348) := X"6E742073";
        ram_buffer(73349) := X"616D706C";
        ram_buffer(73350) := X"696E6720";
        ram_buffer(73351) := X"66616374";
        ram_buffer(73352) := X"6F72730A";
        ram_buffer(73353) := X"00000000";
        ram_buffer(73354) := X"20202D73";
        ram_buffer(73355) := X"63616E73";
        ram_buffer(73356) := X"2066696C";
        ram_buffer(73357) := X"65202020";
        ram_buffer(73358) := X"20437265";
        ram_buffer(73359) := X"61746520";
        ram_buffer(73360) := X"6D756C74";
        ram_buffer(73361) := X"692D7363";
        ram_buffer(73362) := X"616E204A";
        ram_buffer(73363) := X"50454720";
        ram_buffer(73364) := X"70657220";
        ram_buffer(73365) := X"73637269";
        ram_buffer(73366) := X"70742066";
        ram_buffer(73367) := X"696C650A";
        ram_buffer(73368) := X"00000000";
        ram_buffer(73369) := X"61726974";
        ram_buffer(73370) := X"686D6574";
        ram_buffer(73371) := X"69630000";
        ram_buffer(73372) := X"25733A20";
        ram_buffer(73373) := X"736F7272";
        ram_buffer(73374) := X"792C2061";
        ram_buffer(73375) := X"72697468";
        ram_buffer(73376) := X"6D657469";
        ram_buffer(73377) := X"6320636F";
        ram_buffer(73378) := X"64696E67";
        ram_buffer(73379) := X"206E6F74";
        ram_buffer(73380) := X"20737570";
        ram_buffer(73381) := X"706F7274";
        ram_buffer(73382) := X"65640A00";
        ram_buffer(73383) := X"62617365";
        ram_buffer(73384) := X"6C696E65";
        ram_buffer(73385) := X"00000000";
        ram_buffer(73386) := X"64637400";
        ram_buffer(73387) := X"696E7400";
        ram_buffer(73388) := X"66617374";
        ram_buffer(73389) := X"00000000";
        ram_buffer(73390) := X"666C6F61";
        ram_buffer(73391) := X"74000000";
        ram_buffer(73392) := X"64656275";
        ram_buffer(73393) := X"67000000";
        ram_buffer(73394) := X"76657262";
        ram_buffer(73395) := X"6F736500";
        ram_buffer(73396) := X"436F7079";
        ram_buffer(73397) := X"72696768";
        ram_buffer(73398) := X"74202843";
        ram_buffer(73399) := X"29203139";
        ram_buffer(73400) := X"39362C20";
        ram_buffer(73401) := X"54686F6D";
        ram_buffer(73402) := X"61732047";
        ram_buffer(73403) := X"2E204C61";
        ram_buffer(73404) := X"6E650000";
        ram_buffer(73405) := X"36612020";
        ram_buffer(73406) := X"372D4665";
        ram_buffer(73407) := X"622D3936";
        ram_buffer(73408) := X"00000000";
        ram_buffer(73409) := X"496E6465";
        ram_buffer(73410) := X"70656E64";
        ram_buffer(73411) := X"656E7420";
        ram_buffer(73412) := X"4A504547";
        ram_buffer(73413) := X"2047726F";
        ram_buffer(73414) := X"75702773";
        ram_buffer(73415) := X"20434A50";
        ram_buffer(73416) := X"45472C20";
        ram_buffer(73417) := X"76657273";
        ram_buffer(73418) := X"696F6E20";
        ram_buffer(73419) := X"25730A25";
        ram_buffer(73420) := X"730A0000";
        ram_buffer(73421) := X"67726179";
        ram_buffer(73422) := X"7363616C";
        ram_buffer(73423) := X"65000000";
        ram_buffer(73424) := X"67726579";
        ram_buffer(73425) := X"7363616C";
        ram_buffer(73426) := X"65000000";
        ram_buffer(73427) := X"6D61786D";
        ram_buffer(73428) := X"656D6F72";
        ram_buffer(73429) := X"79000000";
        ram_buffer(73430) := X"256C6425";
        ram_buffer(73431) := X"63000000";
        ram_buffer(73432) := X"6F707469";
        ram_buffer(73433) := X"6D697A65";
        ram_buffer(73434) := X"00000000";
        ram_buffer(73435) := X"6F707469";
        ram_buffer(73436) := X"6D697365";
        ram_buffer(73437) := X"00000000";
        ram_buffer(73438) := X"6F757466";
        ram_buffer(73439) := X"696C6500";
        ram_buffer(73440) := X"70726F67";
        ram_buffer(73441) := X"72657373";
        ram_buffer(73442) := X"69766500";
        ram_buffer(73443) := X"7175616C";
        ram_buffer(73444) := X"69747900";
        ram_buffer(73445) := X"71736C6F";
        ram_buffer(73446) := X"74730000";
        ram_buffer(73447) := X"71746162";
        ram_buffer(73448) := X"6C657300";
        ram_buffer(73449) := X"72657374";
        ram_buffer(73450) := X"61727400";
        ram_buffer(73451) := X"73616D70";
        ram_buffer(73452) := X"6C650000";
        ram_buffer(73453) := X"7363616E";
        ram_buffer(73454) := X"73000000";
        ram_buffer(73455) := X"736D6F6F";
        ram_buffer(73456) := X"74680000";
        ram_buffer(73457) := X"74617267";
        ram_buffer(73458) := X"61000000";
        ram_buffer(73459) := X"636A7065";
        ram_buffer(73460) := X"67000000";
        ram_buffer(73461) := X"25733A20";
        ram_buffer(73462) := X"6F6E6C79";
        ram_buffer(73463) := X"206F6E65";
        ram_buffer(73464) := X"20696E70";
        ram_buffer(73465) := X"75742066";
        ram_buffer(73466) := X"696C650A";
        ram_buffer(73467) := X"00000000";
        ram_buffer(73468) := X"72620000";
        ram_buffer(73469) := X"25733A20";
        ram_buffer(73470) := X"63616E27";
        ram_buffer(73471) := X"74206F70";
        ram_buffer(73472) := X"656E2025";
        ram_buffer(73473) := X"730A0000";
        ram_buffer(73474) := X"77620000";
        ram_buffer(73475) := X"2D717561";
        ram_buffer(73476) := X"6C697479";
        ram_buffer(73477) := X"00000000";
        ram_buffer(73478) := X"39300000";
        ram_buffer(73479) := X"2D6F7574";
        ram_buffer(73480) := X"66696C65";
        ram_buffer(73481) := X"00000000";
        ram_buffer(73482) := X"4C656E6E";
        ram_buffer(73483) := X"61313630";
        ram_buffer(73484) := X"2E70706D";
        ram_buffer(73485) := X"00000000";
        ram_buffer(73486) := X"53746172";
        ram_buffer(73487) := X"74696E67";
        ram_buffer(73488) := X"204A5045";
        ram_buffer(73489) := X"4720636F";
        ram_buffer(73490) := X"6D707265";
        ram_buffer(73491) := X"7373696F";
        ram_buffer(73492) := X"6E000000";
        ram_buffer(73493) := X"2D2D2D2D";
        ram_buffer(73494) := X"2D2D2D2D";
        ram_buffer(73495) := X"2D2D2D2D";
        ram_buffer(73496) := X"2D2D2D2D";
        ram_buffer(73497) := X"2D2D2D2D";
        ram_buffer(73498) := X"2D2D2D2D";
        ram_buffer(73499) := X"2D2D2D2D";
        ram_buffer(73500) := X"2D2D2D2D";
        ram_buffer(73501) := X"2D2D2D2D";
        ram_buffer(73502) := X"2D2D2D2D";
        ram_buffer(73503) := X"2D2D2D2D";
        ram_buffer(73504) := X"2D2D2D2D";
        ram_buffer(73505) := X"2D2D2D2D";
        ram_buffer(73506) := X"2D2D2D2D";
        ram_buffer(73507) := X"2D2D0000";
        ram_buffer(73508) := X"434A5045";
        ram_buffer(73509) := X"4720746F";
        ram_buffer(73510) := X"6F6B2025";
        ram_buffer(73511) := X"272E366C";
        ram_buffer(73512) := X"66206D69";
        ram_buffer(73513) := X"6C6C696F";
        ram_buffer(73514) := X"6E20636C";
        ram_buffer(73515) := X"6F636B20";
        ram_buffer(73516) := X"6379636C";
        ram_buffer(73517) := X"65730A00";
        ram_buffer(73518) := X"25630A00";
        ram_buffer(73519) := X"4C656E6E";
        ram_buffer(73520) := X"61313630";
        ram_buffer(73521) := X"2E6A7067";
        ram_buffer(73522) := X"00000000";
        ram_buffer(73523) := X"4C656E6E";
        ram_buffer(73524) := X"61313630";
        ram_buffer(73525) := X"676F6C64";
        ram_buffer(73526) := X"656E2E6A";
        ram_buffer(73527) := X"70670000";
        ram_buffer(73528) := X"556E7375";
        ram_buffer(73529) := X"70706F72";
        ram_buffer(73530) := X"74656420";
        ram_buffer(73531) := X"424D5020";
        ram_buffer(73532) := X"636F6C6F";
        ram_buffer(73533) := X"726D6170";
        ram_buffer(73534) := X"20666F72";
        ram_buffer(73535) := X"6D617400";
        ram_buffer(73536) := X"4F6E6C79";
        ram_buffer(73537) := X"20382D20";
        ram_buffer(73538) := X"616E6420";
        ram_buffer(73539) := X"32342D62";
        ram_buffer(73540) := X"69742042";
        ram_buffer(73541) := X"4D502066";
        ram_buffer(73542) := X"696C6573";
        ram_buffer(73543) := X"20617265";
        ram_buffer(73544) := X"20737570";
        ram_buffer(73545) := X"706F7274";
        ram_buffer(73546) := X"65640000";
        ram_buffer(73547) := X"496E7661";
        ram_buffer(73548) := X"6C696420";
        ram_buffer(73549) := X"424D5020";
        ram_buffer(73550) := X"66696C65";
        ram_buffer(73551) := X"3A206261";
        ram_buffer(73552) := X"64206865";
        ram_buffer(73553) := X"61646572";
        ram_buffer(73554) := X"206C656E";
        ram_buffer(73555) := X"67746800";
        ram_buffer(73556) := X"496E7661";
        ram_buffer(73557) := X"6C696420";
        ram_buffer(73558) := X"424D5020";
        ram_buffer(73559) := X"66696C65";
        ram_buffer(73560) := X"3A206269";
        ram_buffer(73561) := X"506C616E";
        ram_buffer(73562) := X"6573206E";
        ram_buffer(73563) := X"6F742065";
        ram_buffer(73564) := X"7175616C";
        ram_buffer(73565) := X"20746F20";
        ram_buffer(73566) := X"31000000";
        ram_buffer(73567) := X"424D5020";
        ram_buffer(73568) := X"6F757470";
        ram_buffer(73569) := X"7574206D";
        ram_buffer(73570) := X"75737420";
        ram_buffer(73571) := X"62652067";
        ram_buffer(73572) := X"72617973";
        ram_buffer(73573) := X"63616C65";
        ram_buffer(73574) := X"206F7220";
        ram_buffer(73575) := X"52474200";
        ram_buffer(73576) := X"536F7272";
        ram_buffer(73577) := X"792C2063";
        ram_buffer(73578) := X"6F6D7072";
        ram_buffer(73579) := X"65737365";
        ram_buffer(73580) := X"6420424D";
        ram_buffer(73581) := X"5073206E";
        ram_buffer(73582) := X"6F742079";
        ram_buffer(73583) := X"65742073";
        ram_buffer(73584) := X"7570706F";
        ram_buffer(73585) := X"72746564";
        ram_buffer(73586) := X"00000000";
        ram_buffer(73587) := X"4E6F7420";
        ram_buffer(73588) := X"6120424D";
        ram_buffer(73589) := X"50206669";
        ram_buffer(73590) := X"6C65202D";
        ram_buffer(73591) := X"20646F65";
        ram_buffer(73592) := X"73206E6F";
        ram_buffer(73593) := X"74207374";
        ram_buffer(73594) := X"61727420";
        ram_buffer(73595) := X"77697468";
        ram_buffer(73596) := X"20424D00";
        ram_buffer(73597) := X"25757825";
        ram_buffer(73598) := X"75203234";
        ram_buffer(73599) := X"2D626974";
        ram_buffer(73600) := X"20424D50";
        ram_buffer(73601) := X"20696D61";
        ram_buffer(73602) := X"67650000";
        ram_buffer(73603) := X"25757825";
        ram_buffer(73604) := X"7520382D";
        ram_buffer(73605) := X"62697420";
        ram_buffer(73606) := X"636F6C6F";
        ram_buffer(73607) := X"726D6170";
        ram_buffer(73608) := X"70656420";
        ram_buffer(73609) := X"424D5020";
        ram_buffer(73610) := X"696D6167";
        ram_buffer(73611) := X"65000000";
        ram_buffer(73612) := X"25757825";
        ram_buffer(73613) := X"75203234";
        ram_buffer(73614) := X"2D626974";
        ram_buffer(73615) := X"204F5332";
        ram_buffer(73616) := X"20424D50";
        ram_buffer(73617) := X"20696D61";
        ram_buffer(73618) := X"67650000";
        ram_buffer(73619) := X"25757825";
        ram_buffer(73620) := X"7520382D";
        ram_buffer(73621) := X"62697420";
        ram_buffer(73622) := X"636F6C6F";
        ram_buffer(73623) := X"726D6170";
        ram_buffer(73624) := X"70656420";
        ram_buffer(73625) := X"4F533220";
        ram_buffer(73626) := X"424D5020";
        ram_buffer(73627) := X"696D6167";
        ram_buffer(73628) := X"65000000";
        ram_buffer(73629) := X"47494620";
        ram_buffer(73630) := X"6F757470";
        ram_buffer(73631) := X"75742067";
        ram_buffer(73632) := X"6F742063";
        ram_buffer(73633) := X"6F6E6675";
        ram_buffer(73634) := X"73656400";
        ram_buffer(73635) := X"426F6775";
        ram_buffer(73636) := X"73204749";
        ram_buffer(73637) := X"4620636F";
        ram_buffer(73638) := X"64657369";
        ram_buffer(73639) := X"7A652025";
        ram_buffer(73640) := X"64000000";
        ram_buffer(73641) := X"47494620";
        ram_buffer(73642) := X"6F757470";
        ram_buffer(73643) := X"7574206D";
        ram_buffer(73644) := X"75737420";
        ram_buffer(73645) := X"62652067";
        ram_buffer(73646) := X"72617973";
        ram_buffer(73647) := X"63616C65";
        ram_buffer(73648) := X"206F7220";
        ram_buffer(73649) := X"52474200";
        ram_buffer(73650) := X"546F6F20";
        ram_buffer(73651) := X"66657720";
        ram_buffer(73652) := X"696D6167";
        ram_buffer(73653) := X"65732069";
        ram_buffer(73654) := X"6E204749";
        ram_buffer(73655) := X"46206669";
        ram_buffer(73656) := X"6C650000";
        ram_buffer(73657) := X"4E6F7420";
        ram_buffer(73658) := X"61204749";
        ram_buffer(73659) := X"46206669";
        ram_buffer(73660) := X"6C650000";
        ram_buffer(73661) := X"25757825";
        ram_buffer(73662) := X"75782564";
        ram_buffer(73663) := X"20474946";
        ram_buffer(73664) := X"20696D61";
        ram_buffer(73665) := X"67650000";
        ram_buffer(73666) := X"5761726E";
        ram_buffer(73667) := X"696E673A";
        ram_buffer(73668) := X"20756E65";
        ram_buffer(73669) := X"78706563";
        ram_buffer(73670) := X"74656420";
        ram_buffer(73671) := X"47494620";
        ram_buffer(73672) := X"76657273";
        ram_buffer(73673) := X"696F6E20";
        ram_buffer(73674) := X"6E756D62";
        ram_buffer(73675) := X"65722027";
        ram_buffer(73676) := X"25632563";
        ram_buffer(73677) := X"25632700";
        ram_buffer(73678) := X"49676E6F";
        ram_buffer(73679) := X"72696E67";
        ram_buffer(73680) := X"20474946";
        ram_buffer(73681) := X"20657874";
        ram_buffer(73682) := X"656E7369";
        ram_buffer(73683) := X"6F6E2062";
        ram_buffer(73684) := X"6C6F636B";
        ram_buffer(73685) := X"206F6620";
        ram_buffer(73686) := X"74797065";
        ram_buffer(73687) := X"20307825";
        ram_buffer(73688) := X"30327800";
        ram_buffer(73689) := X"43617574";
        ram_buffer(73690) := X"696F6E3A";
        ram_buffer(73691) := X"206E6F6E";
        ram_buffer(73692) := X"73717561";
        ram_buffer(73693) := X"72652070";
        ram_buffer(73694) := X"6978656C";
        ram_buffer(73695) := X"7320696E";
        ram_buffer(73696) := X"20696E70";
        ram_buffer(73697) := X"75740000";
        ram_buffer(73698) := X"436F7272";
        ram_buffer(73699) := X"75707420";
        ram_buffer(73700) := X"64617461";
        ram_buffer(73701) := X"20696E20";
        ram_buffer(73702) := X"47494620";
        ram_buffer(73703) := X"66696C65";
        ram_buffer(73704) := X"00000000";
        ram_buffer(73705) := X"426F6775";
        ram_buffer(73706) := X"73206368";
        ram_buffer(73707) := X"61722030";
        ram_buffer(73708) := X"78253032";
        ram_buffer(73709) := X"7820696E";
        ram_buffer(73710) := X"20474946";
        ram_buffer(73711) := X"2066696C";
        ram_buffer(73712) := X"652C2069";
        ram_buffer(73713) := X"676E6F72";
        ram_buffer(73714) := X"696E6700";
        ram_buffer(73715) := X"5072656D";
        ram_buffer(73716) := X"61747572";
        ram_buffer(73717) := X"6520656E";
        ram_buffer(73718) := X"64206F66";
        ram_buffer(73719) := X"20474946";
        ram_buffer(73720) := X"20696D61";
        ram_buffer(73721) := X"67650000";
        ram_buffer(73722) := X"52616E20";
        ram_buffer(73723) := X"6F757420";
        ram_buffer(73724) := X"6F662047";
        ram_buffer(73725) := X"49462062";
        ram_buffer(73726) := X"69747300";
        ram_buffer(73727) := X"50504D20";
        ram_buffer(73728) := X"6F757470";
        ram_buffer(73729) := X"7574206D";
        ram_buffer(73730) := X"75737420";
        ram_buffer(73731) := X"62652067";
        ram_buffer(73732) := X"72617973";
        ram_buffer(73733) := X"63616C65";
        ram_buffer(73734) := X"206F7220";
        ram_buffer(73735) := X"52474200";
        ram_buffer(73736) := X"4E6F6E6E";
        ram_buffer(73737) := X"756D6572";
        ram_buffer(73738) := X"69632064";
        ram_buffer(73739) := X"61746120";
        ram_buffer(73740) := X"696E2050";
        ram_buffer(73741) := X"504D2066";
        ram_buffer(73742) := X"696C6500";
        ram_buffer(73743) := X"4E6F7420";
        ram_buffer(73744) := X"61205050";
        ram_buffer(73745) := X"4D206669";
        ram_buffer(73746) := X"6C650000";
        ram_buffer(73747) := X"25757825";
        ram_buffer(73748) := X"75205047";
        ram_buffer(73749) := X"4D20696D";
        ram_buffer(73750) := X"61676500";
        ram_buffer(73751) := X"25757825";
        ram_buffer(73752) := X"75207465";
        ram_buffer(73753) := X"78742050";
        ram_buffer(73754) := X"474D2069";
        ram_buffer(73755) := X"6D616765";
        ram_buffer(73756) := X"00000000";
        ram_buffer(73757) := X"25757825";
        ram_buffer(73758) := X"75205050";
        ram_buffer(73759) := X"4D20696D";
        ram_buffer(73760) := X"61676500";
        ram_buffer(73761) := X"25757825";
        ram_buffer(73762) := X"75207465";
        ram_buffer(73763) := X"78742050";
        ram_buffer(73764) := X"504D2069";
        ram_buffer(73765) := X"6D616765";
        ram_buffer(73766) := X"00000000";
        ram_buffer(73767) := X"556E7375";
        ram_buffer(73768) := X"70706F72";
        ram_buffer(73769) := X"74656420";
        ram_buffer(73770) := X"54617267";
        ram_buffer(73771) := X"6120636F";
        ram_buffer(73772) := X"6C6F726D";
        ram_buffer(73773) := X"61702066";
        ram_buffer(73774) := X"6F726D61";
        ram_buffer(73775) := X"74000000";
        ram_buffer(73776) := X"496E7661";
        ram_buffer(73777) := X"6C696420";
        ram_buffer(73778) := X"6F722075";
        ram_buffer(73779) := X"6E737570";
        ram_buffer(73780) := X"706F7274";
        ram_buffer(73781) := X"65642054";
        ram_buffer(73782) := X"61726761";
        ram_buffer(73783) := X"2066696C";
        ram_buffer(73784) := X"65000000";
        ram_buffer(73785) := X"54617267";
        ram_buffer(73786) := X"61206F75";
        ram_buffer(73787) := X"74707574";
        ram_buffer(73788) := X"206D7573";
        ram_buffer(73789) := X"74206265";
        ram_buffer(73790) := X"20677261";
        ram_buffer(73791) := X"79736361";
        ram_buffer(73792) := X"6C65206F";
        ram_buffer(73793) := X"72205247";
        ram_buffer(73794) := X"42000000";
        ram_buffer(73795) := X"25757825";
        ram_buffer(73796) := X"75205247";
        ram_buffer(73797) := X"42205461";
        ram_buffer(73798) := X"72676120";
        ram_buffer(73799) := X"696D6167";
        ram_buffer(73800) := X"65000000";
        ram_buffer(73801) := X"25757825";
        ram_buffer(73802) := X"75206772";
        ram_buffer(73803) := X"61797363";
        ram_buffer(73804) := X"616C6520";
        ram_buffer(73805) := X"54617267";
        ram_buffer(73806) := X"6120696D";
        ram_buffer(73807) := X"61676500";
        ram_buffer(73808) := X"25757825";
        ram_buffer(73809) := X"7520636F";
        ram_buffer(73810) := X"6C6F726D";
        ram_buffer(73811) := X"61707065";
        ram_buffer(73812) := X"64205461";
        ram_buffer(73813) := X"72676120";
        ram_buffer(73814) := X"696D6167";
        ram_buffer(73815) := X"65000000";
        ram_buffer(73816) := X"436F6C6F";
        ram_buffer(73817) := X"72206D61";
        ram_buffer(73818) := X"70206669";
        ram_buffer(73819) := X"6C652069";
        ram_buffer(73820) := X"7320696E";
        ram_buffer(73821) := X"76616C69";
        ram_buffer(73822) := X"64206F72";
        ram_buffer(73823) := X"206F6620";
        ram_buffer(73824) := X"756E7375";
        ram_buffer(73825) := X"70706F72";
        ram_buffer(73826) := X"74656420";
        ram_buffer(73827) := X"666F726D";
        ram_buffer(73828) := X"61740000";
        ram_buffer(73829) := X"4F757470";
        ram_buffer(73830) := X"75742066";
        ram_buffer(73831) := X"696C6520";
        ram_buffer(73832) := X"666F726D";
        ram_buffer(73833) := X"61742063";
        ram_buffer(73834) := X"616E6E6F";
        ram_buffer(73835) := X"74206861";
        ram_buffer(73836) := X"6E646C65";
        ram_buffer(73837) := X"20256420";
        ram_buffer(73838) := X"636F6C6F";
        ram_buffer(73839) := X"726D6170";
        ram_buffer(73840) := X"20656E74";
        ram_buffer(73841) := X"72696573";
        ram_buffer(73842) := X"00000000";
        ram_buffer(73843) := X"756E6765";
        ram_buffer(73844) := X"74632066";
        ram_buffer(73845) := X"61696C65";
        ram_buffer(73846) := X"64000000";
        ram_buffer(73847) := X"556E7265";
        ram_buffer(73848) := X"636F676E";
        ram_buffer(73849) := X"697A6564";
        ram_buffer(73850) := X"20696E70";
        ram_buffer(73851) := X"75742066";
        ram_buffer(73852) := X"696C6520";
        ram_buffer(73853) := X"666F726D";
        ram_buffer(73854) := X"6174202D";
        ram_buffer(73855) := X"2D2D2070";
        ram_buffer(73856) := X"65726861";
        ram_buffer(73857) := X"70732079";
        ram_buffer(73858) := X"6F75206E";
        ram_buffer(73859) := X"65656420";
        ram_buffer(73860) := X"2D746172";
        ram_buffer(73861) := X"67610000";
        ram_buffer(73862) := X"556E7375";
        ram_buffer(73863) := X"70706F72";
        ram_buffer(73864) := X"74656420";
        ram_buffer(73865) := X"6F757470";
        ram_buffer(73866) := X"75742066";
        ram_buffer(73867) := X"696C6520";
        ram_buffer(73868) := X"666F726D";
        ram_buffer(73869) := X"61740000";
        ram_buffer(73870) := X"00000000";
        ram_buffer(73871) := X"100C7CE0";
        ram_buffer(73872) := X"100C7D00";
        ram_buffer(73873) := X"100C7D2C";
        ram_buffer(73874) := X"100C7D50";
        ram_buffer(73875) := X"100C7D7C";
        ram_buffer(73876) := X"100C7DA0";
        ram_buffer(73877) := X"100C7DCC";
        ram_buffer(73878) := X"100C7DF4";
        ram_buffer(73879) := X"100C7E0C";
        ram_buffer(73880) := X"100C7E30";
        ram_buffer(73881) := X"100C7E4C";
        ram_buffer(73882) := X"100C7E74";
        ram_buffer(73883) := X"100C7E8C";
        ram_buffer(73884) := X"100C7EA4";
        ram_buffer(73885) := X"100C7EC8";
        ram_buffer(73886) := X"100C7EE4";
        ram_buffer(73887) := X"100C7EF4";
        ram_buffer(73888) := X"100C7F08";
        ram_buffer(73889) := X"100C7F38";
        ram_buffer(73890) := X"100C7F64";
        ram_buffer(73891) := X"100C7F88";
        ram_buffer(73892) := X"100C7FA4";
        ram_buffer(73893) := X"100C7FCC";
        ram_buffer(73894) := X"100C7FE8";
        ram_buffer(73895) := X"100C7FFC";
        ram_buffer(73896) := X"100C8020";
        ram_buffer(73897) := X"100C803C";
        ram_buffer(73898) := X"100C804C";
        ram_buffer(73899) := X"100C805C";
        ram_buffer(73900) := X"100C8074";
        ram_buffer(73901) := X"100C8084";
        ram_buffer(73902) := X"100C809C";
        ram_buffer(73903) := X"100C80C0";
        ram_buffer(73904) := X"100C80E4";
        ram_buffer(73905) := X"100C810C";
        ram_buffer(73906) := X"100C8124";
        ram_buffer(73907) := X"100C8140";
        ram_buffer(73908) := X"100C8160";
        ram_buffer(73909) := X"100C8194";
        ram_buffer(73910) := X"100C81CC";
        ram_buffer(73911) := X"100C81DC";
        ram_buffer(73912) := X"100C8218";
        ram_buffer(73913) := X"00000000";
        ram_buffer(73914) := X"00081019";
        ram_buffer(73915) := X"2129313A";
        ram_buffer(73916) := X"424A525A";
        ram_buffer(73917) := X"636B737B";
        ram_buffer(73918) := X"848C949C";
        ram_buffer(73919) := X"A5ADB5BD";
        ram_buffer(73920) := X"C5CED6DE";
        ram_buffer(73921) := X"E6EFF7FF";
        ram_buffer(73922) := X"43616E27";
        ram_buffer(73923) := X"74206F70";
        ram_buffer(73924) := X"656E2074";
        ram_buffer(73925) := X"61626C65";
        ram_buffer(73926) := X"2066696C";
        ram_buffer(73927) := X"65202573";
        ram_buffer(73928) := X"0A000000";
        ram_buffer(73929) := X"546F6F20";
        ram_buffer(73930) := X"6D616E79";
        ram_buffer(73931) := X"20746162";
        ram_buffer(73932) := X"6C657320";
        ram_buffer(73933) := X"696E2066";
        ram_buffer(73934) := X"696C6520";
        ram_buffer(73935) := X"25730A00";
        ram_buffer(73936) := X"496E7661";
        ram_buffer(73937) := X"6C696420";
        ram_buffer(73938) := X"7461626C";
        ram_buffer(73939) := X"65206461";
        ram_buffer(73940) := X"74612069";
        ram_buffer(73941) := X"6E206669";
        ram_buffer(73942) := X"6C652025";
        ram_buffer(73943) := X"730A0000";
        ram_buffer(73944) := X"4E6F6E2D";
        ram_buffer(73945) := X"6E756D65";
        ram_buffer(73946) := X"72696320";
        ram_buffer(73947) := X"64617461";
        ram_buffer(73948) := X"20696E20";
        ram_buffer(73949) := X"66696C65";
        ram_buffer(73950) := X"2025730A";
        ram_buffer(73951) := X"00000000";
        ram_buffer(73952) := X"43616E27";
        ram_buffer(73953) := X"74206F70";
        ram_buffer(73954) := X"656E2073";
        ram_buffer(73955) := X"63616E20";
        ram_buffer(73956) := X"64656669";
        ram_buffer(73957) := X"6E697469";
        ram_buffer(73958) := X"6F6E2066";
        ram_buffer(73959) := X"696C6520";
        ram_buffer(73960) := X"25730A00";
        ram_buffer(73961) := X"546F6F20";
        ram_buffer(73962) := X"6D616E79";
        ram_buffer(73963) := X"20736361";
        ram_buffer(73964) := X"6E732064";
        ram_buffer(73965) := X"6566696E";
        ram_buffer(73966) := X"65642069";
        ram_buffer(73967) := X"6E206669";
        ram_buffer(73968) := X"6C652025";
        ram_buffer(73969) := X"730A0000";
        ram_buffer(73970) := X"546F6F20";
        ram_buffer(73971) := X"6D616E79";
        ram_buffer(73972) := X"20636F6D";
        ram_buffer(73973) := X"706F6E65";
        ram_buffer(73974) := X"6E747320";
        ram_buffer(73975) := X"696E206F";
        ram_buffer(73976) := X"6E652073";
        ram_buffer(73977) := X"63616E20";
        ram_buffer(73978) := X"696E2066";
        ram_buffer(73979) := X"696C6520";
        ram_buffer(73980) := X"25730A00";
        ram_buffer(73981) := X"496E7661";
        ram_buffer(73982) := X"6C696420";
        ram_buffer(73983) := X"7363616E";
        ram_buffer(73984) := X"20656E74";
        ram_buffer(73985) := X"72792066";
        ram_buffer(73986) := X"6F726D61";
        ram_buffer(73987) := X"7420696E";
        ram_buffer(73988) := X"2066696C";
        ram_buffer(73989) := X"65202573";
        ram_buffer(73990) := X"0A000000";
        ram_buffer(73991) := X"4A504547";
        ram_buffer(73992) := X"20717561";
        ram_buffer(73993) := X"6E74697A";
        ram_buffer(73994) := X"6174696F";
        ram_buffer(73995) := X"6E207461";
        ram_buffer(73996) := X"626C6573";
        ram_buffer(73997) := X"20617265";
        ram_buffer(73998) := X"206E756D";
        ram_buffer(73999) := X"62657265";
        ram_buffer(74000) := X"6420302E";
        ram_buffer(74001) := X"2E25640A";
        ram_buffer(74002) := X"00000000";
        ram_buffer(74003) := X"25642563";
        ram_buffer(74004) := X"25642563";
        ram_buffer(74005) := X"00000000";
        ram_buffer(74006) := X"4A504547";
        ram_buffer(74007) := X"2073616D";
        ram_buffer(74008) := X"706C696E";
        ram_buffer(74009) := X"67206661";
        ram_buffer(74010) := X"63746F72";
        ram_buffer(74011) := X"73206D75";
        ram_buffer(74012) := X"73742062";
        ram_buffer(74013) := X"6520312E";
        ram_buffer(74014) := X"2E340A00";
        ram_buffer(74015) := X"100877B0";
        ram_buffer(74016) := X"10087844";
        ram_buffer(74017) := X"10087638";
        ram_buffer(74018) := X"10087638";
        ram_buffer(74019) := X"100878B8";
        ram_buffer(74020) := X"100876E4";
        ram_buffer(74021) := X"10087B98";
        ram_buffer(74022) := X"10087BF4";
        ram_buffer(74023) := X"10087C30";
        ram_buffer(74024) := X"10087CAC";
        ram_buffer(74025) := X"10087A70";
        ram_buffer(74026) := X"10087B08";
        ram_buffer(74027) := X"10088290";
        ram_buffer(74028) := X"10088204";
        ram_buffer(74029) := X"10088158";
        ram_buffer(74030) := X"10088158";
        ram_buffer(74031) := X"100882A8";
        ram_buffer(74032) := X"10088278";
        ram_buffer(74033) := X"00010203";
        ram_buffer(74034) := X"11040521";
        ram_buffer(74035) := X"31061241";
        ram_buffer(74036) := X"51076171";
        ram_buffer(74037) := X"13223281";
        ram_buffer(74038) := X"08144291";
        ram_buffer(74039) := X"A1B1C109";
        ram_buffer(74040) := X"233352F0";
        ram_buffer(74041) := X"156272D1";
        ram_buffer(74042) := X"0A162434";
        ram_buffer(74043) := X"E125F117";
        ram_buffer(74044) := X"18191A26";
        ram_buffer(74045) := X"2728292A";
        ram_buffer(74046) := X"35363738";
        ram_buffer(74047) := X"393A4344";
        ram_buffer(74048) := X"45464748";
        ram_buffer(74049) := X"494A5354";
        ram_buffer(74050) := X"55565758";
        ram_buffer(74051) := X"595A6364";
        ram_buffer(74052) := X"65666768";
        ram_buffer(74053) := X"696A7374";
        ram_buffer(74054) := X"75767778";
        ram_buffer(74055) := X"797A8283";
        ram_buffer(74056) := X"84858687";
        ram_buffer(74057) := X"88898A92";
        ram_buffer(74058) := X"93949596";
        ram_buffer(74059) := X"9798999A";
        ram_buffer(74060) := X"A2A3A4A5";
        ram_buffer(74061) := X"A6A7A8A9";
        ram_buffer(74062) := X"AAB2B3B4";
        ram_buffer(74063) := X"B5B6B7B8";
        ram_buffer(74064) := X"B9BAC2C3";
        ram_buffer(74065) := X"C4C5C6C7";
        ram_buffer(74066) := X"C8C9CAD2";
        ram_buffer(74067) := X"D3D4D5D6";
        ram_buffer(74068) := X"D7D8D9DA";
        ram_buffer(74069) := X"E2E3E4E5";
        ram_buffer(74070) := X"E6E7E8E9";
        ram_buffer(74071) := X"EAF2F3F4";
        ram_buffer(74072) := X"F5F6F7F8";
        ram_buffer(74073) := X"F9FA0000";
        ram_buffer(74074) := X"00000201";
        ram_buffer(74075) := X"02040403";
        ram_buffer(74076) := X"04070504";
        ram_buffer(74077) := X"04000102";
        ram_buffer(74078) := X"77000000";
        ram_buffer(74079) := X"00010203";
        ram_buffer(74080) := X"04050607";
        ram_buffer(74081) := X"08090A0B";
        ram_buffer(74082) := X"00000301";
        ram_buffer(74083) := X"01010101";
        ram_buffer(74084) := X"01010101";
        ram_buffer(74085) := X"00000000";
        ram_buffer(74086) := X"00000000";
        ram_buffer(74087) := X"01020300";
        ram_buffer(74088) := X"04110512";
        ram_buffer(74089) := X"21314106";
        ram_buffer(74090) := X"13516107";
        ram_buffer(74091) := X"22711432";
        ram_buffer(74092) := X"8191A108";
        ram_buffer(74093) := X"2342B1C1";
        ram_buffer(74094) := X"1552D1F0";
        ram_buffer(74095) := X"24336272";
        ram_buffer(74096) := X"82090A16";
        ram_buffer(74097) := X"1718191A";
        ram_buffer(74098) := X"25262728";
        ram_buffer(74099) := X"292A3435";
        ram_buffer(74100) := X"36373839";
        ram_buffer(74101) := X"3A434445";
        ram_buffer(74102) := X"46474849";
        ram_buffer(74103) := X"4A535455";
        ram_buffer(74104) := X"56575859";
        ram_buffer(74105) := X"5A636465";
        ram_buffer(74106) := X"66676869";
        ram_buffer(74107) := X"6A737475";
        ram_buffer(74108) := X"76777879";
        ram_buffer(74109) := X"7A838485";
        ram_buffer(74110) := X"86878889";
        ram_buffer(74111) := X"8A929394";
        ram_buffer(74112) := X"95969798";
        ram_buffer(74113) := X"999AA2A3";
        ram_buffer(74114) := X"A4A5A6A7";
        ram_buffer(74115) := X"A8A9AAB2";
        ram_buffer(74116) := X"B3B4B5B6";
        ram_buffer(74117) := X"B7B8B9BA";
        ram_buffer(74118) := X"C2C3C4C5";
        ram_buffer(74119) := X"C6C7C8C9";
        ram_buffer(74120) := X"CAD2D3D4";
        ram_buffer(74121) := X"D5D6D7D8";
        ram_buffer(74122) := X"D9DAE1E2";
        ram_buffer(74123) := X"E3E4E5E6";
        ram_buffer(74124) := X"E7E8E9EA";
        ram_buffer(74125) := X"F1F2F3F4";
        ram_buffer(74126) := X"F5F6F7F8";
        ram_buffer(74127) := X"F9FA0000";
        ram_buffer(74128) := X"00000201";
        ram_buffer(74129) := X"03030204";
        ram_buffer(74130) := X"03050504";
        ram_buffer(74131) := X"04000001";
        ram_buffer(74132) := X"7D000000";
        ram_buffer(74133) := X"00010203";
        ram_buffer(74134) := X"04050607";
        ram_buffer(74135) := X"08090A0B";
        ram_buffer(74136) := X"00000105";
        ram_buffer(74137) := X"01010101";
        ram_buffer(74138) := X"01010000";
        ram_buffer(74139) := X"00000000";
        ram_buffer(74140) := X"00000000";
        ram_buffer(74141) := X"00000011";
        ram_buffer(74142) := X"00000012";
        ram_buffer(74143) := X"00000018";
        ram_buffer(74144) := X"0000002F";
        ram_buffer(74145) := X"00000063";
        ram_buffer(74146) := X"00000063";
        ram_buffer(74147) := X"00000063";
        ram_buffer(74148) := X"00000063";
        ram_buffer(74149) := X"00000012";
        ram_buffer(74150) := X"00000015";
        ram_buffer(74151) := X"0000001A";
        ram_buffer(74152) := X"00000042";
        ram_buffer(74153) := X"00000063";
        ram_buffer(74154) := X"00000063";
        ram_buffer(74155) := X"00000063";
        ram_buffer(74156) := X"00000063";
        ram_buffer(74157) := X"00000018";
        ram_buffer(74158) := X"0000001A";
        ram_buffer(74159) := X"00000038";
        ram_buffer(74160) := X"00000063";
        ram_buffer(74161) := X"00000063";
        ram_buffer(74162) := X"00000063";
        ram_buffer(74163) := X"00000063";
        ram_buffer(74164) := X"00000063";
        ram_buffer(74165) := X"0000002F";
        ram_buffer(74166) := X"00000042";
        ram_buffer(74167) := X"00000063";
        ram_buffer(74168) := X"00000063";
        ram_buffer(74169) := X"00000063";
        ram_buffer(74170) := X"00000063";
        ram_buffer(74171) := X"00000063";
        ram_buffer(74172) := X"00000063";
        ram_buffer(74173) := X"00000063";
        ram_buffer(74174) := X"00000063";
        ram_buffer(74175) := X"00000063";
        ram_buffer(74176) := X"00000063";
        ram_buffer(74177) := X"00000063";
        ram_buffer(74178) := X"00000063";
        ram_buffer(74179) := X"00000063";
        ram_buffer(74180) := X"00000063";
        ram_buffer(74181) := X"00000063";
        ram_buffer(74182) := X"00000063";
        ram_buffer(74183) := X"00000063";
        ram_buffer(74184) := X"00000063";
        ram_buffer(74185) := X"00000063";
        ram_buffer(74186) := X"00000063";
        ram_buffer(74187) := X"00000063";
        ram_buffer(74188) := X"00000063";
        ram_buffer(74189) := X"00000063";
        ram_buffer(74190) := X"00000063";
        ram_buffer(74191) := X"00000063";
        ram_buffer(74192) := X"00000063";
        ram_buffer(74193) := X"00000063";
        ram_buffer(74194) := X"00000063";
        ram_buffer(74195) := X"00000063";
        ram_buffer(74196) := X"00000063";
        ram_buffer(74197) := X"00000063";
        ram_buffer(74198) := X"00000063";
        ram_buffer(74199) := X"00000063";
        ram_buffer(74200) := X"00000063";
        ram_buffer(74201) := X"00000063";
        ram_buffer(74202) := X"00000063";
        ram_buffer(74203) := X"00000063";
        ram_buffer(74204) := X"00000063";
        ram_buffer(74205) := X"00000010";
        ram_buffer(74206) := X"0000000B";
        ram_buffer(74207) := X"0000000A";
        ram_buffer(74208) := X"00000010";
        ram_buffer(74209) := X"00000018";
        ram_buffer(74210) := X"00000028";
        ram_buffer(74211) := X"00000033";
        ram_buffer(74212) := X"0000003D";
        ram_buffer(74213) := X"0000000C";
        ram_buffer(74214) := X"0000000C";
        ram_buffer(74215) := X"0000000E";
        ram_buffer(74216) := X"00000013";
        ram_buffer(74217) := X"0000001A";
        ram_buffer(74218) := X"0000003A";
        ram_buffer(74219) := X"0000003C";
        ram_buffer(74220) := X"00000037";
        ram_buffer(74221) := X"0000000E";
        ram_buffer(74222) := X"0000000D";
        ram_buffer(74223) := X"00000010";
        ram_buffer(74224) := X"00000018";
        ram_buffer(74225) := X"00000028";
        ram_buffer(74226) := X"00000039";
        ram_buffer(74227) := X"00000045";
        ram_buffer(74228) := X"00000038";
        ram_buffer(74229) := X"0000000E";
        ram_buffer(74230) := X"00000011";
        ram_buffer(74231) := X"00000016";
        ram_buffer(74232) := X"0000001D";
        ram_buffer(74233) := X"00000033";
        ram_buffer(74234) := X"00000057";
        ram_buffer(74235) := X"00000050";
        ram_buffer(74236) := X"0000003E";
        ram_buffer(74237) := X"00000012";
        ram_buffer(74238) := X"00000016";
        ram_buffer(74239) := X"00000025";
        ram_buffer(74240) := X"00000038";
        ram_buffer(74241) := X"00000044";
        ram_buffer(74242) := X"0000006D";
        ram_buffer(74243) := X"00000067";
        ram_buffer(74244) := X"0000004D";
        ram_buffer(74245) := X"00000018";
        ram_buffer(74246) := X"00000023";
        ram_buffer(74247) := X"00000037";
        ram_buffer(74248) := X"00000040";
        ram_buffer(74249) := X"00000051";
        ram_buffer(74250) := X"00000068";
        ram_buffer(74251) := X"00000071";
        ram_buffer(74252) := X"0000005C";
        ram_buffer(74253) := X"00000031";
        ram_buffer(74254) := X"00000040";
        ram_buffer(74255) := X"0000004E";
        ram_buffer(74256) := X"00000057";
        ram_buffer(74257) := X"00000067";
        ram_buffer(74258) := X"00000079";
        ram_buffer(74259) := X"00000078";
        ram_buffer(74260) := X"00000065";
        ram_buffer(74261) := X"00000048";
        ram_buffer(74262) := X"0000005C";
        ram_buffer(74263) := X"0000005F";
        ram_buffer(74264) := X"00000062";
        ram_buffer(74265) := X"00000070";
        ram_buffer(74266) := X"00000064";
        ram_buffer(74267) := X"00000067";
        ram_buffer(74268) := X"00000063";
        ram_buffer(74269) := X"1008FED8";
        ram_buffer(74270) := X"1008FEC0";
        ram_buffer(74271) := X"1008FEA8";
        ram_buffer(74272) := X"1008FEA8";
        ram_buffer(74273) := X"1008FE50";
        ram_buffer(74274) := X"1008FE50";
        ram_buffer(74275) := X"10090090";
        ram_buffer(74276) := X"10090038";
        ram_buffer(74277) := X"1008FFF8";
        ram_buffer(74278) := X"1008FFB0";
        ram_buffer(74279) := X"1008FF58";
        ram_buffer(74280) := X"1008FEF0";
        ram_buffer(74281) := X"00000000";
        ram_buffer(74282) := X"3FF00000";
        ram_buffer(74283) := X"00000000";
        ram_buffer(74284) := X"3FF63150";
        ram_buffer(74285) := X"B14861EF";
        ram_buffer(74286) := X"3FF4E7AE";
        ram_buffer(74287) := X"914D6FCA";
        ram_buffer(74288) := X"3FF2D062";
        ram_buffer(74289) := X"EF6C11AA";
        ram_buffer(74290) := X"3FF00000";
        ram_buffer(74291) := X"00000000";
        ram_buffer(74292) := X"3FE92469";
        ram_buffer(74293) := X"C0A7BF3B";
        ram_buffer(74294) := X"3FE1517A";
        ram_buffer(74295) := X"7BC720BB";
        ram_buffer(74296) := X"3FD1A855";
        ram_buffer(74297) := X"DE72AB5D";
        ram_buffer(74298) := X"400058C5";
        ram_buffer(74299) := X"539F4B42";
        ram_buffer(74300) := X"40003249";
        ram_buffer(74301) := X"22A311A8";
        ram_buffer(74302) := X"58C57B21";
        ram_buffer(74303) := X"73FC6862";
        ram_buffer(74304) := X"58C545BF";
        ram_buffer(74305) := X"300B187E";
        ram_buffer(74306) := X"539F73FC";
        ram_buffer(74307) := X"6D416254";
        ram_buffer(74308) := X"539F41B3";
        ram_buffer(74309) := X"2D411712";
        ram_buffer(74310) := X"4B426862";
        ram_buffer(74311) := X"6254587E";
        ram_buffer(74312) := X"4B423B21";
        ram_buffer(74313) := X"28BA14C3";
        ram_buffer(74314) := X"400058C5";
        ram_buffer(74315) := X"539F4B42";
        ram_buffer(74316) := X"40003249";
        ram_buffer(74317) := X"22A311A8";
        ram_buffer(74318) := X"324945BF";
        ram_buffer(74319) := X"41B33B21";
        ram_buffer(74320) := X"32492782";
        ram_buffer(74321) := X"1B370DE0";
        ram_buffer(74322) := X"22A3300B";
        ram_buffer(74323) := X"2D4128BA";
        ram_buffer(74324) := X"22A31B37";
        ram_buffer(74325) := X"12BF098E";
        ram_buffer(74326) := X"11A8187E";
        ram_buffer(74327) := X"171214C3";
        ram_buffer(74328) := X"11A80DE0";
        ram_buffer(74329) := X"098E04DF";
        ram_buffer(74330) := X"00000000";
        ram_buffer(74331) := X"00000001";
        ram_buffer(74332) := X"00000008";
        ram_buffer(74333) := X"00000010";
        ram_buffer(74334) := X"00000009";
        ram_buffer(74335) := X"00000002";
        ram_buffer(74336) := X"00000003";
        ram_buffer(74337) := X"0000000A";
        ram_buffer(74338) := X"00000011";
        ram_buffer(74339) := X"00000018";
        ram_buffer(74340) := X"00000020";
        ram_buffer(74341) := X"00000019";
        ram_buffer(74342) := X"00000012";
        ram_buffer(74343) := X"0000000B";
        ram_buffer(74344) := X"00000004";
        ram_buffer(74345) := X"00000005";
        ram_buffer(74346) := X"0000000C";
        ram_buffer(74347) := X"00000013";
        ram_buffer(74348) := X"0000001A";
        ram_buffer(74349) := X"00000021";
        ram_buffer(74350) := X"00000028";
        ram_buffer(74351) := X"00000030";
        ram_buffer(74352) := X"00000029";
        ram_buffer(74353) := X"00000022";
        ram_buffer(74354) := X"0000001B";
        ram_buffer(74355) := X"00000014";
        ram_buffer(74356) := X"0000000D";
        ram_buffer(74357) := X"00000006";
        ram_buffer(74358) := X"00000007";
        ram_buffer(74359) := X"0000000E";
        ram_buffer(74360) := X"00000015";
        ram_buffer(74361) := X"0000001C";
        ram_buffer(74362) := X"00000023";
        ram_buffer(74363) := X"0000002A";
        ram_buffer(74364) := X"00000031";
        ram_buffer(74365) := X"00000038";
        ram_buffer(74366) := X"00000039";
        ram_buffer(74367) := X"00000032";
        ram_buffer(74368) := X"0000002B";
        ram_buffer(74369) := X"00000024";
        ram_buffer(74370) := X"0000001D";
        ram_buffer(74371) := X"00000016";
        ram_buffer(74372) := X"0000000F";
        ram_buffer(74373) := X"00000017";
        ram_buffer(74374) := X"0000001E";
        ram_buffer(74375) := X"00000025";
        ram_buffer(74376) := X"0000002C";
        ram_buffer(74377) := X"00000033";
        ram_buffer(74378) := X"0000003A";
        ram_buffer(74379) := X"0000003B";
        ram_buffer(74380) := X"00000034";
        ram_buffer(74381) := X"0000002D";
        ram_buffer(74382) := X"00000026";
        ram_buffer(74383) := X"0000001F";
        ram_buffer(74384) := X"00000027";
        ram_buffer(74385) := X"0000002E";
        ram_buffer(74386) := X"00000035";
        ram_buffer(74387) := X"0000003C";
        ram_buffer(74388) := X"0000003D";
        ram_buffer(74389) := X"00000036";
        ram_buffer(74390) := X"0000002F";
        ram_buffer(74391) := X"00000037";
        ram_buffer(74392) := X"0000003E";
        ram_buffer(74393) := X"0000003F";
        ram_buffer(74394) := X"0000003F";
        ram_buffer(74395) := X"0000003F";
        ram_buffer(74396) := X"0000003F";
        ram_buffer(74397) := X"0000003F";
        ram_buffer(74398) := X"0000003F";
        ram_buffer(74399) := X"0000003F";
        ram_buffer(74400) := X"0000003F";
        ram_buffer(74401) := X"0000003F";
        ram_buffer(74402) := X"0000003F";
        ram_buffer(74403) := X"0000003F";
        ram_buffer(74404) := X"0000003F";
        ram_buffer(74405) := X"0000003F";
        ram_buffer(74406) := X"0000003F";
        ram_buffer(74407) := X"0000003F";
        ram_buffer(74408) := X"0000003F";
        ram_buffer(74409) := X"0000003F";
        ram_buffer(74410) := X"426F6775";
        ram_buffer(74411) := X"73206D65";
        ram_buffer(74412) := X"73736167";
        ram_buffer(74413) := X"6520636F";
        ram_buffer(74414) := X"64652025";
        ram_buffer(74415) := X"64000000";
        ram_buffer(74416) := X"536F7272";
        ram_buffer(74417) := X"792C2074";
        ram_buffer(74418) := X"68657265";
        ram_buffer(74419) := X"20617265";
        ram_buffer(74420) := X"206C6567";
        ram_buffer(74421) := X"616C2072";
        ram_buffer(74422) := X"65737472";
        ram_buffer(74423) := X"69637469";
        ram_buffer(74424) := X"6F6E7320";
        ram_buffer(74425) := X"6F6E2061";
        ram_buffer(74426) := X"72697468";
        ram_buffer(74427) := X"6D657469";
        ram_buffer(74428) := X"6320636F";
        ram_buffer(74429) := X"64696E67";
        ram_buffer(74430) := X"00000000";
        ram_buffer(74431) := X"414C4947";
        ram_buffer(74432) := X"4E5F5459";
        ram_buffer(74433) := X"50452069";
        ram_buffer(74434) := X"73207772";
        ram_buffer(74435) := X"6F6E672C";
        ram_buffer(74436) := X"20706C65";
        ram_buffer(74437) := X"61736520";
        ram_buffer(74438) := X"66697800";
        ram_buffer(74439) := X"4D41585F";
        ram_buffer(74440) := X"414C4C4F";
        ram_buffer(74441) := X"435F4348";
        ram_buffer(74442) := X"554E4B20";
        ram_buffer(74443) := X"69732077";
        ram_buffer(74444) := X"726F6E67";
        ram_buffer(74445) := X"2C20706C";
        ram_buffer(74446) := X"65617365";
        ram_buffer(74447) := X"20666978";
        ram_buffer(74448) := X"00000000";
        ram_buffer(74449) := X"426F6775";
        ram_buffer(74450) := X"73206275";
        ram_buffer(74451) := X"66666572";
        ram_buffer(74452) := X"20636F6E";
        ram_buffer(74453) := X"74726F6C";
        ram_buffer(74454) := X"206D6F64";
        ram_buffer(74455) := X"65000000";
        ram_buffer(74456) := X"496E7661";
        ram_buffer(74457) := X"6C696420";
        ram_buffer(74458) := X"636F6D70";
        ram_buffer(74459) := X"6F6E656E";
        ram_buffer(74460) := X"74204944";
        ram_buffer(74461) := X"20256420";
        ram_buffer(74462) := X"696E2053";
        ram_buffer(74463) := X"4F530000";
        ram_buffer(74464) := X"49444354";
        ram_buffer(74465) := X"206F7574";
        ram_buffer(74466) := X"70757420";
        ram_buffer(74467) := X"626C6F63";
        ram_buffer(74468) := X"6B207369";
        ram_buffer(74469) := X"7A652025";
        ram_buffer(74470) := X"64206E6F";
        ram_buffer(74471) := X"74207375";
        ram_buffer(74472) := X"70706F72";
        ram_buffer(74473) := X"74656400";
        ram_buffer(74474) := X"426F6775";
        ram_buffer(74475) := X"7320696E";
        ram_buffer(74476) := X"70757420";
        ram_buffer(74477) := X"636F6C6F";
        ram_buffer(74478) := X"72737061";
        ram_buffer(74479) := X"63650000";
        ram_buffer(74480) := X"426F6775";
        ram_buffer(74481) := X"73204A50";
        ram_buffer(74482) := X"45472063";
        ram_buffer(74483) := X"6F6C6F72";
        ram_buffer(74484) := X"73706163";
        ram_buffer(74485) := X"65000000";
        ram_buffer(74486) := X"426F6775";
        ram_buffer(74487) := X"73206D61";
        ram_buffer(74488) := X"726B6572";
        ram_buffer(74489) := X"206C656E";
        ram_buffer(74490) := X"67746800";
        ram_buffer(74491) := X"57726F6E";
        ram_buffer(74492) := X"67204A50";
        ram_buffer(74493) := X"4547206C";
        ram_buffer(74494) := X"69627261";
        ram_buffer(74495) := X"72792076";
        ram_buffer(74496) := X"65727369";
        ram_buffer(74497) := X"6F6E3A20";
        ram_buffer(74498) := X"6C696272";
        ram_buffer(74499) := X"61727920";
        ram_buffer(74500) := X"69732025";
        ram_buffer(74501) := X"642C2063";
        ram_buffer(74502) := X"616C6C65";
        ram_buffer(74503) := X"72206578";
        ram_buffer(74504) := X"70656374";
        ram_buffer(74505) := X"73202564";
        ram_buffer(74506) := X"00000000";
        ram_buffer(74507) := X"53616D70";
        ram_buffer(74508) := X"6C696E67";
        ram_buffer(74509) := X"20666163";
        ram_buffer(74510) := X"746F7273";
        ram_buffer(74511) := X"20746F6F";
        ram_buffer(74512) := X"206C6172";
        ram_buffer(74513) := X"67652066";
        ram_buffer(74514) := X"6F722069";
        ram_buffer(74515) := X"6E746572";
        ram_buffer(74516) := X"6C656176";
        ram_buffer(74517) := X"65642073";
        ram_buffer(74518) := X"63616E00";
        ram_buffer(74519) := X"496E7661";
        ram_buffer(74520) := X"6C696420";
        ram_buffer(74521) := X"6D656D6F";
        ram_buffer(74522) := X"72792070";
        ram_buffer(74523) := X"6F6F6C20";
        ram_buffer(74524) := X"636F6465";
        ram_buffer(74525) := X"20256400";
        ram_buffer(74526) := X"556E7375";
        ram_buffer(74527) := X"70706F72";
        ram_buffer(74528) := X"74656420";
        ram_buffer(74529) := X"4A504547";
        ram_buffer(74530) := X"20646174";
        ram_buffer(74531) := X"61207072";
        ram_buffer(74532) := X"65636973";
        ram_buffer(74533) := X"696F6E20";
        ram_buffer(74534) := X"25640000";
        ram_buffer(74535) := X"496E7661";
        ram_buffer(74536) := X"6C696420";
        ram_buffer(74537) := X"70726F67";
        ram_buffer(74538) := X"72657373";
        ram_buffer(74539) := X"69766520";
        ram_buffer(74540) := X"70617261";
        ram_buffer(74541) := X"6D657465";
        ram_buffer(74542) := X"72732053";
        ram_buffer(74543) := X"733D2564";
        ram_buffer(74544) := X"2053653D";
        ram_buffer(74545) := X"25642041";
        ram_buffer(74546) := X"683D2564";
        ram_buffer(74547) := X"20416C3D";
        ram_buffer(74548) := X"25640000";
        ram_buffer(74549) := X"496E7661";
        ram_buffer(74550) := X"6C696420";
        ram_buffer(74551) := X"70726F67";
        ram_buffer(74552) := X"72657373";
        ram_buffer(74553) := X"69766520";
        ram_buffer(74554) := X"70617261";
        ram_buffer(74555) := X"6D657465";
        ram_buffer(74556) := X"72732061";
        ram_buffer(74557) := X"74207363";
        ram_buffer(74558) := X"616E2073";
        ram_buffer(74559) := X"63726970";
        ram_buffer(74560) := X"7420656E";
        ram_buffer(74561) := X"74727920";
        ram_buffer(74562) := X"25640000";
        ram_buffer(74563) := X"426F6775";
        ram_buffer(74564) := X"73207361";
        ram_buffer(74565) := X"6D706C69";
        ram_buffer(74566) := X"6E672066";
        ram_buffer(74567) := X"6163746F";
        ram_buffer(74568) := X"72730000";
        ram_buffer(74569) := X"496E7661";
        ram_buffer(74570) := X"6C696420";
        ram_buffer(74571) := X"7363616E";
        ram_buffer(74572) := X"20736372";
        ram_buffer(74573) := X"69707420";
        ram_buffer(74574) := X"61742065";
        ram_buffer(74575) := X"6E747279";
        ram_buffer(74576) := X"20256400";
        ram_buffer(74577) := X"496D7072";
        ram_buffer(74578) := X"6F706572";
        ram_buffer(74579) := X"2063616C";
        ram_buffer(74580) := X"6C20746F";
        ram_buffer(74581) := X"204A5045";
        ram_buffer(74582) := X"47206C69";
        ram_buffer(74583) := X"62726172";
        ram_buffer(74584) := X"7920696E";
        ram_buffer(74585) := X"20737461";
        ram_buffer(74586) := X"74652025";
        ram_buffer(74587) := X"64000000";
        ram_buffer(74588) := X"4A504547";
        ram_buffer(74589) := X"20706172";
        ram_buffer(74590) := X"616D6574";
        ram_buffer(74591) := X"65722073";
        ram_buffer(74592) := X"74727563";
        ram_buffer(74593) := X"74206D69";
        ram_buffer(74594) := X"736D6174";
        ram_buffer(74595) := X"63683A20";
        ram_buffer(74596) := X"6C696272";
        ram_buffer(74597) := X"61727920";
        ram_buffer(74598) := X"7468696E";
        ram_buffer(74599) := X"6B732073";
        ram_buffer(74600) := X"697A6520";
        ram_buffer(74601) := X"69732025";
        ram_buffer(74602) := X"752C2063";
        ram_buffer(74603) := X"616C6C65";
        ram_buffer(74604) := X"72206578";
        ram_buffer(74605) := X"70656374";
        ram_buffer(74606) := X"73202575";
        ram_buffer(74607) := X"00000000";
        ram_buffer(74608) := X"426F6775";
        ram_buffer(74609) := X"73207669";
        ram_buffer(74610) := X"72747561";
        ram_buffer(74611) := X"6C206172";
        ram_buffer(74612) := X"72617920";
        ram_buffer(74613) := X"61636365";
        ram_buffer(74614) := X"73730000";
        ram_buffer(74615) := X"42756666";
        ram_buffer(74616) := X"65722070";
        ram_buffer(74617) := X"61737365";
        ram_buffer(74618) := X"6420746F";
        ram_buffer(74619) := X"204A5045";
        ram_buffer(74620) := X"47206C69";
        ram_buffer(74621) := X"62726172";
        ram_buffer(74622) := X"79206973";
        ram_buffer(74623) := X"20746F6F";
        ram_buffer(74624) := X"20736D61";
        ram_buffer(74625) := X"6C6C0000";
        ram_buffer(74626) := X"53757370";
        ram_buffer(74627) := X"656E7369";
        ram_buffer(74628) := X"6F6E206E";
        ram_buffer(74629) := X"6F742061";
        ram_buffer(74630) := X"6C6C6F77";
        ram_buffer(74631) := X"65642068";
        ram_buffer(74632) := X"65726500";
        ram_buffer(74633) := X"43434952";
        ram_buffer(74634) := X"36303120";
        ram_buffer(74635) := X"73616D70";
        ram_buffer(74636) := X"6C696E67";
        ram_buffer(74637) := X"206E6F74";
        ram_buffer(74638) := X"20696D70";
        ram_buffer(74639) := X"6C656D65";
        ram_buffer(74640) := X"6E746564";
        ram_buffer(74641) := X"20796574";
        ram_buffer(74642) := X"00000000";
        ram_buffer(74643) := X"546F6F20";
        ram_buffer(74644) := X"6D616E79";
        ram_buffer(74645) := X"20636F6C";
        ram_buffer(74646) := X"6F722063";
        ram_buffer(74647) := X"6F6D706F";
        ram_buffer(74648) := X"6E656E74";
        ram_buffer(74649) := X"733A2025";
        ram_buffer(74650) := X"642C206D";
        ram_buffer(74651) := X"61782025";
        ram_buffer(74652) := X"64000000";
        ram_buffer(74653) := X"556E7375";
        ram_buffer(74654) := X"70706F72";
        ram_buffer(74655) := X"74656420";
        ram_buffer(74656) := X"636F6C6F";
        ram_buffer(74657) := X"7220636F";
        ram_buffer(74658) := X"6E766572";
        ram_buffer(74659) := X"73696F6E";
        ram_buffer(74660) := X"20726571";
        ram_buffer(74661) := X"75657374";
        ram_buffer(74662) := X"00000000";
        ram_buffer(74663) := X"426F6775";
        ram_buffer(74664) := X"73204441";
        ram_buffer(74665) := X"4320696E";
        ram_buffer(74666) := X"64657820";
        ram_buffer(74667) := X"25640000";
        ram_buffer(74668) := X"426F6775";
        ram_buffer(74669) := X"73204441";
        ram_buffer(74670) := X"43207661";
        ram_buffer(74671) := X"6C756520";
        ram_buffer(74672) := X"30782578";
        ram_buffer(74673) := X"00000000";
        ram_buffer(74674) := X"426F6775";
        ram_buffer(74675) := X"73204448";
        ram_buffer(74676) := X"5420636F";
        ram_buffer(74677) := X"756E7473";
        ram_buffer(74678) := X"00000000";
        ram_buffer(74679) := X"426F6775";
        ram_buffer(74680) := X"73204448";
        ram_buffer(74681) := X"5420696E";
        ram_buffer(74682) := X"64657820";
        ram_buffer(74683) := X"25640000";
        ram_buffer(74684) := X"426F6775";
        ram_buffer(74685) := X"73204451";
        ram_buffer(74686) := X"5420696E";
        ram_buffer(74687) := X"64657820";
        ram_buffer(74688) := X"25640000";
        ram_buffer(74689) := X"456D7074";
        ram_buffer(74690) := X"79204A50";
        ram_buffer(74691) := X"45472069";
        ram_buffer(74692) := X"6D616765";
        ram_buffer(74693) := X"2028444E";
        ram_buffer(74694) := X"4C206E6F";
        ram_buffer(74695) := X"74207375";
        ram_buffer(74696) := X"70706F72";
        ram_buffer(74697) := X"74656429";
        ram_buffer(74698) := X"00000000";
        ram_buffer(74699) := X"52656164";
        ram_buffer(74700) := X"2066726F";
        ram_buffer(74701) := X"6D20454D";
        ram_buffer(74702) := X"53206661";
        ram_buffer(74703) := X"696C6564";
        ram_buffer(74704) := X"00000000";
        ram_buffer(74705) := X"57726974";
        ram_buffer(74706) := X"6520746F";
        ram_buffer(74707) := X"20454D53";
        ram_buffer(74708) := X"20666169";
        ram_buffer(74709) := X"6C656400";
        ram_buffer(74710) := X"4469646E";
        ram_buffer(74711) := X"27742065";
        ram_buffer(74712) := X"78706563";
        ram_buffer(74713) := X"74206D6F";
        ram_buffer(74714) := X"72652074";
        ram_buffer(74715) := X"68616E20";
        ram_buffer(74716) := X"6F6E6520";
        ram_buffer(74717) := X"7363616E";
        ram_buffer(74718) := X"00000000";
        ram_buffer(74719) := X"496E7075";
        ram_buffer(74720) := X"74206669";
        ram_buffer(74721) := X"6C652072";
        ram_buffer(74722) := X"65616420";
        ram_buffer(74723) := X"6572726F";
        ram_buffer(74724) := X"72000000";
        ram_buffer(74725) := X"4F757470";
        ram_buffer(74726) := X"75742066";
        ram_buffer(74727) := X"696C6520";
        ram_buffer(74728) := X"77726974";
        ram_buffer(74729) := X"65206572";
        ram_buffer(74730) := X"726F7220";
        ram_buffer(74731) := X"2D2D2D20";
        ram_buffer(74732) := X"6F757420";
        ram_buffer(74733) := X"6F662064";
        ram_buffer(74734) := X"69736B20";
        ram_buffer(74735) := X"73706163";
        ram_buffer(74736) := X"653F0000";
        ram_buffer(74737) := X"46726163";
        ram_buffer(74738) := X"74696F6E";
        ram_buffer(74739) := X"616C2073";
        ram_buffer(74740) := X"616D706C";
        ram_buffer(74741) := X"696E6720";
        ram_buffer(74742) := X"6E6F7420";
        ram_buffer(74743) := X"696D706C";
        ram_buffer(74744) := X"656D656E";
        ram_buffer(74745) := X"74656420";
        ram_buffer(74746) := X"79657400";
        ram_buffer(74747) := X"48756666";
        ram_buffer(74748) := X"6D616E20";
        ram_buffer(74749) := X"636F6465";
        ram_buffer(74750) := X"2073697A";
        ram_buffer(74751) := X"65207461";
        ram_buffer(74752) := X"626C6520";
        ram_buffer(74753) := X"6F766572";
        ram_buffer(74754) := X"666C6F77";
        ram_buffer(74755) := X"00000000";
        ram_buffer(74756) := X"4D697373";
        ram_buffer(74757) := X"696E6720";
        ram_buffer(74758) := X"48756666";
        ram_buffer(74759) := X"6D616E20";
        ram_buffer(74760) := X"636F6465";
        ram_buffer(74761) := X"20746162";
        ram_buffer(74762) := X"6C652065";
        ram_buffer(74763) := X"6E747279";
        ram_buffer(74764) := X"00000000";
        ram_buffer(74765) := X"4D617869";
        ram_buffer(74766) := X"6D756D20";
        ram_buffer(74767) := X"73757070";
        ram_buffer(74768) := X"6F727465";
        ram_buffer(74769) := X"6420696D";
        ram_buffer(74770) := X"61676520";
        ram_buffer(74771) := X"64696D65";
        ram_buffer(74772) := X"6E73696F";
        ram_buffer(74773) := X"6E206973";
        ram_buffer(74774) := X"20257520";
        ram_buffer(74775) := X"70697865";
        ram_buffer(74776) := X"6C730000";
        ram_buffer(74777) := X"456D7074";
        ram_buffer(74778) := X"7920696E";
        ram_buffer(74779) := X"70757420";
        ram_buffer(74780) := X"66696C65";
        ram_buffer(74781) := X"00000000";
        ram_buffer(74782) := X"5072656D";
        ram_buffer(74783) := X"61747572";
        ram_buffer(74784) := X"6520656E";
        ram_buffer(74785) := X"64206F66";
        ram_buffer(74786) := X"20696E70";
        ram_buffer(74787) := X"75742066";
        ram_buffer(74788) := X"696C6500";
        ram_buffer(74789) := X"43616E6E";
        ram_buffer(74790) := X"6F742074";
        ram_buffer(74791) := X"72616E73";
        ram_buffer(74792) := X"636F6465";
        ram_buffer(74793) := X"20647565";
        ram_buffer(74794) := X"20746F20";
        ram_buffer(74795) := X"6D756C74";
        ram_buffer(74796) := X"69706C65";
        ram_buffer(74797) := X"20757365";
        ram_buffer(74798) := X"206F6620";
        ram_buffer(74799) := X"7175616E";
        ram_buffer(74800) := X"74697A61";
        ram_buffer(74801) := X"74696F6E";
        ram_buffer(74802) := X"20746162";
        ram_buffer(74803) := X"6C652025";
        ram_buffer(74804) := X"64000000";
        ram_buffer(74805) := X"5363616E";
        ram_buffer(74806) := X"20736372";
        ram_buffer(74807) := X"69707420";
        ram_buffer(74808) := X"646F6573";
        ram_buffer(74809) := X"206E6F74";
        ram_buffer(74810) := X"20747261";
        ram_buffer(74811) := X"6E736D69";
        ram_buffer(74812) := X"7420616C";
        ram_buffer(74813) := X"6C206461";
        ram_buffer(74814) := X"74610000";
        ram_buffer(74815) := X"496E7661";
        ram_buffer(74816) := X"6C696420";
        ram_buffer(74817) := X"636F6C6F";
        ram_buffer(74818) := X"72207175";
        ram_buffer(74819) := X"616E7469";
        ram_buffer(74820) := X"7A617469";
        ram_buffer(74821) := X"6F6E206D";
        ram_buffer(74822) := X"6F646520";
        ram_buffer(74823) := X"6368616E";
        ram_buffer(74824) := X"67650000";
        ram_buffer(74825) := X"4E6F7420";
        ram_buffer(74826) := X"696D706C";
        ram_buffer(74827) := X"656D656E";
        ram_buffer(74828) := X"74656420";
        ram_buffer(74829) := X"79657400";
        ram_buffer(74830) := X"52657175";
        ram_buffer(74831) := X"65737465";
        ram_buffer(74832) := X"64206665";
        ram_buffer(74833) := X"61747572";
        ram_buffer(74834) := X"65207761";
        ram_buffer(74835) := X"73206F6D";
        ram_buffer(74836) := X"69747465";
        ram_buffer(74837) := X"64206174";
        ram_buffer(74838) := X"20636F6D";
        ram_buffer(74839) := X"70696C65";
        ram_buffer(74840) := X"2074696D";
        ram_buffer(74841) := X"65000000";
        ram_buffer(74842) := X"4261636B";
        ram_buffer(74843) := X"696E6720";
        ram_buffer(74844) := X"73746F72";
        ram_buffer(74845) := X"65206E6F";
        ram_buffer(74846) := X"74207375";
        ram_buffer(74847) := X"70706F72";
        ram_buffer(74848) := X"74656400";
        ram_buffer(74849) := X"48756666";
        ram_buffer(74850) := X"6D616E20";
        ram_buffer(74851) := X"7461626C";
        ram_buffer(74852) := X"65203078";
        ram_buffer(74853) := X"25303278";
        ram_buffer(74854) := X"20776173";
        ram_buffer(74855) := X"206E6F74";
        ram_buffer(74856) := X"20646566";
        ram_buffer(74857) := X"696E6564";
        ram_buffer(74858) := X"00000000";
        ram_buffer(74859) := X"4A504547";
        ram_buffer(74860) := X"20646174";
        ram_buffer(74861) := X"61737472";
        ram_buffer(74862) := X"65616D20";
        ram_buffer(74863) := X"636F6E74";
        ram_buffer(74864) := X"61696E73";
        ram_buffer(74865) := X"206E6F20";
        ram_buffer(74866) := X"696D6167";
        ram_buffer(74867) := X"65000000";
        ram_buffer(74868) := X"5175616E";
        ram_buffer(74869) := X"74697A61";
        ram_buffer(74870) := X"74696F6E";
        ram_buffer(74871) := X"20746162";
        ram_buffer(74872) := X"6C652030";
        ram_buffer(74873) := X"78253032";
        ram_buffer(74874) := X"78207761";
        ram_buffer(74875) := X"73206E6F";
        ram_buffer(74876) := X"74206465";
        ram_buffer(74877) := X"66696E65";
        ram_buffer(74878) := X"64000000";
        ram_buffer(74879) := X"4E6F7420";
        ram_buffer(74880) := X"61204A50";
        ram_buffer(74881) := X"45472066";
        ram_buffer(74882) := X"696C653A";
        ram_buffer(74883) := X"20737461";
        ram_buffer(74884) := X"72747320";
        ram_buffer(74885) := X"77697468";
        ram_buffer(74886) := X"20307825";
        ram_buffer(74887) := X"30327820";
        ram_buffer(74888) := X"30782530";
        ram_buffer(74889) := X"32780000";
        ram_buffer(74890) := X"496E7375";
        ram_buffer(74891) := X"66666963";
        ram_buffer(74892) := X"69656E74";
        ram_buffer(74893) := X"206D656D";
        ram_buffer(74894) := X"6F727920";
        ram_buffer(74895) := X"28636173";
        ram_buffer(74896) := X"65202564";
        ram_buffer(74897) := X"29000000";
        ram_buffer(74898) := X"43616E6E";
        ram_buffer(74899) := X"6F742071";
        ram_buffer(74900) := X"75616E74";
        ram_buffer(74901) := X"697A6520";
        ram_buffer(74902) := X"6D6F7265";
        ram_buffer(74903) := X"20746861";
        ram_buffer(74904) := X"6E202564";
        ram_buffer(74905) := X"20636F6C";
        ram_buffer(74906) := X"6F722063";
        ram_buffer(74907) := X"6F6D706F";
        ram_buffer(74908) := X"6E656E74";
        ram_buffer(74909) := X"73000000";
        ram_buffer(74910) := X"43616E6E";
        ram_buffer(74911) := X"6F742071";
        ram_buffer(74912) := X"75616E74";
        ram_buffer(74913) := X"697A6520";
        ram_buffer(74914) := X"746F2066";
        ram_buffer(74915) := X"65776572";
        ram_buffer(74916) := X"20746861";
        ram_buffer(74917) := X"6E202564";
        ram_buffer(74918) := X"20636F6C";
        ram_buffer(74919) := X"6F727300";
        ram_buffer(74920) := X"43616E6E";
        ram_buffer(74921) := X"6F742071";
        ram_buffer(74922) := X"75616E74";
        ram_buffer(74923) := X"697A6520";
        ram_buffer(74924) := X"746F206D";
        ram_buffer(74925) := X"6F726520";
        ram_buffer(74926) := X"7468616E";
        ram_buffer(74927) := X"20256420";
        ram_buffer(74928) := X"636F6C6F";
        ram_buffer(74929) := X"72730000";
        ram_buffer(74930) := X"496E7661";
        ram_buffer(74931) := X"6C696420";
        ram_buffer(74932) := X"4A504547";
        ram_buffer(74933) := X"2066696C";
        ram_buffer(74934) := X"65207374";
        ram_buffer(74935) := X"72756374";
        ram_buffer(74936) := X"7572653A";
        ram_buffer(74937) := X"2074776F";
        ram_buffer(74938) := X"20534F46";
        ram_buffer(74939) := X"206D6172";
        ram_buffer(74940) := X"6B657273";
        ram_buffer(74941) := X"00000000";
        ram_buffer(74942) := X"496E7661";
        ram_buffer(74943) := X"6C696420";
        ram_buffer(74944) := X"4A504547";
        ram_buffer(74945) := X"2066696C";
        ram_buffer(74946) := X"65207374";
        ram_buffer(74947) := X"72756374";
        ram_buffer(74948) := X"7572653A";
        ram_buffer(74949) := X"206D6973";
        ram_buffer(74950) := X"73696E67";
        ram_buffer(74951) := X"20534F53";
        ram_buffer(74952) := X"206D6172";
        ram_buffer(74953) := X"6B657200";
        ram_buffer(74954) := X"556E7375";
        ram_buffer(74955) := X"70706F72";
        ram_buffer(74956) := X"74656420";
        ram_buffer(74957) := X"4A504547";
        ram_buffer(74958) := X"2070726F";
        ram_buffer(74959) := X"63657373";
        ram_buffer(74960) := X"3A20534F";
        ram_buffer(74961) := X"46207479";
        ram_buffer(74962) := X"70652030";
        ram_buffer(74963) := X"78253032";
        ram_buffer(74964) := X"78000000";
        ram_buffer(74965) := X"496E7661";
        ram_buffer(74966) := X"6C696420";
        ram_buffer(74967) := X"4A504547";
        ram_buffer(74968) := X"2066696C";
        ram_buffer(74969) := X"65207374";
        ram_buffer(74970) := X"72756374";
        ram_buffer(74971) := X"7572653A";
        ram_buffer(74972) := X"2074776F";
        ram_buffer(74973) := X"20534F49";
        ram_buffer(74974) := X"206D6172";
        ram_buffer(74975) := X"6B657273";
        ram_buffer(74976) := X"00000000";
        ram_buffer(74977) := X"496E7661";
        ram_buffer(74978) := X"6C696420";
        ram_buffer(74979) := X"4A504547";
        ram_buffer(74980) := X"2066696C";
        ram_buffer(74981) := X"65207374";
        ram_buffer(74982) := X"72756374";
        ram_buffer(74983) := X"7572653A";
        ram_buffer(74984) := X"20534F53";
        ram_buffer(74985) := X"20626566";
        ram_buffer(74986) := X"6F726520";
        ram_buffer(74987) := X"534F4600";
        ram_buffer(74988) := X"4661696C";
        ram_buffer(74989) := X"65642074";
        ram_buffer(74990) := X"6F206372";
        ram_buffer(74991) := X"65617465";
        ram_buffer(74992) := X"2074656D";
        ram_buffer(74993) := X"706F7261";
        ram_buffer(74994) := X"72792066";
        ram_buffer(74995) := X"696C6520";
        ram_buffer(74996) := X"25730000";
        ram_buffer(74997) := X"52656164";
        ram_buffer(74998) := X"20666169";
        ram_buffer(74999) := X"6C656420";
        ram_buffer(75000) := X"6F6E2074";
        ram_buffer(75001) := X"656D706F";
        ram_buffer(75002) := X"72617279";
        ram_buffer(75003) := X"2066696C";
        ram_buffer(75004) := X"65000000";
        ram_buffer(75005) := X"5365656B";
        ram_buffer(75006) := X"20666169";
        ram_buffer(75007) := X"6C656420";
        ram_buffer(75008) := X"6F6E2074";
        ram_buffer(75009) := X"656D706F";
        ram_buffer(75010) := X"72617279";
        ram_buffer(75011) := X"2066696C";
        ram_buffer(75012) := X"65000000";
        ram_buffer(75013) := X"57726974";
        ram_buffer(75014) := X"65206661";
        ram_buffer(75015) := X"696C6564";
        ram_buffer(75016) := X"206F6E20";
        ram_buffer(75017) := X"74656D70";
        ram_buffer(75018) := X"6F726172";
        ram_buffer(75019) := X"79206669";
        ram_buffer(75020) := X"6C65202D";
        ram_buffer(75021) := X"2D2D206F";
        ram_buffer(75022) := X"7574206F";
        ram_buffer(75023) := X"66206469";
        ram_buffer(75024) := X"736B2073";
        ram_buffer(75025) := X"70616365";
        ram_buffer(75026) := X"3F000000";
        ram_buffer(75027) := X"4170706C";
        ram_buffer(75028) := X"69636174";
        ram_buffer(75029) := X"696F6E20";
        ram_buffer(75030) := X"7472616E";
        ram_buffer(75031) := X"73666572";
        ram_buffer(75032) := X"72656420";
        ram_buffer(75033) := X"746F6F20";
        ram_buffer(75034) := X"66657720";
        ram_buffer(75035) := X"7363616E";
        ram_buffer(75036) := X"6C696E65";
        ram_buffer(75037) := X"73000000";
        ram_buffer(75038) := X"556E7375";
        ram_buffer(75039) := X"70706F72";
        ram_buffer(75040) := X"74656420";
        ram_buffer(75041) := X"6D61726B";
        ram_buffer(75042) := X"65722074";
        ram_buffer(75043) := X"79706520";
        ram_buffer(75044) := X"30782530";
        ram_buffer(75045) := X"32780000";
        ram_buffer(75046) := X"56697274";
        ram_buffer(75047) := X"75616C20";
        ram_buffer(75048) := X"61727261";
        ram_buffer(75049) := X"7920636F";
        ram_buffer(75050) := X"6E74726F";
        ram_buffer(75051) := X"6C6C6572";
        ram_buffer(75052) := X"206D6573";
        ram_buffer(75053) := X"73656420";
        ram_buffer(75054) := X"75700000";
        ram_buffer(75055) := X"496D6167";
        ram_buffer(75056) := X"6520746F";
        ram_buffer(75057) := X"6F207769";
        ram_buffer(75058) := X"64652066";
        ram_buffer(75059) := X"6F722074";
        ram_buffer(75060) := X"68697320";
        ram_buffer(75061) := X"696D706C";
        ram_buffer(75062) := X"656D656E";
        ram_buffer(75063) := X"74617469";
        ram_buffer(75064) := X"6F6E0000";
        ram_buffer(75065) := X"52656164";
        ram_buffer(75066) := X"2066726F";
        ram_buffer(75067) := X"6D20584D";
        ram_buffer(75068) := X"53206661";
        ram_buffer(75069) := X"696C6564";
        ram_buffer(75070) := X"00000000";
        ram_buffer(75071) := X"57726974";
        ram_buffer(75072) := X"6520746F";
        ram_buffer(75073) := X"20584D53";
        ram_buffer(75074) := X"20666169";
        ram_buffer(75075) := X"6C656400";
        ram_buffer(75076) := X"43617574";
        ram_buffer(75077) := X"696F6E3A";
        ram_buffer(75078) := X"20717561";
        ram_buffer(75079) := X"6E74697A";
        ram_buffer(75080) := X"6174696F";
        ram_buffer(75081) := X"6E207461";
        ram_buffer(75082) := X"626C6573";
        ram_buffer(75083) := X"20617265";
        ram_buffer(75084) := X"20746F6F";
        ram_buffer(75085) := X"20636F61";
        ram_buffer(75086) := X"72736520";
        ram_buffer(75087) := X"666F7220";
        ram_buffer(75088) := X"62617365";
        ram_buffer(75089) := X"6C696E65";
        ram_buffer(75090) := X"204A5045";
        ram_buffer(75091) := X"47000000";
        ram_buffer(75092) := X"41646F62";
        ram_buffer(75093) := X"65204150";
        ram_buffer(75094) := X"50313420";
        ram_buffer(75095) := X"6D61726B";
        ram_buffer(75096) := X"65723A20";
        ram_buffer(75097) := X"76657273";
        ram_buffer(75098) := X"696F6E20";
        ram_buffer(75099) := X"25642C20";
        ram_buffer(75100) := X"666C6167";
        ram_buffer(75101) := X"73203078";
        ram_buffer(75102) := X"25303478";
        ram_buffer(75103) := X"20307825";
        ram_buffer(75104) := X"3034782C";
        ram_buffer(75105) := X"20747261";
        ram_buffer(75106) := X"6E73666F";
        ram_buffer(75107) := X"726D2025";
        ram_buffer(75108) := X"64000000";
        ram_buffer(75109) := X"556E6B6E";
        ram_buffer(75110) := X"6F776E20";
        ram_buffer(75111) := X"41505030";
        ram_buffer(75112) := X"206D6172";
        ram_buffer(75113) := X"6B657220";
        ram_buffer(75114) := X"286E6F74";
        ram_buffer(75115) := X"204A4649";
        ram_buffer(75116) := X"46292C20";
        ram_buffer(75117) := X"6C656E67";
        ram_buffer(75118) := X"74682025";
        ram_buffer(75119) := X"75000000";
        ram_buffer(75120) := X"556E6B6E";
        ram_buffer(75121) := X"6F776E20";
        ram_buffer(75122) := X"41505031";
        ram_buffer(75123) := X"34206D61";
        ram_buffer(75124) := X"726B6572";
        ram_buffer(75125) := X"20286E6F";
        ram_buffer(75126) := X"74204164";
        ram_buffer(75127) := X"6F626529";
        ram_buffer(75128) := X"2C206C65";
        ram_buffer(75129) := X"6E677468";
        ram_buffer(75130) := X"20257500";
        ram_buffer(75131) := X"44656669";
        ram_buffer(75132) := X"6E652041";
        ram_buffer(75133) := X"72697468";
        ram_buffer(75134) := X"6D657469";
        ram_buffer(75135) := X"63205461";
        ram_buffer(75136) := X"626C6520";
        ram_buffer(75137) := X"30782530";
        ram_buffer(75138) := X"32783A20";
        ram_buffer(75139) := X"30782530";
        ram_buffer(75140) := X"32780000";
        ram_buffer(75141) := X"44656669";
        ram_buffer(75142) := X"6E652048";
        ram_buffer(75143) := X"7566666D";
        ram_buffer(75144) := X"616E2054";
        ram_buffer(75145) := X"61626C65";
        ram_buffer(75146) := X"20307825";
        ram_buffer(75147) := X"30327800";
        ram_buffer(75148) := X"44656669";
        ram_buffer(75149) := X"6E652051";
        ram_buffer(75150) := X"75616E74";
        ram_buffer(75151) := X"697A6174";
        ram_buffer(75152) := X"696F6E20";
        ram_buffer(75153) := X"5461626C";
        ram_buffer(75154) := X"65202564";
        ram_buffer(75155) := X"20207072";
        ram_buffer(75156) := X"65636973";
        ram_buffer(75157) := X"696F6E20";
        ram_buffer(75158) := X"25640000";
        ram_buffer(75159) := X"44656669";
        ram_buffer(75160) := X"6E652052";
        ram_buffer(75161) := X"65737461";
        ram_buffer(75162) := X"72742049";
        ram_buffer(75163) := X"6E746572";
        ram_buffer(75164) := X"76616C20";
        ram_buffer(75165) := X"25750000";
        ram_buffer(75166) := X"46726565";
        ram_buffer(75167) := X"6420454D";
        ram_buffer(75168) := X"53206861";
        ram_buffer(75169) := X"6E646C65";
        ram_buffer(75170) := X"20257500";
        ram_buffer(75171) := X"4F627461";
        ram_buffer(75172) := X"696E6564";
        ram_buffer(75173) := X"20454D53";
        ram_buffer(75174) := X"2068616E";
        ram_buffer(75175) := X"646C6520";
        ram_buffer(75176) := X"25750000";
        ram_buffer(75177) := X"456E6420";
        ram_buffer(75178) := X"4F662049";
        ram_buffer(75179) := X"6D616765";
        ram_buffer(75180) := X"00000000";
        ram_buffer(75181) := X"20202020";
        ram_buffer(75182) := X"20202020";
        ram_buffer(75183) := X"25336420";
        ram_buffer(75184) := X"25336420";
        ram_buffer(75185) := X"25336420";
        ram_buffer(75186) := X"25336420";
        ram_buffer(75187) := X"25336420";
        ram_buffer(75188) := X"25336420";
        ram_buffer(75189) := X"25336420";
        ram_buffer(75190) := X"25336400";
        ram_buffer(75191) := X"4A464946";
        ram_buffer(75192) := X"20415050";
        ram_buffer(75193) := X"30206D61";
        ram_buffer(75194) := X"726B6572";
        ram_buffer(75195) := X"2C206465";
        ram_buffer(75196) := X"6E736974";
        ram_buffer(75197) := X"79202564";
        ram_buffer(75198) := X"78256420";
        ram_buffer(75199) := X"20256400";
        ram_buffer(75200) := X"5761726E";
        ram_buffer(75201) := X"696E673A";
        ram_buffer(75202) := X"20746875";
        ram_buffer(75203) := X"6D626E61";
        ram_buffer(75204) := X"696C2069";
        ram_buffer(75205) := X"6D616765";
        ram_buffer(75206) := X"2073697A";
        ram_buffer(75207) := X"6520646F";
        ram_buffer(75208) := X"6573206E";
        ram_buffer(75209) := X"6F74206D";
        ram_buffer(75210) := X"61746368";
        ram_buffer(75211) := X"20646174";
        ram_buffer(75212) := X"61206C65";
        ram_buffer(75213) := X"6E677468";
        ram_buffer(75214) := X"20257500";
        ram_buffer(75215) := X"556E6B6E";
        ram_buffer(75216) := X"6F776E20";
        ram_buffer(75217) := X"4A464946";
        ram_buffer(75218) := X"206D696E";
        ram_buffer(75219) := X"6F722072";
        ram_buffer(75220) := X"65766973";
        ram_buffer(75221) := X"696F6E20";
        ram_buffer(75222) := X"6E756D62";
        ram_buffer(75223) := X"65722025";
        ram_buffer(75224) := X"642E2530";
        ram_buffer(75225) := X"32640000";
        ram_buffer(75226) := X"20202020";
        ram_buffer(75227) := X"77697468";
        ram_buffer(75228) := X"20256420";
        ram_buffer(75229) := X"78202564";
        ram_buffer(75230) := X"20746875";
        ram_buffer(75231) := X"6D626E61";
        ram_buffer(75232) := X"696C2069";
        ram_buffer(75233) := X"6D616765";
        ram_buffer(75234) := X"00000000";
        ram_buffer(75235) := X"536B6970";
        ram_buffer(75236) := X"70696E67";
        ram_buffer(75237) := X"206D6172";
        ram_buffer(75238) := X"6B657220";
        ram_buffer(75239) := X"30782530";
        ram_buffer(75240) := X"32782C20";
        ram_buffer(75241) := X"6C656E67";
        ram_buffer(75242) := X"74682025";
        ram_buffer(75243) := X"75000000";
        ram_buffer(75244) := X"556E6578";
        ram_buffer(75245) := X"70656374";
        ram_buffer(75246) := X"6564206D";
        ram_buffer(75247) := X"61726B65";
        ram_buffer(75248) := X"72203078";
        ram_buffer(75249) := X"25303278";
        ram_buffer(75250) := X"00000000";
        ram_buffer(75251) := X"20202020";
        ram_buffer(75252) := X"20202020";
        ram_buffer(75253) := X"25347520";
        ram_buffer(75254) := X"25347520";
        ram_buffer(75255) := X"25347520";
        ram_buffer(75256) := X"25347520";
        ram_buffer(75257) := X"25347520";
        ram_buffer(75258) := X"25347520";
        ram_buffer(75259) := X"25347520";
        ram_buffer(75260) := X"25347500";
        ram_buffer(75261) := X"5175616E";
        ram_buffer(75262) := X"74697A69";
        ram_buffer(75263) := X"6E672074";
        ram_buffer(75264) := X"6F202564";
        ram_buffer(75265) := X"203D2025";
        ram_buffer(75266) := X"642A2564";
        ram_buffer(75267) := X"2A256420";
        ram_buffer(75268) := X"636F6C6F";
        ram_buffer(75269) := X"72730000";
        ram_buffer(75270) := X"5175616E";
        ram_buffer(75271) := X"74697A69";
        ram_buffer(75272) := X"6E672074";
        ram_buffer(75273) := X"6F202564";
        ram_buffer(75274) := X"20636F6C";
        ram_buffer(75275) := X"6F727300";
        ram_buffer(75276) := X"53656C65";
        ram_buffer(75277) := X"63746564";
        ram_buffer(75278) := X"20256420";
        ram_buffer(75279) := X"636F6C6F";
        ram_buffer(75280) := X"72732066";
        ram_buffer(75281) := X"6F722071";
        ram_buffer(75282) := X"75616E74";
        ram_buffer(75283) := X"697A6174";
        ram_buffer(75284) := X"696F6E00";
        ram_buffer(75285) := X"4174206D";
        ram_buffer(75286) := X"61726B65";
        ram_buffer(75287) := X"72203078";
        ram_buffer(75288) := X"25303278";
        ram_buffer(75289) := X"2C207265";
        ram_buffer(75290) := X"636F7665";
        ram_buffer(75291) := X"72792061";
        ram_buffer(75292) := X"6374696F";
        ram_buffer(75293) := X"6E202564";
        ram_buffer(75294) := X"00000000";
        ram_buffer(75295) := X"52535425";
        ram_buffer(75296) := X"64000000";
        ram_buffer(75297) := X"536D6F6F";
        ram_buffer(75298) := X"7468696E";
        ram_buffer(75299) := X"67206E6F";
        ram_buffer(75300) := X"74207375";
        ram_buffer(75301) := X"70706F72";
        ram_buffer(75302) := X"74656420";
        ram_buffer(75303) := X"77697468";
        ram_buffer(75304) := X"206E6F6E";
        ram_buffer(75305) := X"7374616E";
        ram_buffer(75306) := X"64617264";
        ram_buffer(75307) := X"2073616D";
        ram_buffer(75308) := X"706C696E";
        ram_buffer(75309) := X"67207261";
        ram_buffer(75310) := X"74696F73";
        ram_buffer(75311) := X"00000000";
        ram_buffer(75312) := X"53746172";
        ram_buffer(75313) := X"74204F66";
        ram_buffer(75314) := X"20467261";
        ram_buffer(75315) := X"6D652030";
        ram_buffer(75316) := X"78253032";
        ram_buffer(75317) := X"783A2077";
        ram_buffer(75318) := X"69647468";
        ram_buffer(75319) := X"3D25752C";
        ram_buffer(75320) := X"20686569";
        ram_buffer(75321) := X"6768743D";
        ram_buffer(75322) := X"25752C20";
        ram_buffer(75323) := X"636F6D70";
        ram_buffer(75324) := X"6F6E656E";
        ram_buffer(75325) := X"74733D25";
        ram_buffer(75326) := X"64000000";
        ram_buffer(75327) := X"20202020";
        ram_buffer(75328) := X"436F6D70";
        ram_buffer(75329) := X"6F6E656E";
        ram_buffer(75330) := X"74202564";
        ram_buffer(75331) := X"3A202564";
        ram_buffer(75332) := X"68782564";
        ram_buffer(75333) := X"7620713D";
        ram_buffer(75334) := X"25640000";
        ram_buffer(75335) := X"53746172";
        ram_buffer(75336) := X"74206F66";
        ram_buffer(75337) := X"20496D61";
        ram_buffer(75338) := X"67650000";
        ram_buffer(75339) := X"53746172";
        ram_buffer(75340) := X"74204F66";
        ram_buffer(75341) := X"20536361";
        ram_buffer(75342) := X"6E3A2025";
        ram_buffer(75343) := X"6420636F";
        ram_buffer(75344) := X"6D706F6E";
        ram_buffer(75345) := X"656E7473";
        ram_buffer(75346) := X"00000000";
        ram_buffer(75347) := X"20202020";
        ram_buffer(75348) := X"436F6D70";
        ram_buffer(75349) := X"6F6E656E";
        ram_buffer(75350) := X"74202564";
        ram_buffer(75351) := X"3A206463";
        ram_buffer(75352) := X"3D256420";
        ram_buffer(75353) := X"61633D25";
        ram_buffer(75354) := X"64000000";
        ram_buffer(75355) := X"20205373";
        ram_buffer(75356) := X"3D25642C";
        ram_buffer(75357) := X"2053653D";
        ram_buffer(75358) := X"25642C20";
        ram_buffer(75359) := X"41683D25";
        ram_buffer(75360) := X"642C2041";
        ram_buffer(75361) := X"6C3D2564";
        ram_buffer(75362) := X"00000000";
        ram_buffer(75363) := X"436C6F73";
        ram_buffer(75364) := X"65642074";
        ram_buffer(75365) := X"656D706F";
        ram_buffer(75366) := X"72617279";
        ram_buffer(75367) := X"2066696C";
        ram_buffer(75368) := X"65202573";
        ram_buffer(75369) := X"00000000";
        ram_buffer(75370) := X"4F70656E";
        ram_buffer(75371) := X"65642074";
        ram_buffer(75372) := X"656D706F";
        ram_buffer(75373) := X"72617279";
        ram_buffer(75374) := X"2066696C";
        ram_buffer(75375) := X"65202573";
        ram_buffer(75376) := X"00000000";
        ram_buffer(75377) := X"556E7265";
        ram_buffer(75378) := X"636F676E";
        ram_buffer(75379) := X"697A6564";
        ram_buffer(75380) := X"20636F6D";
        ram_buffer(75381) := X"706F6E65";
        ram_buffer(75382) := X"6E742049";
        ram_buffer(75383) := X"44732025";
        ram_buffer(75384) := X"64202564";
        ram_buffer(75385) := X"2025642C";
        ram_buffer(75386) := X"20617373";
        ram_buffer(75387) := X"756D696E";
        ram_buffer(75388) := X"67205943";
        ram_buffer(75389) := X"62437200";
        ram_buffer(75390) := X"46726565";
        ram_buffer(75391) := X"6420584D";
        ram_buffer(75392) := X"53206861";
        ram_buffer(75393) := X"6E646C65";
        ram_buffer(75394) := X"20257500";
        ram_buffer(75395) := X"4F627461";
        ram_buffer(75396) := X"696E6564";
        ram_buffer(75397) := X"20584D53";
        ram_buffer(75398) := X"2068616E";
        ram_buffer(75399) := X"646C6520";
        ram_buffer(75400) := X"25750000";
        ram_buffer(75401) := X"556E6B6E";
        ram_buffer(75402) := X"6F776E20";
        ram_buffer(75403) := X"41646F62";
        ram_buffer(75404) := X"6520636F";
        ram_buffer(75405) := X"6C6F7220";
        ram_buffer(75406) := X"7472616E";
        ram_buffer(75407) := X"73666F72";
        ram_buffer(75408) := X"6D20636F";
        ram_buffer(75409) := X"64652025";
        ram_buffer(75410) := X"64000000";
        ram_buffer(75411) := X"496E636F";
        ram_buffer(75412) := X"6E736973";
        ram_buffer(75413) := X"74656E74";
        ram_buffer(75414) := X"2070726F";
        ram_buffer(75415) := X"67726573";
        ram_buffer(75416) := X"73696F6E";
        ram_buffer(75417) := X"20736571";
        ram_buffer(75418) := X"75656E63";
        ram_buffer(75419) := X"6520666F";
        ram_buffer(75420) := X"7220636F";
        ram_buffer(75421) := X"6D706F6E";
        ram_buffer(75422) := X"656E7420";
        ram_buffer(75423) := X"25642063";
        ram_buffer(75424) := X"6F656666";
        ram_buffer(75425) := X"69636965";
        ram_buffer(75426) := X"6E742025";
        ram_buffer(75427) := X"64000000";
        ram_buffer(75428) := X"436F7272";
        ram_buffer(75429) := X"75707420";
        ram_buffer(75430) := X"4A504547";
        ram_buffer(75431) := X"20646174";
        ram_buffer(75432) := X"613A2025";
        ram_buffer(75433) := X"75206578";
        ram_buffer(75434) := X"7472616E";
        ram_buffer(75435) := X"656F7573";
        ram_buffer(75436) := X"20627974";
        ram_buffer(75437) := X"65732062";
        ram_buffer(75438) := X"65666F72";
        ram_buffer(75439) := X"65206D61";
        ram_buffer(75440) := X"726B6572";
        ram_buffer(75441) := X"20307825";
        ram_buffer(75442) := X"30327800";
        ram_buffer(75443) := X"436F7272";
        ram_buffer(75444) := X"75707420";
        ram_buffer(75445) := X"4A504547";
        ram_buffer(75446) := X"20646174";
        ram_buffer(75447) := X"613A2070";
        ram_buffer(75448) := X"72656D61";
        ram_buffer(75449) := X"74757265";
        ram_buffer(75450) := X"20656E64";
        ram_buffer(75451) := X"206F6620";
        ram_buffer(75452) := X"64617461";
        ram_buffer(75453) := X"20736567";
        ram_buffer(75454) := X"6D656E74";
        ram_buffer(75455) := X"00000000";
        ram_buffer(75456) := X"436F7272";
        ram_buffer(75457) := X"75707420";
        ram_buffer(75458) := X"4A504547";
        ram_buffer(75459) := X"20646174";
        ram_buffer(75460) := X"613A2062";
        ram_buffer(75461) := X"61642048";
        ram_buffer(75462) := X"7566666D";
        ram_buffer(75463) := X"616E2063";
        ram_buffer(75464) := X"6F646500";
        ram_buffer(75465) := X"5761726E";
        ram_buffer(75466) := X"696E673A";
        ram_buffer(75467) := X"20756E6B";
        ram_buffer(75468) := X"6E6F776E";
        ram_buffer(75469) := X"204A4649";
        ram_buffer(75470) := X"46207265";
        ram_buffer(75471) := X"76697369";
        ram_buffer(75472) := X"6F6E206E";
        ram_buffer(75473) := X"756D6265";
        ram_buffer(75474) := X"72202564";
        ram_buffer(75475) := X"2E253032";
        ram_buffer(75476) := X"64000000";
        ram_buffer(75477) := X"5072656D";
        ram_buffer(75478) := X"61747572";
        ram_buffer(75479) := X"6520656E";
        ram_buffer(75480) := X"64206F66";
        ram_buffer(75481) := X"204A5045";
        ram_buffer(75482) := X"47206669";
        ram_buffer(75483) := X"6C650000";
        ram_buffer(75484) := X"436F7272";
        ram_buffer(75485) := X"75707420";
        ram_buffer(75486) := X"4A504547";
        ram_buffer(75487) := X"20646174";
        ram_buffer(75488) := X"613A2066";
        ram_buffer(75489) := X"6F756E64";
        ram_buffer(75490) := X"206D6172";
        ram_buffer(75491) := X"6B657220";
        ram_buffer(75492) := X"30782530";
        ram_buffer(75493) := X"32782069";
        ram_buffer(75494) := X"6E737465";
        ram_buffer(75495) := X"6164206F";
        ram_buffer(75496) := X"66205253";
        ram_buffer(75497) := X"54256400";
        ram_buffer(75498) := X"496E7661";
        ram_buffer(75499) := X"6C696420";
        ram_buffer(75500) := X"534F5320";
        ram_buffer(75501) := X"70617261";
        ram_buffer(75502) := X"6D657465";
        ram_buffer(75503) := X"72732066";
        ram_buffer(75504) := X"6F722073";
        ram_buffer(75505) := X"65717565";
        ram_buffer(75506) := X"6E746961";
        ram_buffer(75507) := X"6C204A50";
        ram_buffer(75508) := X"45470000";
        ram_buffer(75509) := X"4170706C";
        ram_buffer(75510) := X"69636174";
        ram_buffer(75511) := X"696F6E20";
        ram_buffer(75512) := X"7472616E";
        ram_buffer(75513) := X"73666572";
        ram_buffer(75514) := X"72656420";
        ram_buffer(75515) := X"746F6F20";
        ram_buffer(75516) := X"6D616E79";
        ram_buffer(75517) := X"20736361";
        ram_buffer(75518) := X"6E6C696E";
        ram_buffer(75519) := X"65730000";
        ram_buffer(75520) := X"100C8AA8";
        ram_buffer(75521) := X"100C8AC0";
        ram_buffer(75522) := X"100C8AFC";
        ram_buffer(75523) := X"100C8B1C";
        ram_buffer(75524) := X"100C8B44";
        ram_buffer(75525) := X"100C8B60";
        ram_buffer(75526) := X"100C8B80";
        ram_buffer(75527) := X"100C8BA8";
        ram_buffer(75528) := X"100C8BC0";
        ram_buffer(75529) := X"100C8BD8";
        ram_buffer(75530) := X"100C8BEC";
        ram_buffer(75531) := X"100C8C2C";
        ram_buffer(75532) := X"100C8C5C";
        ram_buffer(75533) := X"100C8C78";
        ram_buffer(75534) := X"100C8C9C";
        ram_buffer(75535) := X"100C8CD4";
        ram_buffer(75536) := X"100C8D0C";
        ram_buffer(75537) := X"100C8D24";
        ram_buffer(75538) := X"100C8D44";
        ram_buffer(75539) := X"100C8D70";
        ram_buffer(75540) := X"100C8DC0";
        ram_buffer(75541) := X"100C8DDC";
        ram_buffer(75542) := X"100C8E08";
        ram_buffer(75543) := X"100C8E24";
        ram_buffer(75544) := X"100C8E4C";
        ram_buffer(75545) := X"100C8E74";
        ram_buffer(75546) := X"100C8E9C";
        ram_buffer(75547) := X"100C8EB0";
        ram_buffer(75548) := X"100C8EC8";
        ram_buffer(75549) := X"100C8EDC";
        ram_buffer(75550) := X"100C8EF0";
        ram_buffer(75551) := X"100C8F04";
        ram_buffer(75552) := X"100C8F2C";
        ram_buffer(75553) := X"100C8F44";
        ram_buffer(75554) := X"100C8F58";
        ram_buffer(75555) := X"100C8F7C";
        ram_buffer(75556) := X"100C8F94";
        ram_buffer(75557) := X"100C8FC4";
        ram_buffer(75558) := X"100C8FEC";
        ram_buffer(75559) := X"100C9010";
        ram_buffer(75560) := X"100C9034";
        ram_buffer(75561) := X"100C9064";
        ram_buffer(75562) := X"100C9078";
        ram_buffer(75563) := X"100C9094";
        ram_buffer(75564) := X"100C90D4";
        ram_buffer(75565) := X"100C90FC";
        ram_buffer(75566) := X"100C9124";
        ram_buffer(75567) := X"100C9138";
        ram_buffer(75568) := X"100C9168";
        ram_buffer(75569) := X"100C9184";
        ram_buffer(75570) := X"100C91AC";
        ram_buffer(75571) := X"100C91D0";
        ram_buffer(75572) := X"100C91FC";
        ram_buffer(75573) := X"100C9228";
        ram_buffer(75574) := X"100C9248";
        ram_buffer(75575) := X"100C9278";
        ram_buffer(75576) := X"100C92A0";
        ram_buffer(75577) := X"100C92C8";
        ram_buffer(75578) := X"100C92F8";
        ram_buffer(75579) := X"100C9328";
        ram_buffer(75580) := X"100C9354";
        ram_buffer(75581) := X"100C9384";
        ram_buffer(75582) := X"100C93B0";
        ram_buffer(75583) := X"100C93D4";
        ram_buffer(75584) := X"100C93F4";
        ram_buffer(75585) := X"100C9414";
        ram_buffer(75586) := X"100C944C";
        ram_buffer(75587) := X"100C9478";
        ram_buffer(75588) := X"100C9498";
        ram_buffer(75589) := X"100C94BC";
        ram_buffer(75590) := X"100C94E4";
        ram_buffer(75591) := X"100C94FC";
        ram_buffer(75592) := X"100C7AD0";
        ram_buffer(75593) := X"100C7AF4";
        ram_buffer(75594) := X"100C9510";
        ram_buffer(75595) := X"100C9550";
        ram_buffer(75596) := X"100C9594";
        ram_buffer(75597) := X"100C95C0";
        ram_buffer(75598) := X"100C95EC";
        ram_buffer(75599) := X"100C9614";
        ram_buffer(75600) := X"100C9630";
        ram_buffer(75601) := X"100C965C";
        ram_buffer(75602) := X"100C9678";
        ram_buffer(75603) := X"100C968C";
        ram_buffer(75604) := X"100C96A4";
        ram_buffer(75605) := X"100C96B4";
        ram_buffer(75606) := X"100C96DC";
        ram_buffer(75607) := X"100C9700";
        ram_buffer(75608) := X"100C973C";
        ram_buffer(75609) := X"100C9768";
        ram_buffer(75610) := X"100C978C";
        ram_buffer(75611) := X"100C97B0";
        ram_buffer(75612) := X"100C97CC";
        ram_buffer(75613) := X"100C97F4";
        ram_buffer(75614) := X"100C9818";
        ram_buffer(75615) := X"100C9830";
        ram_buffer(75616) := X"100C9854";
        ram_buffer(75617) := X"100C987C";
        ram_buffer(75618) := X"100C9884";
        ram_buffer(75619) := X"100C98C0";
        ram_buffer(75620) := X"100C98FC";
        ram_buffer(75621) := X"100C991C";
        ram_buffer(75622) := X"100C992C";
        ram_buffer(75623) := X"100C994C";
        ram_buffer(75624) := X"100C996C";
        ram_buffer(75625) := X"100C998C";
        ram_buffer(75626) := X"100C99A8";
        ram_buffer(75627) := X"100C99C4";
        ram_buffer(75628) := X"100C99F8";
        ram_buffer(75629) := X"100C9A0C";
        ram_buffer(75630) := X"100C9A24";
        ram_buffer(75631) := X"100C9A4C";
        ram_buffer(75632) := X"100C9A90";
        ram_buffer(75633) := X"100C9ACC";
        ram_buffer(75634) := X"100C9B00";
        ram_buffer(75635) := X"100C9B24";
        ram_buffer(75636) := X"100C9B54";
        ram_buffer(75637) := X"100C9B70";
        ram_buffer(75638) := X"100C9BA8";
        ram_buffer(75639) := X"100C9BD4";
        ram_buffer(75640) := X"00000000";
        ram_buffer(75641) := X"4A504547";
        ram_buffer(75642) := X"4D454D00";
        ram_buffer(75643) := X"00000000";
        ram_buffer(75644) := X"00000000";
        ram_buffer(75645) := X"00000000";
        ram_buffer(75646) := X"00000000";
        ram_buffer(75647) := X"00000000";
        ram_buffer(75648) := X"00000000";
        ram_buffer(75649) := X"00000000";
        ram_buffer(75650) := X"00000000";
        ram_buffer(75651) := X"00000000";
        ram_buffer(75652) := X"00000000";
        ram_buffer(75653) := X"00000000";
        ram_buffer(75654) := X"00000000";
        ram_buffer(75655) := X"00000000";
        ram_buffer(75656) := X"00000000";
        ram_buffer(75657) := X"00000000";
        ram_buffer(75658) := X"00000000";
        ram_buffer(75659) := X"00000000";
        ram_buffer(75660) := X"00000000";
        ram_buffer(75661) := X"00000000";
        ram_buffer(75662) := X"00000000";
        ram_buffer(75663) := X"00000000";
        ram_buffer(75664) := X"00000000";
        ram_buffer(75665) := X"00000000";
        ram_buffer(75666) := X"00000000";
        ram_buffer(75667) := X"00000000";
        ram_buffer(75668) := X"00000000";
        ram_buffer(75669) := X"00000000";
        ram_buffer(75670) := X"00000000";
        ram_buffer(75671) := X"00000000";
        ram_buffer(75672) := X"00000000";
        ram_buffer(75673) := X"00000000";
        ram_buffer(75674) := X"00000000";
        ram_buffer(75675) := X"20202020";
        ram_buffer(75676) := X"20202020";
        ram_buffer(75677) := X"20282828";
        ram_buffer(75678) := X"28282020";
        ram_buffer(75679) := X"20202020";
        ram_buffer(75680) := X"20202020";
        ram_buffer(75681) := X"20202020";
        ram_buffer(75682) := X"20202020";
        ram_buffer(75683) := X"88101010";
        ram_buffer(75684) := X"10101010";
        ram_buffer(75685) := X"10101010";
        ram_buffer(75686) := X"10101010";
        ram_buffer(75687) := X"04040404";
        ram_buffer(75688) := X"04040404";
        ram_buffer(75689) := X"04041010";
        ram_buffer(75690) := X"10101010";
        ram_buffer(75691) := X"10414141";
        ram_buffer(75692) := X"41414101";
        ram_buffer(75693) := X"01010101";
        ram_buffer(75694) := X"01010101";
        ram_buffer(75695) := X"01010101";
        ram_buffer(75696) := X"01010101";
        ram_buffer(75697) := X"01010110";
        ram_buffer(75698) := X"10101010";
        ram_buffer(75699) := X"10424242";
        ram_buffer(75700) := X"42424202";
        ram_buffer(75701) := X"02020202";
        ram_buffer(75702) := X"02020202";
        ram_buffer(75703) := X"02020202";
        ram_buffer(75704) := X"02020202";
        ram_buffer(75705) := X"02020210";
        ram_buffer(75706) := X"10101020";
        ram_buffer(75707) := X"00000000";
        ram_buffer(75708) := X"00000000";
        ram_buffer(75709) := X"00000000";
        ram_buffer(75710) := X"00000000";
        ram_buffer(75711) := X"00000000";
        ram_buffer(75712) := X"00000000";
        ram_buffer(75713) := X"00000000";
        ram_buffer(75714) := X"00000000";
        ram_buffer(75715) := X"00000000";
        ram_buffer(75716) := X"00000000";
        ram_buffer(75717) := X"00000000";
        ram_buffer(75718) := X"00000000";
        ram_buffer(75719) := X"00000000";
        ram_buffer(75720) := X"00000000";
        ram_buffer(75721) := X"00000000";
        ram_buffer(75722) := X"00000000";
        ram_buffer(75723) := X"00000000";
        ram_buffer(75724) := X"00000000";
        ram_buffer(75725) := X"00000000";
        ram_buffer(75726) := X"00000000";
        ram_buffer(75727) := X"00000000";
        ram_buffer(75728) := X"00000000";
        ram_buffer(75729) := X"00000000";
        ram_buffer(75730) := X"00000000";
        ram_buffer(75731) := X"00000000";
        ram_buffer(75732) := X"00000000";
        ram_buffer(75733) := X"00000000";
        ram_buffer(75734) := X"00000000";
        ram_buffer(75735) := X"00000000";
        ram_buffer(75736) := X"00000000";
        ram_buffer(75737) := X"00000000";
        ram_buffer(75738) := X"00000000";
        ram_buffer(75739) := X"00202020";
        ram_buffer(75740) := X"20202020";
        ram_buffer(75741) := X"20202828";
        ram_buffer(75742) := X"28282820";
        ram_buffer(75743) := X"20202020";
        ram_buffer(75744) := X"20202020";
        ram_buffer(75745) := X"20202020";
        ram_buffer(75746) := X"20202020";
        ram_buffer(75747) := X"20881010";
        ram_buffer(75748) := X"10101010";
        ram_buffer(75749) := X"10101010";
        ram_buffer(75750) := X"10101010";
        ram_buffer(75751) := X"10040404";
        ram_buffer(75752) := X"04040404";
        ram_buffer(75753) := X"04040410";
        ram_buffer(75754) := X"10101010";
        ram_buffer(75755) := X"10104141";
        ram_buffer(75756) := X"41414141";
        ram_buffer(75757) := X"01010101";
        ram_buffer(75758) := X"01010101";
        ram_buffer(75759) := X"01010101";
        ram_buffer(75760) := X"01010101";
        ram_buffer(75761) := X"01010101";
        ram_buffer(75762) := X"10101010";
        ram_buffer(75763) := X"10104242";
        ram_buffer(75764) := X"42424242";
        ram_buffer(75765) := X"02020202";
        ram_buffer(75766) := X"02020202";
        ram_buffer(75767) := X"02020202";
        ram_buffer(75768) := X"02020202";
        ram_buffer(75769) := X"02020202";
        ram_buffer(75770) := X"10101010";
        ram_buffer(75771) := X"20000000";
        ram_buffer(75772) := X"00000000";
        ram_buffer(75773) := X"00000000";
        ram_buffer(75774) := X"00000000";
        ram_buffer(75775) := X"00000000";
        ram_buffer(75776) := X"00000000";
        ram_buffer(75777) := X"00000000";
        ram_buffer(75778) := X"00000000";
        ram_buffer(75779) := X"00000000";
        ram_buffer(75780) := X"00000000";
        ram_buffer(75781) := X"00000000";
        ram_buffer(75782) := X"00000000";
        ram_buffer(75783) := X"00000000";
        ram_buffer(75784) := X"00000000";
        ram_buffer(75785) := X"00000000";
        ram_buffer(75786) := X"00000000";
        ram_buffer(75787) := X"00000000";
        ram_buffer(75788) := X"00000000";
        ram_buffer(75789) := X"00000000";
        ram_buffer(75790) := X"00000000";
        ram_buffer(75791) := X"00000000";
        ram_buffer(75792) := X"00000000";
        ram_buffer(75793) := X"00000000";
        ram_buffer(75794) := X"00000000";
        ram_buffer(75795) := X"00000000";
        ram_buffer(75796) := X"00000000";
        ram_buffer(75797) := X"00000000";
        ram_buffer(75798) := X"00000000";
        ram_buffer(75799) := X"00000000";
        ram_buffer(75800) := X"00000000";
        ram_buffer(75801) := X"00000000";
        ram_buffer(75802) := X"00000000";
        ram_buffer(75803) := X"00000000";
        ram_buffer(75804) := X"43000000";
        ram_buffer(75805) := X"0A000000";
        ram_buffer(75806) := X"494E4600";
        ram_buffer(75807) := X"696E6600";
        ram_buffer(75808) := X"4E414E00";
        ram_buffer(75809) := X"6E616E00";
        ram_buffer(75810) := X"30313233";
        ram_buffer(75811) := X"34353637";
        ram_buffer(75812) := X"38396162";
        ram_buffer(75813) := X"63646566";
        ram_buffer(75814) := X"00000000";
        ram_buffer(75815) := X"286E756C";
        ram_buffer(75816) := X"6C290000";
        ram_buffer(75817) := X"30313233";
        ram_buffer(75818) := X"34353637";
        ram_buffer(75819) := X"38394142";
        ram_buffer(75820) := X"43444546";
        ram_buffer(75821) := X"00000000";
        ram_buffer(75822) := X"62756720";
        ram_buffer(75823) := X"696E2076";
        ram_buffer(75824) := X"66707269";
        ram_buffer(75825) := X"6E74663A";
        ram_buffer(75826) := X"20626164";
        ram_buffer(75827) := X"20626173";
        ram_buffer(75828) := X"65000000";
        ram_buffer(75829) := X"30000000";
        ram_buffer(75830) := X"100A19D8";
        ram_buffer(75831) := X"100A2E9C";
        ram_buffer(75832) := X"100A2E9C";
        ram_buffer(75833) := X"100A19F8";
        ram_buffer(75834) := X"100A2E9C";
        ram_buffer(75835) := X"100A2E9C";
        ram_buffer(75836) := X"100A2E9C";
        ram_buffer(75837) := X"100A1954";
        ram_buffer(75838) := X"100A2E9C";
        ram_buffer(75839) := X"100A2E9C";
        ram_buffer(75840) := X"100A1A04";
        ram_buffer(75841) := X"100A1A54";
        ram_buffer(75842) := X"100A2E9C";
        ram_buffer(75843) := X"100A1A48";
        ram_buffer(75844) := X"100A1A64";
        ram_buffer(75845) := X"100A2E9C";
        ram_buffer(75846) := X"100A1B28";
        ram_buffer(75847) := X"100A1B34";
        ram_buffer(75848) := X"100A1B34";
        ram_buffer(75849) := X"100A1B34";
        ram_buffer(75850) := X"100A1B34";
        ram_buffer(75851) := X"100A1B34";
        ram_buffer(75852) := X"100A1B34";
        ram_buffer(75853) := X"100A1B34";
        ram_buffer(75854) := X"100A1B34";
        ram_buffer(75855) := X"100A1B34";
        ram_buffer(75856) := X"100A2E9C";
        ram_buffer(75857) := X"100A2E9C";
        ram_buffer(75858) := X"100A2E9C";
        ram_buffer(75859) := X"100A2E9C";
        ram_buffer(75860) := X"100A2E9C";
        ram_buffer(75861) := X"100A2E9C";
        ram_buffer(75862) := X"100A2E9C";
        ram_buffer(75863) := X"100A1DC4";
        ram_buffer(75864) := X"100A2E9C";
        ram_buffer(75865) := X"100A1C00";
        ram_buffer(75866) := X"100A1C3C";
        ram_buffer(75867) := X"100A1DC4";
        ram_buffer(75868) := X"100A1DC4";
        ram_buffer(75869) := X"100A1DC4";
        ram_buffer(75870) := X"100A2E9C";
        ram_buffer(75871) := X"100A2E9C";
        ram_buffer(75872) := X"100A2E9C";
        ram_buffer(75873) := X"100A2E9C";
        ram_buffer(75874) := X"100A1B84";
        ram_buffer(75875) := X"100A2E9C";
        ram_buffer(75876) := X"100A2E9C";
        ram_buffer(75877) := X"100A2548";
        ram_buffer(75878) := X"100A2E9C";
        ram_buffer(75879) := X"100A2E9C";
        ram_buffer(75880) := X"100A2E9C";
        ram_buffer(75881) := X"100A26E0";
        ram_buffer(75882) := X"100A2E9C";
        ram_buffer(75883) := X"100A27B4";
        ram_buffer(75884) := X"100A2E9C";
        ram_buffer(75885) := X"100A2E9C";
        ram_buffer(75886) := X"100A2914";
        ram_buffer(75887) := X"100A2E9C";
        ram_buffer(75888) := X"100A2E9C";
        ram_buffer(75889) := X"100A2E9C";
        ram_buffer(75890) := X"100A2E9C";
        ram_buffer(75891) := X"100A2E9C";
        ram_buffer(75892) := X"100A2E9C";
        ram_buffer(75893) := X"100A2E9C";
        ram_buffer(75894) := X"100A2E9C";
        ram_buffer(75895) := X"100A1DC4";
        ram_buffer(75896) := X"100A2E9C";
        ram_buffer(75897) := X"100A1C00";
        ram_buffer(75898) := X"100A1C40";
        ram_buffer(75899) := X"100A1DC4";
        ram_buffer(75900) := X"100A1DC4";
        ram_buffer(75901) := X"100A1DC4";
        ram_buffer(75902) := X"100A1B90";
        ram_buffer(75903) := X"100A1C40";
        ram_buffer(75904) := X"100A1BF4";
        ram_buffer(75905) := X"100A2E9C";
        ram_buffer(75906) := X"100A1BBC";
        ram_buffer(75907) := X"100A2E9C";
        ram_buffer(75908) := X"100A2428";
        ram_buffer(75909) := X"100A254C";
        ram_buffer(75910) := X"100A268C";
        ram_buffer(75911) := X"100A1BE8";
        ram_buffer(75912) := X"100A2E9C";
        ram_buffer(75913) := X"100A26E0";
        ram_buffer(75914) := X"100A1910";
        ram_buffer(75915) := X"100A27B8";
        ram_buffer(75916) := X"100A2E9C";
        ram_buffer(75917) := X"100A2E9C";
        ram_buffer(75918) := X"100A2928";
        ram_buffer(75919) := X"100A2E9C";
        ram_buffer(75920) := X"100A1910";
        ram_buffer(75921) := X"20202020";
        ram_buffer(75922) := X"20202020";
        ram_buffer(75923) := X"20202020";
        ram_buffer(75924) := X"20202020";
        ram_buffer(75925) := X"30303030";
        ram_buffer(75926) := X"30303030";
        ram_buffer(75927) := X"30303030";
        ram_buffer(75928) := X"30303030";
        ram_buffer(75929) := X"65256C64";
        ram_buffer(75930) := X"00000000";
        ram_buffer(75931) := X"100A5744";
        ram_buffer(75932) := X"100A5750";
        ram_buffer(75933) := X"100A5750";
        ram_buffer(75934) := X"100A5750";
        ram_buffer(75935) := X"100A5750";
        ram_buffer(75936) := X"100A5750";
        ram_buffer(75937) := X"100A5750";
        ram_buffer(75938) := X"100A5750";
        ram_buffer(75939) := X"100A5750";
        ram_buffer(75940) := X"100A5750";
        ram_buffer(75941) := X"100A5750";
        ram_buffer(75942) := X"100A5750";
        ram_buffer(75943) := X"100A5750";
        ram_buffer(75944) := X"100A5750";
        ram_buffer(75945) := X"100A5750";
        ram_buffer(75946) := X"100A5750";
        ram_buffer(75947) := X"100A5750";
        ram_buffer(75948) := X"100A5750";
        ram_buffer(75949) := X"100A5750";
        ram_buffer(75950) := X"100A5750";
        ram_buffer(75951) := X"100A5750";
        ram_buffer(75952) := X"100A5750";
        ram_buffer(75953) := X"100A5750";
        ram_buffer(75954) := X"100A5750";
        ram_buffer(75955) := X"100A5750";
        ram_buffer(75956) := X"100A5750";
        ram_buffer(75957) := X"100A5750";
        ram_buffer(75958) := X"100A5750";
        ram_buffer(75959) := X"100A5750";
        ram_buffer(75960) := X"100A5750";
        ram_buffer(75961) := X"100A5750";
        ram_buffer(75962) := X"100A5750";
        ram_buffer(75963) := X"100A5750";
        ram_buffer(75964) := X"100A5750";
        ram_buffer(75965) := X"100A5750";
        ram_buffer(75966) := X"100A5750";
        ram_buffer(75967) := X"100A5750";
        ram_buffer(75968) := X"100A5348";
        ram_buffer(75969) := X"100A5750";
        ram_buffer(75970) := X"100A5750";
        ram_buffer(75971) := X"100A5750";
        ram_buffer(75972) := X"100A5750";
        ram_buffer(75973) := X"100A5414";
        ram_buffer(75974) := X"100A5750";
        ram_buffer(75975) := X"100A5750";
        ram_buffer(75976) := X"100A5750";
        ram_buffer(75977) := X"100A5750";
        ram_buffer(75978) := X"100A5750";
        ram_buffer(75979) := X"100A5490";
        ram_buffer(75980) := X"100A5490";
        ram_buffer(75981) := X"100A5490";
        ram_buffer(75982) := X"100A5490";
        ram_buffer(75983) := X"100A5490";
        ram_buffer(75984) := X"100A5490";
        ram_buffer(75985) := X"100A5490";
        ram_buffer(75986) := X"100A5490";
        ram_buffer(75987) := X"100A5490";
        ram_buffer(75988) := X"100A5490";
        ram_buffer(75989) := X"100A5750";
        ram_buffer(75990) := X"100A5750";
        ram_buffer(75991) := X"100A5750";
        ram_buffer(75992) := X"100A5750";
        ram_buffer(75993) := X"100A5750";
        ram_buffer(75994) := X"100A5750";
        ram_buffer(75995) := X"100A5750";
        ram_buffer(75996) := X"100A555C";
        ram_buffer(75997) := X"100A5750";
        ram_buffer(75998) := X"100A55A0";
        ram_buffer(75999) := X"100A54B4";
        ram_buffer(76000) := X"100A555C";
        ram_buffer(76001) := X"100A555C";
        ram_buffer(76002) := X"100A555C";
        ram_buffer(76003) := X"100A5750";
        ram_buffer(76004) := X"100A5750";
        ram_buffer(76005) := X"100A5750";
        ram_buffer(76006) := X"100A5750";
        ram_buffer(76007) := X"100A544C";
        ram_buffer(76008) := X"100A5750";
        ram_buffer(76009) := X"100A5750";
        ram_buffer(76010) := X"100A54F4";
        ram_buffer(76011) := X"100A5750";
        ram_buffer(76012) := X"100A5750";
        ram_buffer(76013) := X"100A5750";
        ram_buffer(76014) := X"100A5568";
        ram_buffer(76015) := X"100A5750";
        ram_buffer(76016) := X"100A5750";
        ram_buffer(76017) := X"100A5750";
        ram_buffer(76018) := X"100A5750";
        ram_buffer(76019) := X"100A5538";
        ram_buffer(76020) := X"100A5750";
        ram_buffer(76021) := X"100A5750";
        ram_buffer(76022) := X"100A5578";
        ram_buffer(76023) := X"100A5750";
        ram_buffer(76024) := X"100A5750";
        ram_buffer(76025) := X"100A5750";
        ram_buffer(76026) := X"100A5750";
        ram_buffer(76027) := X"100A5750";
        ram_buffer(76028) := X"100A555C";
        ram_buffer(76029) := X"100A5750";
        ram_buffer(76030) := X"100A55A4";
        ram_buffer(76031) := X"100A54B8";
        ram_buffer(76032) := X"100A555C";
        ram_buffer(76033) := X"100A555C";
        ram_buffer(76034) := X"100A555C";
        ram_buffer(76035) := X"100A5458";
        ram_buffer(76036) := X"100A54D8";
        ram_buffer(76037) := X"100A5484";
        ram_buffer(76038) := X"100A5750";
        ram_buffer(76039) := X"100A5420";
        ram_buffer(76040) := X"100A5750";
        ram_buffer(76041) := X"100A55D8";
        ram_buffer(76042) := X"100A54F8";
        ram_buffer(76043) := X"100A55B4";
        ram_buffer(76044) := X"100A5750";
        ram_buffer(76045) := X"100A5750";
        ram_buffer(76046) := X"100A556C";
        ram_buffer(76047) := X"100A5304";
        ram_buffer(76048) := X"100A5518";
        ram_buffer(76049) := X"100A5750";
        ram_buffer(76050) := X"100A5750";
        ram_buffer(76051) := X"100A5538";
        ram_buffer(76052) := X"100A5750";
        ram_buffer(76053) := X"100A5304";
        ram_buffer(76054) := X"100A5898";
        ram_buffer(76055) := X"100A5BC4";
        ram_buffer(76056) := X"100A5DCC";
        ram_buffer(76057) := X"100A623C";
        ram_buffer(76058) := X"100A6788";
        ram_buffer(76059) := X"100A63DC";
        ram_buffer(76060) := X"100A64D0";
        ram_buffer(76061) := X"100A63DC";
        ram_buffer(76062) := X"100A64D0";
        ram_buffer(76063) := X"100A64D0";
        ram_buffer(76064) := X"100A62B4";
        ram_buffer(76065) := X"100A633C";
        ram_buffer(76066) := X"100A633C";
        ram_buffer(76067) := X"100A633C";
        ram_buffer(76068) := X"100A633C";
        ram_buffer(76069) := X"100A633C";
        ram_buffer(76070) := X"100A633C";
        ram_buffer(76071) := X"100A633C";
        ram_buffer(76072) := X"100A6370";
        ram_buffer(76073) := X"100A6370";
        ram_buffer(76074) := X"100A64D0";
        ram_buffer(76075) := X"100A64D0";
        ram_buffer(76076) := X"100A64D0";
        ram_buffer(76077) := X"100A64D0";
        ram_buffer(76078) := X"100A64D0";
        ram_buffer(76079) := X"100A64D0";
        ram_buffer(76080) := X"100A64D0";
        ram_buffer(76081) := X"100A63B8";
        ram_buffer(76082) := X"100A63B8";
        ram_buffer(76083) := X"100A63B8";
        ram_buffer(76084) := X"100A63B8";
        ram_buffer(76085) := X"100A63B8";
        ram_buffer(76086) := X"100A63B8";
        ram_buffer(76087) := X"100A64D0";
        ram_buffer(76088) := X"100A64D0";
        ram_buffer(76089) := X"100A64D0";
        ram_buffer(76090) := X"100A64D0";
        ram_buffer(76091) := X"100A64D0";
        ram_buffer(76092) := X"100A64D0";
        ram_buffer(76093) := X"100A64D0";
        ram_buffer(76094) := X"100A64D0";
        ram_buffer(76095) := X"100A64D0";
        ram_buffer(76096) := X"100A64D0";
        ram_buffer(76097) := X"100A64D0";
        ram_buffer(76098) := X"100A64D0";
        ram_buffer(76099) := X"100A64D0";
        ram_buffer(76100) := X"100A64D0";
        ram_buffer(76101) := X"100A64D0";
        ram_buffer(76102) := X"100A64D0";
        ram_buffer(76103) := X"100A64D0";
        ram_buffer(76104) := X"100A63F8";
        ram_buffer(76105) := X"100A64D0";
        ram_buffer(76106) := X"100A64D0";
        ram_buffer(76107) := X"100A64D0";
        ram_buffer(76108) := X"100A64D0";
        ram_buffer(76109) := X"100A64D0";
        ram_buffer(76110) := X"100A64D0";
        ram_buffer(76111) := X"100A64D0";
        ram_buffer(76112) := X"100A64D0";
        ram_buffer(76113) := X"100A63B8";
        ram_buffer(76114) := X"100A63B8";
        ram_buffer(76115) := X"100A63B8";
        ram_buffer(76116) := X"100A63B8";
        ram_buffer(76117) := X"100A63B8";
        ram_buffer(76118) := X"100A63B8";
        ram_buffer(76119) := X"100A64D0";
        ram_buffer(76120) := X"100A64D0";
        ram_buffer(76121) := X"100A64D0";
        ram_buffer(76122) := X"100A64D0";
        ram_buffer(76123) := X"100A64D0";
        ram_buffer(76124) := X"100A64D0";
        ram_buffer(76125) := X"100A64D0";
        ram_buffer(76126) := X"100A64D0";
        ram_buffer(76127) := X"100A64D0";
        ram_buffer(76128) := X"100A64D0";
        ram_buffer(76129) := X"100A64D0";
        ram_buffer(76130) := X"100A64D0";
        ram_buffer(76131) := X"100A64D0";
        ram_buffer(76132) := X"100A64D0";
        ram_buffer(76133) := X"100A64D0";
        ram_buffer(76134) := X"100A64D0";
        ram_buffer(76135) := X"100A64D0";
        ram_buffer(76136) := X"100A63F8";
        ram_buffer(76137) := X"100A68A4";
        ram_buffer(76138) := X"100A6AD8";
        ram_buffer(76139) := X"100A68A4";
        ram_buffer(76140) := X"100A6AD8";
        ram_buffer(76141) := X"100A6AD8";
        ram_buffer(76142) := X"100A682C";
        ram_buffer(76143) := X"100A687C";
        ram_buffer(76144) := X"100A687C";
        ram_buffer(76145) := X"100A687C";
        ram_buffer(76146) := X"100A687C";
        ram_buffer(76147) := X"100A687C";
        ram_buffer(76148) := X"100A687C";
        ram_buffer(76149) := X"100A687C";
        ram_buffer(76150) := X"100A687C";
        ram_buffer(76151) := X"100A687C";
        ram_buffer(76152) := X"100A6AD8";
        ram_buffer(76153) := X"100A6AD8";
        ram_buffer(76154) := X"100A6AD8";
        ram_buffer(76155) := X"100A6AD8";
        ram_buffer(76156) := X"100A6AD8";
        ram_buffer(76157) := X"100A6AD8";
        ram_buffer(76158) := X"100A6AD8";
        ram_buffer(76159) := X"100A6968";
        ram_buffer(76160) := X"100A6AD8";
        ram_buffer(76161) := X"100A6AD8";
        ram_buffer(76162) := X"100A6AD8";
        ram_buffer(76163) := X"100A6A70";
        ram_buffer(76164) := X"100A6A10";
        ram_buffer(76165) := X"100A6AD8";
        ram_buffer(76166) := X"100A6AD8";
        ram_buffer(76167) := X"100A6988";
        ram_buffer(76168) := X"100A6AD8";
        ram_buffer(76169) := X"100A6AD8";
        ram_buffer(76170) := X"100A6AD8";
        ram_buffer(76171) := X"100A6AD8";
        ram_buffer(76172) := X"100A68C0";
        ram_buffer(76173) := X"100A6AD8";
        ram_buffer(76174) := X"100A6AD8";
        ram_buffer(76175) := X"100A6AD8";
        ram_buffer(76176) := X"100A6AD8";
        ram_buffer(76177) := X"100A6AD8";
        ram_buffer(76178) := X"100A6A30";
        ram_buffer(76179) := X"100A6AD8";
        ram_buffer(76180) := X"100A6AD8";
        ram_buffer(76181) := X"100A6AD8";
        ram_buffer(76182) := X"100A6AD8";
        ram_buffer(76183) := X"100A6A50";
        ram_buffer(76184) := X"100A6AD8";
        ram_buffer(76185) := X"100A6AD8";
        ram_buffer(76186) := X"100A6AD8";
        ram_buffer(76187) := X"100A6AD8";
        ram_buffer(76188) := X"100A6AD8";
        ram_buffer(76189) := X"100A6AD8";
        ram_buffer(76190) := X"100A6AD8";
        ram_buffer(76191) := X"100A6968";
        ram_buffer(76192) := X"100A6AD8";
        ram_buffer(76193) := X"100A6AD8";
        ram_buffer(76194) := X"100A6AD8";
        ram_buffer(76195) := X"100A6A70";
        ram_buffer(76196) := X"100A6A10";
        ram_buffer(76197) := X"100A6AD8";
        ram_buffer(76198) := X"100A6AD8";
        ram_buffer(76199) := X"100A6988";
        ram_buffer(76200) := X"100A6AD8";
        ram_buffer(76201) := X"100A6AD8";
        ram_buffer(76202) := X"100A6AD8";
        ram_buffer(76203) := X"100A6AD8";
        ram_buffer(76204) := X"100A68C0";
        ram_buffer(76205) := X"100A6AD8";
        ram_buffer(76206) := X"100A6AD8";
        ram_buffer(76207) := X"100A6AD8";
        ram_buffer(76208) := X"100A6AD8";
        ram_buffer(76209) := X"100A6AD8";
        ram_buffer(76210) := X"100A6A30";
        ram_buffer(76211) := X"100A6AD8";
        ram_buffer(76212) := X"100A6AD8";
        ram_buffer(76213) := X"100A6AD8";
        ram_buffer(76214) := X"100A6AD8";
        ram_buffer(76215) := X"100A6A50";
        ram_buffer(76216) := X"000A0001";
        ram_buffer(76217) := X"00020003";
        ram_buffer(76218) := X"00040005";
        ram_buffer(76219) := X"00060007";
        ram_buffer(76220) := X"00080009";
        ram_buffer(76221) := X"000A000B";
        ram_buffer(76222) := X"000C000D";
        ram_buffer(76223) := X"000E000F";
        ram_buffer(76224) := X"00100000";
        ram_buffer(76225) := X"494E4600";
        ram_buffer(76226) := X"696E6600";
        ram_buffer(76227) := X"4E414E00";
        ram_buffer(76228) := X"6E616E00";
        ram_buffer(76229) := X"30313233";
        ram_buffer(76230) := X"34353637";
        ram_buffer(76231) := X"38396162";
        ram_buffer(76232) := X"63646566";
        ram_buffer(76233) := X"00000000";
        ram_buffer(76234) := X"286E756C";
        ram_buffer(76235) := X"6C290000";
        ram_buffer(76236) := X"30313233";
        ram_buffer(76237) := X"34353637";
        ram_buffer(76238) := X"38394142";
        ram_buffer(76239) := X"43444546";
        ram_buffer(76240) := X"00000000";
        ram_buffer(76241) := X"62756720";
        ram_buffer(76242) := X"696E2076";
        ram_buffer(76243) := X"66707269";
        ram_buffer(76244) := X"6E74663A";
        ram_buffer(76245) := X"20626164";
        ram_buffer(76246) := X"20626173";
        ram_buffer(76247) := X"65000000";
        ram_buffer(76248) := X"30000000";
        ram_buffer(76249) := X"100A7BBC";
        ram_buffer(76250) := X"100A9080";
        ram_buffer(76251) := X"100A9080";
        ram_buffer(76252) := X"100A7BDC";
        ram_buffer(76253) := X"100A9080";
        ram_buffer(76254) := X"100A9080";
        ram_buffer(76255) := X"100A9080";
        ram_buffer(76256) := X"100A7B38";
        ram_buffer(76257) := X"100A9080";
        ram_buffer(76258) := X"100A9080";
        ram_buffer(76259) := X"100A7BE8";
        ram_buffer(76260) := X"100A7C38";
        ram_buffer(76261) := X"100A9080";
        ram_buffer(76262) := X"100A7C2C";
        ram_buffer(76263) := X"100A7C48";
        ram_buffer(76264) := X"100A9080";
        ram_buffer(76265) := X"100A7D0C";
        ram_buffer(76266) := X"100A7D18";
        ram_buffer(76267) := X"100A7D18";
        ram_buffer(76268) := X"100A7D18";
        ram_buffer(76269) := X"100A7D18";
        ram_buffer(76270) := X"100A7D18";
        ram_buffer(76271) := X"100A7D18";
        ram_buffer(76272) := X"100A7D18";
        ram_buffer(76273) := X"100A7D18";
        ram_buffer(76274) := X"100A7D18";
        ram_buffer(76275) := X"100A9080";
        ram_buffer(76276) := X"100A9080";
        ram_buffer(76277) := X"100A9080";
        ram_buffer(76278) := X"100A9080";
        ram_buffer(76279) := X"100A9080";
        ram_buffer(76280) := X"100A9080";
        ram_buffer(76281) := X"100A9080";
        ram_buffer(76282) := X"100A7FA8";
        ram_buffer(76283) := X"100A9080";
        ram_buffer(76284) := X"100A7DE4";
        ram_buffer(76285) := X"100A7E20";
        ram_buffer(76286) := X"100A7FA8";
        ram_buffer(76287) := X"100A7FA8";
        ram_buffer(76288) := X"100A7FA8";
        ram_buffer(76289) := X"100A9080";
        ram_buffer(76290) := X"100A9080";
        ram_buffer(76291) := X"100A9080";
        ram_buffer(76292) := X"100A9080";
        ram_buffer(76293) := X"100A7D68";
        ram_buffer(76294) := X"100A9080";
        ram_buffer(76295) := X"100A9080";
        ram_buffer(76296) := X"100A872C";
        ram_buffer(76297) := X"100A9080";
        ram_buffer(76298) := X"100A9080";
        ram_buffer(76299) := X"100A9080";
        ram_buffer(76300) := X"100A88C4";
        ram_buffer(76301) := X"100A9080";
        ram_buffer(76302) := X"100A8998";
        ram_buffer(76303) := X"100A9080";
        ram_buffer(76304) := X"100A9080";
        ram_buffer(76305) := X"100A8AF8";
        ram_buffer(76306) := X"100A9080";
        ram_buffer(76307) := X"100A9080";
        ram_buffer(76308) := X"100A9080";
        ram_buffer(76309) := X"100A9080";
        ram_buffer(76310) := X"100A9080";
        ram_buffer(76311) := X"100A9080";
        ram_buffer(76312) := X"100A9080";
        ram_buffer(76313) := X"100A9080";
        ram_buffer(76314) := X"100A7FA8";
        ram_buffer(76315) := X"100A9080";
        ram_buffer(76316) := X"100A7DE4";
        ram_buffer(76317) := X"100A7E24";
        ram_buffer(76318) := X"100A7FA8";
        ram_buffer(76319) := X"100A7FA8";
        ram_buffer(76320) := X"100A7FA8";
        ram_buffer(76321) := X"100A7D74";
        ram_buffer(76322) := X"100A7E24";
        ram_buffer(76323) := X"100A7DD8";
        ram_buffer(76324) := X"100A9080";
        ram_buffer(76325) := X"100A7DA0";
        ram_buffer(76326) := X"100A9080";
        ram_buffer(76327) := X"100A860C";
        ram_buffer(76328) := X"100A8730";
        ram_buffer(76329) := X"100A8870";
        ram_buffer(76330) := X"100A7DCC";
        ram_buffer(76331) := X"100A9080";
        ram_buffer(76332) := X"100A88C4";
        ram_buffer(76333) := X"100A7AF4";
        ram_buffer(76334) := X"100A899C";
        ram_buffer(76335) := X"100A9080";
        ram_buffer(76336) := X"100A9080";
        ram_buffer(76337) := X"100A8B0C";
        ram_buffer(76338) := X"100A9080";
        ram_buffer(76339) := X"100A7AF4";
        ram_buffer(76340) := X"20202020";
        ram_buffer(76341) := X"20202020";
        ram_buffer(76342) := X"20202020";
        ram_buffer(76343) := X"20202020";
        ram_buffer(76344) := X"30303030";
        ram_buffer(76345) := X"30303030";
        ram_buffer(76346) := X"30303030";
        ram_buffer(76347) := X"30303030";
        ram_buffer(76348) := X"496E6669";
        ram_buffer(76349) := X"6E697479";
        ram_buffer(76350) := X"00000000";
        ram_buffer(76351) := X"4E614E00";
        ram_buffer(76352) := X"30000000";
        ram_buffer(76353) := X"100AC534";
        ram_buffer(76354) := X"100AC534";
        ram_buffer(76355) := X"100AC548";
        ram_buffer(76356) := X"100AC590";
        ram_buffer(76357) := X"100AC54C";
        ram_buffer(76358) := X"100AC594";
        ram_buffer(76359) := X"2E000000";
        ram_buffer(76360) := X"00000000";
        ram_buffer(76361) := X"504F5349";
        ram_buffer(76362) := X"58000000";
        ram_buffer(76363) := X"43000000";
        ram_buffer(76364) := X"00000000";
        ram_buffer(76365) := X"00000000";
        ram_buffer(76366) := X"3FF00000";
        ram_buffer(76367) := X"00000000";
        ram_buffer(76368) := X"40240000";
        ram_buffer(76369) := X"00000000";
        ram_buffer(76370) := X"40590000";
        ram_buffer(76371) := X"00000000";
        ram_buffer(76372) := X"408F4000";
        ram_buffer(76373) := X"00000000";
        ram_buffer(76374) := X"40C38800";
        ram_buffer(76375) := X"00000000";
        ram_buffer(76376) := X"40F86A00";
        ram_buffer(76377) := X"00000000";
        ram_buffer(76378) := X"412E8480";
        ram_buffer(76379) := X"00000000";
        ram_buffer(76380) := X"416312D0";
        ram_buffer(76381) := X"00000000";
        ram_buffer(76382) := X"4197D784";
        ram_buffer(76383) := X"00000000";
        ram_buffer(76384) := X"41CDCD65";
        ram_buffer(76385) := X"00000000";
        ram_buffer(76386) := X"4202A05F";
        ram_buffer(76387) := X"20000000";
        ram_buffer(76388) := X"42374876";
        ram_buffer(76389) := X"E8000000";
        ram_buffer(76390) := X"426D1A94";
        ram_buffer(76391) := X"A2000000";
        ram_buffer(76392) := X"42A2309C";
        ram_buffer(76393) := X"E5400000";
        ram_buffer(76394) := X"42D6BCC4";
        ram_buffer(76395) := X"1E900000";
        ram_buffer(76396) := X"430C6BF5";
        ram_buffer(76397) := X"26340000";
        ram_buffer(76398) := X"4341C379";
        ram_buffer(76399) := X"37E08000";
        ram_buffer(76400) := X"43763457";
        ram_buffer(76401) := X"85D8A000";
        ram_buffer(76402) := X"43ABC16D";
        ram_buffer(76403) := X"674EC800";
        ram_buffer(76404) := X"43E158E4";
        ram_buffer(76405) := X"60913D00";
        ram_buffer(76406) := X"4415AF1D";
        ram_buffer(76407) := X"78B58C40";
        ram_buffer(76408) := X"444B1AE4";
        ram_buffer(76409) := X"D6E2EF50";
        ram_buffer(76410) := X"4480F0CF";
        ram_buffer(76411) := X"064DD592";
        ram_buffer(76412) := X"44B52D02";
        ram_buffer(76413) := X"C7E14AF6";
        ram_buffer(76414) := X"44EA7843";
        ram_buffer(76415) := X"79D99DB4";
        ram_buffer(76416) := X"4341C379";
        ram_buffer(76417) := X"37E08000";
        ram_buffer(76418) := X"4693B8B5";
        ram_buffer(76419) := X"B5056E17";
        ram_buffer(76420) := X"4D384F03";
        ram_buffer(76421) := X"E93FF9F5";
        ram_buffer(76422) := X"5A827748";
        ram_buffer(76423) := X"F9301D32";
        ram_buffer(76424) := X"75154FDD";
        ram_buffer(76425) := X"7F73BF3C";
        ram_buffer(76426) := X"3C9CD2B2";
        ram_buffer(76427) := X"97D889BC";
        ram_buffer(76428) := X"3949F623";
        ram_buffer(76429) := X"D5A8A733";
        ram_buffer(76430) := X"32A50FFD";
        ram_buffer(76431) := X"44F4A73D";
        ram_buffer(76432) := X"255BBA08";
        ram_buffer(76433) := X"CF8C979D";
        ram_buffer(76434) := X"0AC80628";
        ram_buffer(76435) := X"64AC6F43";
        ram_buffer(76436) := X"00000005";
        ram_buffer(76437) := X"00000019";
        ram_buffer(76438) := X"0000007D";
        ram_buffer(76439) := X"00000000";
        ram_buffer(76440) := X"3C9CD2B2";
        ram_buffer(76441) := X"97D889BC";
        ram_buffer(76442) := X"3949F623";
        ram_buffer(76443) := X"D5A8A733";
        ram_buffer(76444) := X"32A50FFD";
        ram_buffer(76445) := X"44F4A73D";
        ram_buffer(76446) := X"255BBA08";
        ram_buffer(76447) := X"CF8C979D";
        ram_buffer(76448) := X"11680628";
        ram_buffer(76449) := X"64AC6F43";
        ram_buffer(76450) := X"100B3A08";
        ram_buffer(76451) := X"100B3A70";
        ram_buffer(76452) := X"100B3A30";
        ram_buffer(76453) := X"100B3AD4";
        ram_buffer(76454) := X"100B3AF8";
        ram_buffer(76455) := X"100B3A70";
        ram_buffer(76456) := X"100B3A08";
        ram_buffer(76457) := X"6E660000";
        ram_buffer(76458) := X"696E6974";
        ram_buffer(76459) := X"79000000";
        ram_buffer(76460) := X"616E0000";
        ram_buffer(76461) := X"100B4794";
        ram_buffer(76462) := X"100B3DA0";
        ram_buffer(76463) := X"100B3DA0";
        ram_buffer(76464) := X"100B3DA0";
        ram_buffer(76465) := X"100B3DA0";
        ram_buffer(76466) := X"100B3DA0";
        ram_buffer(76467) := X"100B3DA0";
        ram_buffer(76468) := X"100B3DA0";
        ram_buffer(76469) := X"100B3DA0";
        ram_buffer(76470) := X"100B3D88";
        ram_buffer(76471) := X"100B3D88";
        ram_buffer(76472) := X"100B3D88";
        ram_buffer(76473) := X"100B3D88";
        ram_buffer(76474) := X"100B3D88";
        ram_buffer(76475) := X"100B3DA0";
        ram_buffer(76476) := X"100B3DA0";
        ram_buffer(76477) := X"100B3DA0";
        ram_buffer(76478) := X"100B3DA0";
        ram_buffer(76479) := X"100B3DA0";
        ram_buffer(76480) := X"100B3DA0";
        ram_buffer(76481) := X"100B3DA0";
        ram_buffer(76482) := X"100B3DA0";
        ram_buffer(76483) := X"100B3DA0";
        ram_buffer(76484) := X"100B3DA0";
        ram_buffer(76485) := X"100B3DA0";
        ram_buffer(76486) := X"100B3DA0";
        ram_buffer(76487) := X"100B3DA0";
        ram_buffer(76488) := X"100B3DA0";
        ram_buffer(76489) := X"100B3DA0";
        ram_buffer(76490) := X"100B3DA0";
        ram_buffer(76491) := X"100B3DA0";
        ram_buffer(76492) := X"100B3DA0";
        ram_buffer(76493) := X"100B3D88";
        ram_buffer(76494) := X"100B3DA0";
        ram_buffer(76495) := X"100B3DA0";
        ram_buffer(76496) := X"100B3DA0";
        ram_buffer(76497) := X"100B3DA0";
        ram_buffer(76498) := X"100B3DA0";
        ram_buffer(76499) := X"100B3DA0";
        ram_buffer(76500) := X"100B3DA0";
        ram_buffer(76501) := X"100B3DA0";
        ram_buffer(76502) := X"100B3DA0";
        ram_buffer(76503) := X"100B3DA0";
        ram_buffer(76504) := X"100B3D58";
        ram_buffer(76505) := X"100B3DA0";
        ram_buffer(76506) := X"100B3D50";
        ram_buffer(76507) := X"00000035";
        ram_buffer(76508) := X"FFFFFBCE";
        ram_buffer(76509) := X"000003CB";
        ram_buffer(76510) := X"00000001";
        ram_buffer(76511) := X"00000000";
        ram_buffer(76512) := X"00000034";
        ram_buffer(76513) := X"FFFFFBCE";
        ram_buffer(76514) := X"000003CB";
        ram_buffer(76515) := X"00000001";
        ram_buffer(76516) := X"00000000";
        ram_buffer(76517) := X"00000000";
        ram_buffer(76518) := X"30313233";
        ram_buffer(76519) := X"34353637";
        ram_buffer(76520) := X"38396162";
        ram_buffer(76521) := X"63646566";
        ram_buffer(76522) := X"00000000";
        ram_buffer(76523) := X"286E756C";
        ram_buffer(76524) := X"6C290000";
        ram_buffer(76525) := X"30313233";
        ram_buffer(76526) := X"34353637";
        ram_buffer(76527) := X"38394142";
        ram_buffer(76528) := X"43444546";
        ram_buffer(76529) := X"00000000";
        ram_buffer(76530) := X"62756720";
        ram_buffer(76531) := X"696E2076";
        ram_buffer(76532) := X"66707269";
        ram_buffer(76533) := X"6E74663A";
        ram_buffer(76534) := X"20626164";
        ram_buffer(76535) := X"20626173";
        ram_buffer(76536) := X"65000000";
        ram_buffer(76537) := X"100B7958";
        ram_buffer(76538) := X"100B87AC";
        ram_buffer(76539) := X"100B87AC";
        ram_buffer(76540) := X"100B7978";
        ram_buffer(76541) := X"100B87AC";
        ram_buffer(76542) := X"100B87AC";
        ram_buffer(76543) := X"100B87AC";
        ram_buffer(76544) := X"100B78D4";
        ram_buffer(76545) := X"100B87AC";
        ram_buffer(76546) := X"100B87AC";
        ram_buffer(76547) := X"100B7984";
        ram_buffer(76548) := X"100B79D4";
        ram_buffer(76549) := X"100B87AC";
        ram_buffer(76550) := X"100B79C8";
        ram_buffer(76551) := X"100B79E4";
        ram_buffer(76552) := X"100B87AC";
        ram_buffer(76553) := X"100B7AA8";
        ram_buffer(76554) := X"100B7AB4";
        ram_buffer(76555) := X"100B7AB4";
        ram_buffer(76556) := X"100B7AB4";
        ram_buffer(76557) := X"100B7AB4";
        ram_buffer(76558) := X"100B7AB4";
        ram_buffer(76559) := X"100B7AB4";
        ram_buffer(76560) := X"100B7AB4";
        ram_buffer(76561) := X"100B7AB4";
        ram_buffer(76562) := X"100B7AB4";
        ram_buffer(76563) := X"100B87AC";
        ram_buffer(76564) := X"100B87AC";
        ram_buffer(76565) := X"100B87AC";
        ram_buffer(76566) := X"100B87AC";
        ram_buffer(76567) := X"100B87AC";
        ram_buffer(76568) := X"100B87AC";
        ram_buffer(76569) := X"100B87AC";
        ram_buffer(76570) := X"100B87AC";
        ram_buffer(76571) := X"100B87AC";
        ram_buffer(76572) := X"100B7B74";
        ram_buffer(76573) := X"100B7BB0";
        ram_buffer(76574) := X"100B87AC";
        ram_buffer(76575) := X"100B87AC";
        ram_buffer(76576) := X"100B87AC";
        ram_buffer(76577) := X"100B87AC";
        ram_buffer(76578) := X"100B87AC";
        ram_buffer(76579) := X"100B87AC";
        ram_buffer(76580) := X"100B87AC";
        ram_buffer(76581) := X"100B87AC";
        ram_buffer(76582) := X"100B87AC";
        ram_buffer(76583) := X"100B87AC";
        ram_buffer(76584) := X"100B7E58";
        ram_buffer(76585) := X"100B87AC";
        ram_buffer(76586) := X"100B87AC";
        ram_buffer(76587) := X"100B87AC";
        ram_buffer(76588) := X"100B7FF0";
        ram_buffer(76589) := X"100B87AC";
        ram_buffer(76590) := X"100B80C4";
        ram_buffer(76591) := X"100B87AC";
        ram_buffer(76592) := X"100B87AC";
        ram_buffer(76593) := X"100B8224";
        ram_buffer(76594) := X"100B87AC";
        ram_buffer(76595) := X"100B87AC";
        ram_buffer(76596) := X"100B87AC";
        ram_buffer(76597) := X"100B87AC";
        ram_buffer(76598) := X"100B87AC";
        ram_buffer(76599) := X"100B87AC";
        ram_buffer(76600) := X"100B87AC";
        ram_buffer(76601) := X"100B87AC";
        ram_buffer(76602) := X"100B87AC";
        ram_buffer(76603) := X"100B87AC";
        ram_buffer(76604) := X"100B7B74";
        ram_buffer(76605) := X"100B7BB4";
        ram_buffer(76606) := X"100B87AC";
        ram_buffer(76607) := X"100B87AC";
        ram_buffer(76608) := X"100B87AC";
        ram_buffer(76609) := X"100B7B04";
        ram_buffer(76610) := X"100B7BB4";
        ram_buffer(76611) := X"100B7B68";
        ram_buffer(76612) := X"100B87AC";
        ram_buffer(76613) := X"100B7B30";
        ram_buffer(76614) := X"100B87AC";
        ram_buffer(76615) := X"100B7D38";
        ram_buffer(76616) := X"100B7E5C";
        ram_buffer(76617) := X"100B7F9C";
        ram_buffer(76618) := X"100B7B5C";
        ram_buffer(76619) := X"100B87AC";
        ram_buffer(76620) := X"100B7FF0";
        ram_buffer(76621) := X"100B7890";
        ram_buffer(76622) := X"100B80C8";
        ram_buffer(76623) := X"100B87AC";
        ram_buffer(76624) := X"100B87AC";
        ram_buffer(76625) := X"100B8238";
        ram_buffer(76626) := X"100B87AC";
        ram_buffer(76627) := X"100B7890";
        ram_buffer(76628) := X"20202020";
        ram_buffer(76629) := X"20202020";
        ram_buffer(76630) := X"20202020";
        ram_buffer(76631) := X"20202020";
        ram_buffer(76632) := X"30303030";
        ram_buffer(76633) := X"30303030";
        ram_buffer(76634) := X"30303030";
        ram_buffer(76635) := X"30303030";
        ram_buffer(76636) := X"100B9A48";
        ram_buffer(76637) := X"100B9A54";
        ram_buffer(76638) := X"100B9A54";
        ram_buffer(76639) := X"100B9A54";
        ram_buffer(76640) := X"100B9A54";
        ram_buffer(76641) := X"100B9A54";
        ram_buffer(76642) := X"100B9A54";
        ram_buffer(76643) := X"100B9A54";
        ram_buffer(76644) := X"100B9A54";
        ram_buffer(76645) := X"100B9A54";
        ram_buffer(76646) := X"100B9A54";
        ram_buffer(76647) := X"100B9A54";
        ram_buffer(76648) := X"100B9A54";
        ram_buffer(76649) := X"100B9A54";
        ram_buffer(76650) := X"100B9A54";
        ram_buffer(76651) := X"100B9A54";
        ram_buffer(76652) := X"100B9A54";
        ram_buffer(76653) := X"100B9A54";
        ram_buffer(76654) := X"100B9A54";
        ram_buffer(76655) := X"100B9A54";
        ram_buffer(76656) := X"100B9A54";
        ram_buffer(76657) := X"100B9A54";
        ram_buffer(76658) := X"100B9A54";
        ram_buffer(76659) := X"100B9A54";
        ram_buffer(76660) := X"100B9A54";
        ram_buffer(76661) := X"100B9A54";
        ram_buffer(76662) := X"100B9A54";
        ram_buffer(76663) := X"100B9A54";
        ram_buffer(76664) := X"100B9A54";
        ram_buffer(76665) := X"100B9A54";
        ram_buffer(76666) := X"100B9A54";
        ram_buffer(76667) := X"100B9A54";
        ram_buffer(76668) := X"100B9A54";
        ram_buffer(76669) := X"100B9A54";
        ram_buffer(76670) := X"100B9A54";
        ram_buffer(76671) := X"100B9A54";
        ram_buffer(76672) := X"100B9A54";
        ram_buffer(76673) := X"100B9658";
        ram_buffer(76674) := X"100B9A54";
        ram_buffer(76675) := X"100B9A54";
        ram_buffer(76676) := X"100B9A54";
        ram_buffer(76677) := X"100B9A54";
        ram_buffer(76678) := X"100B9724";
        ram_buffer(76679) := X"100B9A54";
        ram_buffer(76680) := X"100B9A54";
        ram_buffer(76681) := X"100B9A54";
        ram_buffer(76682) := X"100B9A54";
        ram_buffer(76683) := X"100B9A54";
        ram_buffer(76684) := X"100B97A0";
        ram_buffer(76685) := X"100B97A0";
        ram_buffer(76686) := X"100B97A0";
        ram_buffer(76687) := X"100B97A0";
        ram_buffer(76688) := X"100B97A0";
        ram_buffer(76689) := X"100B97A0";
        ram_buffer(76690) := X"100B97A0";
        ram_buffer(76691) := X"100B97A0";
        ram_buffer(76692) := X"100B97A0";
        ram_buffer(76693) := X"100B97A0";
        ram_buffer(76694) := X"100B9A54";
        ram_buffer(76695) := X"100B9A54";
        ram_buffer(76696) := X"100B9A54";
        ram_buffer(76697) := X"100B9A54";
        ram_buffer(76698) := X"100B9A54";
        ram_buffer(76699) := X"100B9A54";
        ram_buffer(76700) := X"100B9A54";
        ram_buffer(76701) := X"100B9A54";
        ram_buffer(76702) := X"100B9A54";
        ram_buffer(76703) := X"100B98A4";
        ram_buffer(76704) := X"100B97C4";
        ram_buffer(76705) := X"100B9A54";
        ram_buffer(76706) := X"100B9A54";
        ram_buffer(76707) := X"100B9A54";
        ram_buffer(76708) := X"100B9A54";
        ram_buffer(76709) := X"100B9A54";
        ram_buffer(76710) := X"100B9A54";
        ram_buffer(76711) := X"100B9A54";
        ram_buffer(76712) := X"100B975C";
        ram_buffer(76713) := X"100B9A54";
        ram_buffer(76714) := X"100B9A54";
        ram_buffer(76715) := X"100B9804";
        ram_buffer(76716) := X"100B9A54";
        ram_buffer(76717) := X"100B9A54";
        ram_buffer(76718) := X"100B9A54";
        ram_buffer(76719) := X"100B986C";
        ram_buffer(76720) := X"100B9A54";
        ram_buffer(76721) := X"100B9A54";
        ram_buffer(76722) := X"100B9A54";
        ram_buffer(76723) := X"100B9A54";
        ram_buffer(76724) := X"100B9848";
        ram_buffer(76725) := X"100B9A54";
        ram_buffer(76726) := X"100B9A54";
        ram_buffer(76727) := X"100B987C";
        ram_buffer(76728) := X"100B9A54";
        ram_buffer(76729) := X"100B9A54";
        ram_buffer(76730) := X"100B9A54";
        ram_buffer(76731) := X"100B9A54";
        ram_buffer(76732) := X"100B9A54";
        ram_buffer(76733) := X"100B9A54";
        ram_buffer(76734) := X"100B9A54";
        ram_buffer(76735) := X"100B98A8";
        ram_buffer(76736) := X"100B97C8";
        ram_buffer(76737) := X"100B9A54";
        ram_buffer(76738) := X"100B9A54";
        ram_buffer(76739) := X"100B9A54";
        ram_buffer(76740) := X"100B9768";
        ram_buffer(76741) := X"100B97E8";
        ram_buffer(76742) := X"100B9794";
        ram_buffer(76743) := X"100B9A54";
        ram_buffer(76744) := X"100B9730";
        ram_buffer(76745) := X"100B9A54";
        ram_buffer(76746) := X"100B98DC";
        ram_buffer(76747) := X"100B9808";
        ram_buffer(76748) := X"100B98B8";
        ram_buffer(76749) := X"100B9A54";
        ram_buffer(76750) := X"100B9A54";
        ram_buffer(76751) := X"100B9870";
        ram_buffer(76752) := X"100B9614";
        ram_buffer(76753) := X"100B9828";
        ram_buffer(76754) := X"100B9A54";
        ram_buffer(76755) := X"100B9A54";
        ram_buffer(76756) := X"100B9848";
        ram_buffer(76757) := X"100B9A54";
        ram_buffer(76758) := X"100B9614";
        ram_buffer(76759) := X"100BA6FC";
        ram_buffer(76760) := X"100BA7F0";
        ram_buffer(76761) := X"100BA6FC";
        ram_buffer(76762) := X"100BA7F0";
        ram_buffer(76763) := X"100BA7F0";
        ram_buffer(76764) := X"100BA5D4";
        ram_buffer(76765) := X"100BA65C";
        ram_buffer(76766) := X"100BA65C";
        ram_buffer(76767) := X"100BA65C";
        ram_buffer(76768) := X"100BA65C";
        ram_buffer(76769) := X"100BA65C";
        ram_buffer(76770) := X"100BA65C";
        ram_buffer(76771) := X"100BA65C";
        ram_buffer(76772) := X"100BA690";
        ram_buffer(76773) := X"100BA690";
        ram_buffer(76774) := X"100BA7F0";
        ram_buffer(76775) := X"100BA7F0";
        ram_buffer(76776) := X"100BA7F0";
        ram_buffer(76777) := X"100BA7F0";
        ram_buffer(76778) := X"100BA7F0";
        ram_buffer(76779) := X"100BA7F0";
        ram_buffer(76780) := X"100BA7F0";
        ram_buffer(76781) := X"100BA6D8";
        ram_buffer(76782) := X"100BA6D8";
        ram_buffer(76783) := X"100BA6D8";
        ram_buffer(76784) := X"100BA6D8";
        ram_buffer(76785) := X"100BA6D8";
        ram_buffer(76786) := X"100BA6D8";
        ram_buffer(76787) := X"100BA7F0";
        ram_buffer(76788) := X"100BA7F0";
        ram_buffer(76789) := X"100BA7F0";
        ram_buffer(76790) := X"100BA7F0";
        ram_buffer(76791) := X"100BA7F0";
        ram_buffer(76792) := X"100BA7F0";
        ram_buffer(76793) := X"100BA7F0";
        ram_buffer(76794) := X"100BA7F0";
        ram_buffer(76795) := X"100BA7F0";
        ram_buffer(76796) := X"100BA7F0";
        ram_buffer(76797) := X"100BA7F0";
        ram_buffer(76798) := X"100BA7F0";
        ram_buffer(76799) := X"100BA7F0";
        ram_buffer(76800) := X"100BA7F0";
        ram_buffer(76801) := X"100BA7F0";
        ram_buffer(76802) := X"100BA7F0";
        ram_buffer(76803) := X"100BA7F0";
        ram_buffer(76804) := X"100BA718";
        ram_buffer(76805) := X"100BA7F0";
        ram_buffer(76806) := X"100BA7F0";
        ram_buffer(76807) := X"100BA7F0";
        ram_buffer(76808) := X"100BA7F0";
        ram_buffer(76809) := X"100BA7F0";
        ram_buffer(76810) := X"100BA7F0";
        ram_buffer(76811) := X"100BA7F0";
        ram_buffer(76812) := X"100BA7F0";
        ram_buffer(76813) := X"100BA6D8";
        ram_buffer(76814) := X"100BA6D8";
        ram_buffer(76815) := X"100BA6D8";
        ram_buffer(76816) := X"100BA6D8";
        ram_buffer(76817) := X"100BA6D8";
        ram_buffer(76818) := X"100BA6D8";
        ram_buffer(76819) := X"100BA7F0";
        ram_buffer(76820) := X"100BA7F0";
        ram_buffer(76821) := X"100BA7F0";
        ram_buffer(76822) := X"100BA7F0";
        ram_buffer(76823) := X"100BA7F0";
        ram_buffer(76824) := X"100BA7F0";
        ram_buffer(76825) := X"100BA7F0";
        ram_buffer(76826) := X"100BA7F0";
        ram_buffer(76827) := X"100BA7F0";
        ram_buffer(76828) := X"100BA7F0";
        ram_buffer(76829) := X"100BA7F0";
        ram_buffer(76830) := X"100BA7F0";
        ram_buffer(76831) := X"100BA7F0";
        ram_buffer(76832) := X"100BA7F0";
        ram_buffer(76833) := X"100BA7F0";
        ram_buffer(76834) := X"100BA7F0";
        ram_buffer(76835) := X"100BA7F0";
        ram_buffer(76836) := X"100BA718";
        ram_buffer(76837) := X"000A0001";
        ram_buffer(76838) := X"00020003";
        ram_buffer(76839) := X"00040005";
        ram_buffer(76840) := X"00060007";
        ram_buffer(76841) := X"00080009";
        ram_buffer(76842) := X"000A000B";
        ram_buffer(76843) := X"000C000D";
        ram_buffer(76844) := X"000E000F";
        ram_buffer(76845) := X"00100000";
        ram_buffer(76846) := X"30313233";
        ram_buffer(76847) := X"34353637";
        ram_buffer(76848) := X"38396162";
        ram_buffer(76849) := X"63646566";
        ram_buffer(76850) := X"00000000";
        ram_buffer(76851) := X"286E756C";
        ram_buffer(76852) := X"6C290000";
        ram_buffer(76853) := X"30313233";
        ram_buffer(76854) := X"34353637";
        ram_buffer(76855) := X"38394142";
        ram_buffer(76856) := X"43444546";
        ram_buffer(76857) := X"00000000";
        ram_buffer(76858) := X"62756720";
        ram_buffer(76859) := X"696E2076";
        ram_buffer(76860) := X"66707269";
        ram_buffer(76861) := X"6E74663A";
        ram_buffer(76862) := X"20626164";
        ram_buffer(76863) := X"20626173";
        ram_buffer(76864) := X"65000000";
        ram_buffer(76865) := X"100BB294";
        ram_buffer(76866) := X"100BC0E8";
        ram_buffer(76867) := X"100BC0E8";
        ram_buffer(76868) := X"100BB2B4";
        ram_buffer(76869) := X"100BC0E8";
        ram_buffer(76870) := X"100BC0E8";
        ram_buffer(76871) := X"100BC0E8";
        ram_buffer(76872) := X"100BB210";
        ram_buffer(76873) := X"100BC0E8";
        ram_buffer(76874) := X"100BC0E8";
        ram_buffer(76875) := X"100BB2C0";
        ram_buffer(76876) := X"100BB310";
        ram_buffer(76877) := X"100BC0E8";
        ram_buffer(76878) := X"100BB304";
        ram_buffer(76879) := X"100BB320";
        ram_buffer(76880) := X"100BC0E8";
        ram_buffer(76881) := X"100BB3E4";
        ram_buffer(76882) := X"100BB3F0";
        ram_buffer(76883) := X"100BB3F0";
        ram_buffer(76884) := X"100BB3F0";
        ram_buffer(76885) := X"100BB3F0";
        ram_buffer(76886) := X"100BB3F0";
        ram_buffer(76887) := X"100BB3F0";
        ram_buffer(76888) := X"100BB3F0";
        ram_buffer(76889) := X"100BB3F0";
        ram_buffer(76890) := X"100BB3F0";
        ram_buffer(76891) := X"100BC0E8";
        ram_buffer(76892) := X"100BC0E8";
        ram_buffer(76893) := X"100BC0E8";
        ram_buffer(76894) := X"100BC0E8";
        ram_buffer(76895) := X"100BC0E8";
        ram_buffer(76896) := X"100BC0E8";
        ram_buffer(76897) := X"100BC0E8";
        ram_buffer(76898) := X"100BC0E8";
        ram_buffer(76899) := X"100BC0E8";
        ram_buffer(76900) := X"100BB4B0";
        ram_buffer(76901) := X"100BB4EC";
        ram_buffer(76902) := X"100BC0E8";
        ram_buffer(76903) := X"100BC0E8";
        ram_buffer(76904) := X"100BC0E8";
        ram_buffer(76905) := X"100BC0E8";
        ram_buffer(76906) := X"100BC0E8";
        ram_buffer(76907) := X"100BC0E8";
        ram_buffer(76908) := X"100BC0E8";
        ram_buffer(76909) := X"100BC0E8";
        ram_buffer(76910) := X"100BC0E8";
        ram_buffer(76911) := X"100BC0E8";
        ram_buffer(76912) := X"100BB794";
        ram_buffer(76913) := X"100BC0E8";
        ram_buffer(76914) := X"100BC0E8";
        ram_buffer(76915) := X"100BC0E8";
        ram_buffer(76916) := X"100BB92C";
        ram_buffer(76917) := X"100BC0E8";
        ram_buffer(76918) := X"100BBA00";
        ram_buffer(76919) := X"100BC0E8";
        ram_buffer(76920) := X"100BC0E8";
        ram_buffer(76921) := X"100BBB60";
        ram_buffer(76922) := X"100BC0E8";
        ram_buffer(76923) := X"100BC0E8";
        ram_buffer(76924) := X"100BC0E8";
        ram_buffer(76925) := X"100BC0E8";
        ram_buffer(76926) := X"100BC0E8";
        ram_buffer(76927) := X"100BC0E8";
        ram_buffer(76928) := X"100BC0E8";
        ram_buffer(76929) := X"100BC0E8";
        ram_buffer(76930) := X"100BC0E8";
        ram_buffer(76931) := X"100BC0E8";
        ram_buffer(76932) := X"100BB4B0";
        ram_buffer(76933) := X"100BB4F0";
        ram_buffer(76934) := X"100BC0E8";
        ram_buffer(76935) := X"100BC0E8";
        ram_buffer(76936) := X"100BC0E8";
        ram_buffer(76937) := X"100BB440";
        ram_buffer(76938) := X"100BB4F0";
        ram_buffer(76939) := X"100BB4A4";
        ram_buffer(76940) := X"100BC0E8";
        ram_buffer(76941) := X"100BB46C";
        ram_buffer(76942) := X"100BC0E8";
        ram_buffer(76943) := X"100BB674";
        ram_buffer(76944) := X"100BB798";
        ram_buffer(76945) := X"100BB8D8";
        ram_buffer(76946) := X"100BB498";
        ram_buffer(76947) := X"100BC0E8";
        ram_buffer(76948) := X"100BB92C";
        ram_buffer(76949) := X"100BB1CC";
        ram_buffer(76950) := X"100BBA04";
        ram_buffer(76951) := X"100BC0E8";
        ram_buffer(76952) := X"100BC0E8";
        ram_buffer(76953) := X"100BBB74";
        ram_buffer(76954) := X"100BC0E8";
        ram_buffer(76955) := X"100BB1CC";
        ram_buffer(76956) := X"20202020";
        ram_buffer(76957) := X"20202020";
        ram_buffer(76958) := X"20202020";
        ram_buffer(76959) := X"20202020";
        ram_buffer(76960) := X"30303030";
        ram_buffer(76961) := X"30303030";
        ram_buffer(76962) := X"30303030";
        ram_buffer(76963) := X"30303030";
        ram_buffer(76964) := X"00000000";
        ram_buffer(76965) := X"00000000";
        ram_buffer(76966) := X"00000000";
        ram_buffer(76967) := X"00000000";
        ram_buffer(76968) := X"00000000";
        ram_buffer(76969) := X"00000000";
        ram_buffer(76970) := X"00000000";
        ram_buffer(76971) := X"00000000";
        ram_buffer(76972) := X"00000000";
        ram_buffer(76973) := X"00000000";
        ram_buffer(76974) := X"00000000";
        ram_buffer(76975) := X"00000000";
        ram_buffer(76976) := X"10111213";
        ram_buffer(76977) := X"14151617";
        ram_buffer(76978) := X"18190000";
        ram_buffer(76979) := X"00000000";
        ram_buffer(76980) := X"001A1B1C";
        ram_buffer(76981) := X"1D1E1F00";
        ram_buffer(76982) := X"00000000";
        ram_buffer(76983) := X"00000000";
        ram_buffer(76984) := X"00000000";
        ram_buffer(76985) := X"00000000";
        ram_buffer(76986) := X"00000000";
        ram_buffer(76987) := X"00000000";
        ram_buffer(76988) := X"001A1B1C";
        ram_buffer(76989) := X"1D1E1F00";
        ram_buffer(76990) := X"00000000";
        ram_buffer(76991) := X"00000000";
        ram_buffer(76992) := X"00000000";
        ram_buffer(76993) := X"00000000";
        ram_buffer(76994) := X"00000000";
        ram_buffer(76995) := X"00000000";
        ram_buffer(76996) := X"00000000";
        ram_buffer(76997) := X"00000000";
        ram_buffer(76998) := X"00000000";
        ram_buffer(76999) := X"00000000";
        ram_buffer(77000) := X"00000000";
        ram_buffer(77001) := X"00000000";
        ram_buffer(77002) := X"00000000";
        ram_buffer(77003) := X"00000000";
        ram_buffer(77004) := X"00000000";
        ram_buffer(77005) := X"00000000";
        ram_buffer(77006) := X"00000000";
        ram_buffer(77007) := X"00000000";
        ram_buffer(77008) := X"00000000";
        ram_buffer(77009) := X"00000000";
        ram_buffer(77010) := X"00000000";
        ram_buffer(77011) := X"00000000";
        ram_buffer(77012) := X"00000000";
        ram_buffer(77013) := X"00000000";
        ram_buffer(77014) := X"00000000";
        ram_buffer(77015) := X"00000000";
        ram_buffer(77016) := X"00000000";
        ram_buffer(77017) := X"00000000";
        ram_buffer(77018) := X"00000000";
        ram_buffer(77019) := X"00000000";
        ram_buffer(77020) := X"00000000";
        ram_buffer(77021) := X"00000000";
        ram_buffer(77022) := X"00000000";
        ram_buffer(77023) := X"00000000";
        ram_buffer(77024) := X"00000000";
        ram_buffer(77025) := X"00000000";
        ram_buffer(77026) := X"00000000";
        ram_buffer(77027) := X"00000000";
        ram_buffer(77028) := X"5F657869";
        ram_buffer(77029) := X"74282920";
        ram_buffer(77030) := X"73797363";
        ram_buffer(77031) := X"616C6C00";
        ram_buffer(77032) := X"4F757420";
        ram_buffer(77033) := X"6F662068";
        ram_buffer(77034) := X"65617020";
        ram_buffer(77035) := X"6D656D6F";
        ram_buffer(77036) := X"72790A00";
        ram_buffer(77037) := X"466C6173";
        ram_buffer(77038) := X"68436C65";
        ram_buffer(77039) := X"616E7570";
        ram_buffer(77040) := X"00000000";
        ram_buffer(77041) := X"4F70656E";
        ram_buffer(77042) := X"696E6720";
        ram_buffer(77043) := X"25732064";
        ram_buffer(77044) := X"69726563";
        ram_buffer(77045) := X"746F7279";
        ram_buffer(77046) := X"20666F72";
        ram_buffer(77047) := X"2025730A";
        ram_buffer(77048) := X"00000000";
        ram_buffer(77049) := X"656E646F";
        ram_buffer(77050) := X"6666696C";
        ram_buffer(77051) := X"65000000";
        ram_buffer(77052) := X"2F000000";
        ram_buffer(77053) := X"772B0000";
        ram_buffer(77054) := X"4552524F";
        ram_buffer(77055) := X"523A2043";
        ram_buffer(77056) := X"616E6E6F";
        ram_buffer(77057) := X"74206F70";
        ram_buffer(77058) := X"656E2066";
        ram_buffer(77059) := X"696C6520";
        ram_buffer(77060) := X"25730A00";
        ram_buffer(77061) := X"4552524F";
        ram_buffer(77062) := X"52207768";
        ram_buffer(77063) := X"696C6520";
        ram_buffer(77064) := X"72656164";
        ram_buffer(77065) := X"696E6720";
        ram_buffer(77066) := X"25733A20";
        ram_buffer(77067) := X"72656164";
        ram_buffer(77068) := X"20256420";
        ram_buffer(77069) := X"62797465";
        ram_buffer(77070) := X"732C2066";
        ram_buffer(77071) := X"696C6520";
        ram_buffer(77072) := X"73697A65";
        ram_buffer(77073) := X"20256420";
        ram_buffer(77074) := X"62797465";
        ram_buffer(77075) := X"730A0000";
        ram_buffer(77076) := X"4552524F";
        ram_buffer(77077) := X"523A2057";
        ram_buffer(77078) := X"726F6E67";
        ram_buffer(77079) := X"206F7574";
        ram_buffer(77080) := X"70757420";
        ram_buffer(77081) := X"66696C65";
        ram_buffer(77082) := X"0A000000";
        ram_buffer(77083) := X"434F5252";
        ram_buffer(77084) := X"45435421";
        ram_buffer(77085) := X"0A000000";
        ram_buffer(77086) := X"54727969";
        ram_buffer(77087) := X"6E672074";
        ram_buffer(77088) := X"6F206F70";
        ram_buffer(77089) := X"656E2025";
        ram_buffer(77090) := X"730A0000";
        ram_buffer(77091) := X"4572726F";
        ram_buffer(77092) := X"72206F70";
        ram_buffer(77093) := X"656E696E";
        ram_buffer(77094) := X"67202573";
        ram_buffer(77095) := X"0A000000";
        ram_buffer(77096) := X"52657375";
        ram_buffer(77097) := X"6C74206F";
        ram_buffer(77098) := X"66204F53";
        ram_buffer(77099) := X"5F666469";
        ram_buffer(77100) := X"72282573";
        ram_buffer(77101) := X"293A2025";
        ram_buffer(77102) := X"640A0000";
        ram_buffer(77103) := X"2F257300";
        ram_buffer(77104) := X"25732F25";
        ram_buffer(77105) := X"73000000";
        ram_buffer(77106) := X"456E7465";
        ram_buffer(77107) := X"72696E67";
        ram_buffer(77108) := X"20696E20";
        ram_buffer(77109) := X"64697265";
        ram_buffer(77110) := X"63746F72";
        ram_buffer(77111) := X"79202573";
        ram_buffer(77112) := X"0A000000";
        ram_buffer(77113) := X"25732025";
        ram_buffer(77114) := X"640A0000";
        ram_buffer(77115) := X"2F646972";
        ram_buffer(77116) := X"2F737562";
        ram_buffer(77117) := X"64697200";
        ram_buffer(77118) := X"77000000";
        ram_buffer(77119) := X"2F646972";
        ram_buffer(77120) := X"2F737562";
        ram_buffer(77121) := X"6469722F";
        ram_buffer(77122) := X"74657374";
        ram_buffer(77123) := X"2E747874";
        ram_buffer(77124) := X"00000000";
        ram_buffer(77125) := X"28257329";
        ram_buffer(77126) := X"0A000000";
        ram_buffer(77127) := X"2F646972";
        ram_buffer(77128) := X"25640000";
        ram_buffer(77129) := X"2F646972";
        ram_buffer(77130) := X"25642F66";
        ram_buffer(77131) := X"696C6525";
        ram_buffer(77132) := X"64256400";
        ram_buffer(77133) := X"693D2564";
        ram_buffer(77134) := X"206A3D25";
        ram_buffer(77135) := X"64000000";
        ram_buffer(77136) := X"2F646972";
        ram_buffer(77137) := X"312F6669";
        ram_buffer(77138) := X"6C653132";
        ram_buffer(77139) := X"00000000";
        ram_buffer(77140) := X"2F626164";
        ram_buffer(77141) := X"6469722F";
        ram_buffer(77142) := X"6D796669";
        ram_buffer(77143) := X"6C652E74";
        ram_buffer(77144) := X"78740000";
        ram_buffer(77145) := X"4552524F";
        ram_buffer(77146) := X"52210000";
        ram_buffer(77147) := X"693D2564";
        ram_buffer(77148) := X"206A3D25";
        ram_buffer(77149) := X"6420636F";
        ram_buffer(77150) := X"756E743D";
        ram_buffer(77151) := X"25642028";
        ram_buffer(77152) := X"2573290A";
        ram_buffer(77153) := X"00000000";
        ram_buffer(77154) := X"2F646972";
        ram_buffer(77155) := X"00000000";
        ram_buffer(77156) := X"496E7465";
        ram_buffer(77157) := X"72727570";
        ram_buffer(77158) := X"74212121";
        ram_buffer(77159) := X"21212100";
        ram_buffer(77160) := X"100C3E48";
        ram_buffer(77161) := X"100C3D14";
        ram_buffer(77162) := X"100C3D14";
        ram_buffer(77163) := X"100C3D10";
        ram_buffer(77164) := X"100C3E2C";
        ram_buffer(77165) := X"100C3E2C";
        ram_buffer(77166) := X"100C3E08";
        ram_buffer(77167) := X"100C3D10";
        ram_buffer(77168) := X"100C3E2C";
        ram_buffer(77169) := X"100C3E08";
        ram_buffer(77170) := X"100C3E2C";
        ram_buffer(77171) := X"100C3D10";
        ram_buffer(77172) := X"100C3E38";
        ram_buffer(77173) := X"100C3E38";
        ram_buffer(77174) := X"100C3E38";
        ram_buffer(77175) := X"100C3EEC";
        ram_buffer(77176) := X"100C5448";
        ram_buffer(77177) := X"100C52C0";
        ram_buffer(77178) := X"100C5358";
        ram_buffer(77179) := X"100C5328";
        ram_buffer(77180) := X"100C5358";
        ram_buffer(77181) := X"100C5420";
        ram_buffer(77182) := X"100C5358";
        ram_buffer(77183) := X"100C5328";
        ram_buffer(77184) := X"100C52C0";
        ram_buffer(77185) := X"100C52C0";
        ram_buffer(77186) := X"100C5420";
        ram_buffer(77187) := X"100C5328";
        ram_buffer(77188) := X"100C5338";
        ram_buffer(77189) := X"100C5338";
        ram_buffer(77190) := X"100C5338";
        ram_buffer(77191) := X"100C546C";
        ram_buffer(77192) := X"100C6058";
        ram_buffer(77193) := X"100C5EC0";
        ram_buffer(77194) := X"100C5EC0";
        ram_buffer(77195) := X"100C5EBC";
        ram_buffer(77196) := X"100C6034";
        ram_buffer(77197) := X"100C6034";
        ram_buffer(77198) := X"100C600C";
        ram_buffer(77199) := X"100C5EBC";
        ram_buffer(77200) := X"100C6034";
        ram_buffer(77201) := X"100C600C";
        ram_buffer(77202) := X"100C6034";
        ram_buffer(77203) := X"100C5EBC";
        ram_buffer(77204) := X"100C6044";
        ram_buffer(77205) := X"100C6044";
        ram_buffer(77206) := X"100C6044";
        ram_buffer(77207) := X"100C61A0";
        ram_buffer(77208) := X"00010202";
        ram_buffer(77209) := X"03030303";
        ram_buffer(77210) := X"04040404";
        ram_buffer(77211) := X"04040404";
        ram_buffer(77212) := X"05050505";
        ram_buffer(77213) := X"05050505";
        ram_buffer(77214) := X"05050505";
        ram_buffer(77215) := X"05050505";
        ram_buffer(77216) := X"06060606";
        ram_buffer(77217) := X"06060606";
        ram_buffer(77218) := X"06060606";
        ram_buffer(77219) := X"06060606";
        ram_buffer(77220) := X"06060606";
        ram_buffer(77221) := X"06060606";
        ram_buffer(77222) := X"06060606";
        ram_buffer(77223) := X"06060606";
        ram_buffer(77224) := X"07070707";
        ram_buffer(77225) := X"07070707";
        ram_buffer(77226) := X"07070707";
        ram_buffer(77227) := X"07070707";
        ram_buffer(77228) := X"07070707";
        ram_buffer(77229) := X"07070707";
        ram_buffer(77230) := X"07070707";
        ram_buffer(77231) := X"07070707";
        ram_buffer(77232) := X"07070707";
        ram_buffer(77233) := X"07070707";
        ram_buffer(77234) := X"07070707";
        ram_buffer(77235) := X"07070707";
        ram_buffer(77236) := X"07070707";
        ram_buffer(77237) := X"07070707";
        ram_buffer(77238) := X"07070707";
        ram_buffer(77239) := X"07070707";
        ram_buffer(77240) := X"08080808";
        ram_buffer(77241) := X"08080808";
        ram_buffer(77242) := X"08080808";
        ram_buffer(77243) := X"08080808";
        ram_buffer(77244) := X"08080808";
        ram_buffer(77245) := X"08080808";
        ram_buffer(77246) := X"08080808";
        ram_buffer(77247) := X"08080808";
        ram_buffer(77248) := X"08080808";
        ram_buffer(77249) := X"08080808";
        ram_buffer(77250) := X"08080808";
        ram_buffer(77251) := X"08080808";
        ram_buffer(77252) := X"08080808";
        ram_buffer(77253) := X"08080808";
        ram_buffer(77254) := X"08080808";
        ram_buffer(77255) := X"08080808";
        ram_buffer(77256) := X"08080808";
        ram_buffer(77257) := X"08080808";
        ram_buffer(77258) := X"08080808";
        ram_buffer(77259) := X"08080808";
        ram_buffer(77260) := X"08080808";
        ram_buffer(77261) := X"08080808";
        ram_buffer(77262) := X"08080808";
        ram_buffer(77263) := X"08080808";
        ram_buffer(77264) := X"08080808";
        ram_buffer(77265) := X"08080808";
        ram_buffer(77266) := X"08080808";
        ram_buffer(77267) := X"08080808";
        ram_buffer(77268) := X"08080808";
        ram_buffer(77269) := X"08080808";
        ram_buffer(77270) := X"08080808";
        ram_buffer(77271) := X"08080808";
        ram_buffer(77272) := X"00000010";
        ram_buffer(77273) := X"00000000";
        ram_buffer(77274) := X"017A5200";
        ram_buffer(77275) := X"017C1F01";
        ram_buffer(77276) := X"0B0D1D00";
        ram_buffer(77277) := X"00000010";
        ram_buffer(77278) := X"00000018";
        ram_buffer(77279) := X"100C299C";
        ram_buffer(77280) := X"0000065C";
        ram_buffer(77281) := X"00000000";
        ram_buffer(77282) := X"00000010";
        ram_buffer(77283) := X"0000002C";
        ram_buffer(77284) := X"100C2FF8";
        ram_buffer(77285) := X"0000064C";
        ram_buffer(77286) := X"00000000";
        ram_buffer(77287) := X"00000000";
        ram_buffer(77288) := X"00000000";
        ram_buffer(77289) := X"00000000";
        ram_buffer(77290) := X"00000000";
        ram_buffer(77291) := X"00000000";
        ram_buffer(77292) := X"00000000";
        ram_buffer(77293) := X"00000000";
        ram_buffer(77294) := X"00000000";
        ram_buffer(77295) := X"00000000";
        ram_buffer(77296) := X"00000000";
        ram_buffer(77297) := X"00000000";
        ram_buffer(77298) := X"00000000";
        ram_buffer(77299) := X"00000000";
        ram_buffer(77300) := X"00000000";
        ram_buffer(77301) := X"00000000";
        ram_buffer(77302) := X"00000000";
        ram_buffer(77303) := X"00000000";
        ram_buffer(77304) := X"00000000";
        ram_buffer(77305) := X"00000000";
        ram_buffer(77306) := X"00000000";
        ram_buffer(77307) := X"00000000";
        ram_buffer(77308) := X"00000000";
        ram_buffer(77309) := X"00000000";
        ram_buffer(77310) := X"00000000";
        ram_buffer(77311) := X"00000000";
        ram_buffer(77312) := X"00000000";
        ram_buffer(77313) := X"00000000";
        ram_buffer(77314) := X"00000000";
        ram_buffer(77315) := X"00000000";
        ram_buffer(77316) := X"00000000";
        ram_buffer(77317) := X"00000000";
        ram_buffer(77318) := X"00000000";
        ram_buffer(77319) := X"00000000";
        ram_buffer(77320) := X"00000000";
        ram_buffer(77321) := X"00000000";
        ram_buffer(77322) := X"00000000";
        ram_buffer(77323) := X"00000000";
        ram_buffer(77324) := X"00000000";
        ram_buffer(77325) := X"00000000";
        ram_buffer(77326) := X"00000000";
        ram_buffer(77327) := X"00000000";
        ram_buffer(77328) := X"00000000";
        ram_buffer(77329) := X"00000000";
        ram_buffer(77330) := X"00000000";
        ram_buffer(77331) := X"00000000";
        ram_buffer(77332) := X"00000000";
        ram_buffer(77333) := X"00000000";
        ram_buffer(77334) := X"00000000";
        ram_buffer(77335) := X"00000000";
        ram_buffer(77336) := X"00000000";
        ram_buffer(77337) := X"00000000";
        ram_buffer(77338) := X"00000000";
        ram_buffer(77339) := X"00000000";
        ram_buffer(77340) := X"00000000";
        ram_buffer(77341) := X"00000000";
        ram_buffer(77342) := X"00000000";
        ram_buffer(77343) := X"00000000";
        ram_buffer(77344) := X"00000000";
        ram_buffer(77345) := X"00000000";
        ram_buffer(77346) := X"00000000";
        ram_buffer(77347) := X"00000000";
        ram_buffer(77348) := X"00000000";
        ram_buffer(77349) := X"00000000";
        ram_buffer(77350) := X"00000000";
        ram_buffer(77351) := X"00000000";
        ram_buffer(77352) := X"00000000";
        ram_buffer(77353) := X"00000000";
        ram_buffer(77354) := X"00000000";
        ram_buffer(77355) := X"00000000";
        ram_buffer(77356) := X"00000000";
        ram_buffer(77357) := X"00000000";
        ram_buffer(77358) := X"00000000";
        ram_buffer(77359) := X"00000000";
        ram_buffer(77360) := X"00000000";
        ram_buffer(77361) := X"00000000";
        ram_buffer(77362) := X"00000000";
        ram_buffer(77363) := X"00000000";
        ram_buffer(77364) := X"00000000";
        ram_buffer(77365) := X"00000000";
        ram_buffer(77366) := X"00000000";
        ram_buffer(77367) := X"00000000";
        ram_buffer(77368) := X"00000000";
        ram_buffer(77369) := X"00000000";
        ram_buffer(77370) := X"00000000";
        ram_buffer(77371) := X"00000000";
        ram_buffer(77372) := X"00000000";
        ram_buffer(77373) := X"00000000";
        ram_buffer(77374) := X"00000000";
        ram_buffer(77375) := X"00000000";
        ram_buffer(77376) := X"00000000";
        ram_buffer(77377) := X"00000000";
        ram_buffer(77378) := X"00000000";
        ram_buffer(77379) := X"00000000";
        ram_buffer(77380) := X"00000000";
        ram_buffer(77381) := X"00000000";
        ram_buffer(77382) := X"00000000";
        ram_buffer(77383) := X"00000000";
        ram_buffer(77384) := X"00000000";
        ram_buffer(77385) := X"00000000";
        ram_buffer(77386) := X"00000000";
        ram_buffer(77387) := X"00000000";
        ram_buffer(77388) := X"00000000";
        ram_buffer(77389) := X"00000000";
        ram_buffer(77390) := X"00000000";
        ram_buffer(77391) := X"00000000";
        ram_buffer(77392) := X"00000000";
        ram_buffer(77393) := X"00000000";
        ram_buffer(77394) := X"00000000";
        ram_buffer(77395) := X"00000000";
        ram_buffer(77396) := X"00000000";
        ram_buffer(77397) := X"00000000";
        ram_buffer(77398) := X"00000000";
        ram_buffer(77399) := X"00000000";
        ram_buffer(77400) := X"00000000";
        ram_buffer(77401) := X"00000000";
        ram_buffer(77402) := X"00000000";
        ram_buffer(77403) := X"00000000";
        ram_buffer(77404) := X"00000000";
        ram_buffer(77405) := X"00000000";
        ram_buffer(77406) := X"00000000";
        ram_buffer(77407) := X"00000000";
        ram_buffer(77408) := X"00000000";
        ram_buffer(77409) := X"00000000";
        ram_buffer(77410) := X"00000000";
        ram_buffer(77411) := X"00000000";
        ram_buffer(77412) := X"00000000";
        ram_buffer(77413) := X"00000000";
        ram_buffer(77414) := X"00000000";
        ram_buffer(77415) := X"00000000";
        ram_buffer(77416) := X"00000000";
        ram_buffer(77417) := X"00000000";
        ram_buffer(77418) := X"00000000";
        ram_buffer(77419) := X"00000000";
        ram_buffer(77420) := X"00000000";
        ram_buffer(77421) := X"00000000";
        ram_buffer(77422) := X"00000000";
        ram_buffer(77423) := X"00000000";
        ram_buffer(77424) := X"00000000";
        ram_buffer(77425) := X"00000000";
        ram_buffer(77426) := X"00000000";
        ram_buffer(77427) := X"00000000";
        ram_buffer(77428) := X"00000000";
        ram_buffer(77429) := X"00000000";
        ram_buffer(77430) := X"00000000";
        ram_buffer(77431) := X"00000000";
        ram_buffer(77432) := X"00000000";
        ram_buffer(77433) := X"00000000";
        ram_buffer(77434) := X"00000000";
        ram_buffer(77435) := X"00000000";
        ram_buffer(77436) := X"00000000";
        ram_buffer(77437) := X"00000000";
        ram_buffer(77438) := X"00000000";
        ram_buffer(77439) := X"00000000";
        ram_buffer(77440) := X"00000000";
        ram_buffer(77441) := X"00000000";
        ram_buffer(77442) := X"00000000";
        ram_buffer(77443) := X"00000000";
        ram_buffer(77444) := X"00000000";
        ram_buffer(77445) := X"00000000";
        ram_buffer(77446) := X"00000000";
        ram_buffer(77447) := X"00000000";
        ram_buffer(77448) := X"00000000";
        ram_buffer(77449) := X"00000000";
        ram_buffer(77450) := X"00000000";
        ram_buffer(77451) := X"00000000";
        ram_buffer(77452) := X"00000000";
        ram_buffer(77453) := X"00000000";
        ram_buffer(77454) := X"00000000";
        ram_buffer(77455) := X"00000000";
        ram_buffer(77456) := X"00000000";
        ram_buffer(77457) := X"00000000";
        ram_buffer(77458) := X"00000000";
        ram_buffer(77459) := X"00000000";
        ram_buffer(77460) := X"00000000";
        ram_buffer(77461) := X"00000000";
        ram_buffer(77462) := X"00000000";
        ram_buffer(77463) := X"00000000";
        ram_buffer(77464) := X"00000000";
        ram_buffer(77465) := X"00000000";
        ram_buffer(77466) := X"00000000";
        ram_buffer(77467) := X"00000000";
        ram_buffer(77468) := X"00000000";
        ram_buffer(77469) := X"00000000";
        ram_buffer(77470) := X"00000000";
        ram_buffer(77471) := X"00000000";
        ram_buffer(77472) := X"00000000";
        ram_buffer(77473) := X"00000000";
        ram_buffer(77474) := X"00000000";
        ram_buffer(77475) := X"00000000";
        ram_buffer(77476) := X"00000000";
        ram_buffer(77477) := X"00000000";
        ram_buffer(77478) := X"00000000";
        ram_buffer(77479) := X"00000000";
        ram_buffer(77480) := X"00000000";
        ram_buffer(77481) := X"00000000";
        ram_buffer(77482) := X"00000000";
        ram_buffer(77483) := X"00000000";
        ram_buffer(77484) := X"00000000";
        ram_buffer(77485) := X"00000000";
        ram_buffer(77486) := X"00000000";
        ram_buffer(77487) := X"00000000";
        ram_buffer(77488) := X"00000000";
        ram_buffer(77489) := X"00000000";
        ram_buffer(77490) := X"00000000";
        ram_buffer(77491) := X"00000000";
        ram_buffer(77492) := X"00000000";
        ram_buffer(77493) := X"00000000";
        ram_buffer(77494) := X"00000000";
        ram_buffer(77495) := X"00000000";
        ram_buffer(77496) := X"00000000";
        ram_buffer(77497) := X"00000000";
        ram_buffer(77498) := X"00000000";
        ram_buffer(77499) := X"00000000";
        ram_buffer(77500) := X"00000000";
        ram_buffer(77501) := X"00000000";
        ram_buffer(77502) := X"00000000";
        ram_buffer(77503) := X"00000000";
        ram_buffer(77504) := X"00000000";
        ram_buffer(77505) := X"00000000";
        ram_buffer(77506) := X"00000000";
        ram_buffer(77507) := X"00000000";
        ram_buffer(77508) := X"00000000";
        ram_buffer(77509) := X"00000000";
        ram_buffer(77510) := X"00000000";
        ram_buffer(77511) := X"00000000";
        ram_buffer(77512) := X"00000000";
        ram_buffer(77513) := X"00000000";
        ram_buffer(77514) := X"00000000";
        ram_buffer(77515) := X"00000000";
        ram_buffer(77516) := X"00000000";
        ram_buffer(77517) := X"00000000";
        ram_buffer(77518) := X"00000000";
        ram_buffer(77519) := X"00000000";
        ram_buffer(77520) := X"00000000";
        ram_buffer(77521) := X"00000000";
        ram_buffer(77522) := X"00000000";
        ram_buffer(77523) := X"00000000";
        ram_buffer(77524) := X"00000000";
        ram_buffer(77525) := X"00000000";
        ram_buffer(77526) := X"00000000";
        ram_buffer(77527) := X"00000000";
        ram_buffer(77528) := X"00000000";
        ram_buffer(77529) := X"00000000";
        ram_buffer(77530) := X"00000000";
        ram_buffer(77531) := X"00000000";
        ram_buffer(77532) := X"00000000";
        ram_buffer(77533) := X"00000000";
        ram_buffer(77534) := X"00000000";
        ram_buffer(77535) := X"00000000";
        ram_buffer(77536) := X"00000000";
        ram_buffer(77537) := X"00000000";
        ram_buffer(77538) := X"00000000";
        ram_buffer(77539) := X"00000000";
        ram_buffer(77540) := X"00000000";
        ram_buffer(77541) := X"00000000";
        ram_buffer(77542) := X"00000000";
        ram_buffer(77543) := X"00000000";
        ram_buffer(77544) := X"00000000";
        ram_buffer(77545) := X"00000000";
        ram_buffer(77546) := X"00000000";
        ram_buffer(77547) := X"00000000";
        ram_buffer(77548) := X"00000000";
        ram_buffer(77549) := X"00000000";
        ram_buffer(77550) := X"00000000";
        ram_buffer(77551) := X"00000000";
        ram_buffer(77552) := X"00000000";
        ram_buffer(77553) := X"00000000";
        ram_buffer(77554) := X"00000000";
        ram_buffer(77555) := X"00000000";
        ram_buffer(77556) := X"00000000";
        ram_buffer(77557) := X"00000000";
        ram_buffer(77558) := X"00000000";
        ram_buffer(77559) := X"00000000";
        ram_buffer(77560) := X"00000000";
        ram_buffer(77561) := X"00000000";
        ram_buffer(77562) := X"00000000";
        ram_buffer(77563) := X"00000000";
        ram_buffer(77564) := X"00000000";
        ram_buffer(77565) := X"00000000";
        ram_buffer(77566) := X"00000000";
        ram_buffer(77567) := X"00000000";
        ram_buffer(77568) := X"00000000";
        ram_buffer(77569) := X"00000000";
        ram_buffer(77570) := X"00000000";
        ram_buffer(77571) := X"00000000";
        ram_buffer(77572) := X"00000000";
        ram_buffer(77573) := X"00000000";
        ram_buffer(77574) := X"00000000";
        ram_buffer(77575) := X"00000000";
        ram_buffer(77576) := X"00000000";
        ram_buffer(77577) := X"00000000";
        ram_buffer(77578) := X"00000000";
        ram_buffer(77579) := X"00000000";
        ram_buffer(77580) := X"00000000";
        ram_buffer(77581) := X"00000000";
        ram_buffer(77582) := X"00000000";
        ram_buffer(77583) := X"00000000";
        ram_buffer(77584) := X"00000000";
        ram_buffer(77585) := X"00000000";
        ram_buffer(77586) := X"00000000";
        ram_buffer(77587) := X"00000000";
        ram_buffer(77588) := X"00000000";
        ram_buffer(77589) := X"00000000";
        ram_buffer(77590) := X"00000000";
        ram_buffer(77591) := X"00000000";
        ram_buffer(77592) := X"00000000";
        ram_buffer(77593) := X"00000000";
        ram_buffer(77594) := X"00000000";
        ram_buffer(77595) := X"00000000";
        ram_buffer(77596) := X"00000000";
        ram_buffer(77597) := X"00000000";
        ram_buffer(77598) := X"00000000";
        ram_buffer(77599) := X"00000000";
        ram_buffer(77600) := X"00000000";
        ram_buffer(77601) := X"00000000";
        ram_buffer(77602) := X"00000000";
        ram_buffer(77603) := X"00000000";
        ram_buffer(77604) := X"00000000";
        ram_buffer(77605) := X"00000000";
        ram_buffer(77606) := X"00000000";
        ram_buffer(77607) := X"00000000";
        ram_buffer(77608) := X"00000000";
        ram_buffer(77609) := X"00000000";
        ram_buffer(77610) := X"00000000";
        ram_buffer(77611) := X"00000000";
        ram_buffer(77612) := X"00000000";
        ram_buffer(77613) := X"00000000";
        ram_buffer(77614) := X"00000000";
        ram_buffer(77615) := X"00000000";
        ram_buffer(77616) := X"00000000";
        ram_buffer(77617) := X"00000000";
        ram_buffer(77618) := X"00000000";
        ram_buffer(77619) := X"00000000";
        ram_buffer(77620) := X"00000000";
        ram_buffer(77621) := X"00000000";
        ram_buffer(77622) := X"00000000";
        ram_buffer(77623) := X"00000000";
        ram_buffer(77624) := X"00000000";
        ram_buffer(77625) := X"00000000";
        ram_buffer(77626) := X"00000000";
        ram_buffer(77627) := X"00000000";
        ram_buffer(77628) := X"00000000";
        ram_buffer(77629) := X"00000000";
        ram_buffer(77630) := X"00000000";
        ram_buffer(77631) := X"00000000";
        ram_buffer(77632) := X"00000000";
        ram_buffer(77633) := X"00000000";
        ram_buffer(77634) := X"00000000";
        ram_buffer(77635) := X"00000000";
        ram_buffer(77636) := X"00000000";
        ram_buffer(77637) := X"00000000";
        ram_buffer(77638) := X"00000000";
        ram_buffer(77639) := X"00000000";
        ram_buffer(77640) := X"00000000";
        ram_buffer(77641) := X"00000000";
        ram_buffer(77642) := X"00000000";
        ram_buffer(77643) := X"00000000";
        ram_buffer(77644) := X"00000000";
        ram_buffer(77645) := X"00000000";
        ram_buffer(77646) := X"00000000";
        ram_buffer(77647) := X"00000000";
        ram_buffer(77648) := X"00000000";
        ram_buffer(77649) := X"00000000";
        ram_buffer(77650) := X"00000000";
        ram_buffer(77651) := X"00000000";
        ram_buffer(77652) := X"00000000";
        ram_buffer(77653) := X"00000000";
        ram_buffer(77654) := X"00000000";
        ram_buffer(77655) := X"00000000";
        ram_buffer(77656) := X"00000000";
        ram_buffer(77657) := X"00000000";
        ram_buffer(77658) := X"00000000";
        ram_buffer(77659) := X"00000000";
        ram_buffer(77660) := X"00000000";
        ram_buffer(77661) := X"00000000";
        ram_buffer(77662) := X"00000000";
        ram_buffer(77663) := X"00000000";
        ram_buffer(77664) := X"00000000";
        ram_buffer(77665) := X"00000000";
        ram_buffer(77666) := X"00000000";
        ram_buffer(77667) := X"00000000";
        ram_buffer(77668) := X"00000000";
        ram_buffer(77669) := X"00000000";
        ram_buffer(77670) := X"00000000";
        ram_buffer(77671) := X"00000000";
        ram_buffer(77672) := X"00000000";
        ram_buffer(77673) := X"00000000";
        ram_buffer(77674) := X"00000000";
        ram_buffer(77675) := X"00000000";
        ram_buffer(77676) := X"00000000";
        ram_buffer(77677) := X"00000000";
        ram_buffer(77678) := X"00000000";
        ram_buffer(77679) := X"00000000";
        ram_buffer(77680) := X"00000000";
        ram_buffer(77681) := X"00000000";
        ram_buffer(77682) := X"00000000";
        ram_buffer(77683) := X"00000000";
        ram_buffer(77684) := X"00000000";
        ram_buffer(77685) := X"00000000";
        ram_buffer(77686) := X"00000000";
        ram_buffer(77687) := X"00000000";
        ram_buffer(77688) := X"00000000";
        ram_buffer(77689) := X"00000000";
        ram_buffer(77690) := X"00000000";
        ram_buffer(77691) := X"00000000";
        ram_buffer(77692) := X"00000000";
        ram_buffer(77693) := X"00000000";
        ram_buffer(77694) := X"00000000";
        ram_buffer(77695) := X"00000000";
        ram_buffer(77696) := X"00000000";
        ram_buffer(77697) := X"00000000";
        ram_buffer(77698) := X"00000000";
        ram_buffer(77699) := X"00000000";
        ram_buffer(77700) := X"00000000";
        ram_buffer(77701) := X"00000000";
        ram_buffer(77702) := X"00000000";
        ram_buffer(77703) := X"00000000";
        ram_buffer(77704) := X"00000000";
        ram_buffer(77705) := X"00000000";
        ram_buffer(77706) := X"00000000";
        ram_buffer(77707) := X"00000000";
        ram_buffer(77708) := X"00000000";
        ram_buffer(77709) := X"00000000";
        ram_buffer(77710) := X"00000000";
        ram_buffer(77711) := X"00000000";
        ram_buffer(77712) := X"00000000";
        ram_buffer(77713) := X"00000000";
        ram_buffer(77714) := X"00000000";
        ram_buffer(77715) := X"00000000";
        ram_buffer(77716) := X"00000000";
        ram_buffer(77717) := X"00000000";
        ram_buffer(77718) := X"00000000";
        ram_buffer(77719) := X"00000000";
        ram_buffer(77720) := X"00000000";
        ram_buffer(77721) := X"00000000";
        ram_buffer(77722) := X"00000000";
        ram_buffer(77723) := X"00000000";
        ram_buffer(77724) := X"00000000";
        ram_buffer(77725) := X"00000000";
        ram_buffer(77726) := X"00000000";
        ram_buffer(77727) := X"00000000";
        ram_buffer(77728) := X"00000000";
        ram_buffer(77729) := X"00000000";
        ram_buffer(77730) := X"00000000";
        ram_buffer(77731) := X"00000000";
        ram_buffer(77732) := X"00000000";
        ram_buffer(77733) := X"00000000";
        ram_buffer(77734) := X"00000000";
        ram_buffer(77735) := X"00000000";
        ram_buffer(77736) := X"00000000";
        ram_buffer(77737) := X"00000000";
        ram_buffer(77738) := X"00000000";
        ram_buffer(77739) := X"00000000";
        ram_buffer(77740) := X"00000000";
        ram_buffer(77741) := X"00000000";
        ram_buffer(77742) := X"00000000";
        ram_buffer(77743) := X"00000000";
        ram_buffer(77744) := X"00000000";
        ram_buffer(77745) := X"00000000";
        ram_buffer(77746) := X"00000000";
        ram_buffer(77747) := X"00000000";
        ram_buffer(77748) := X"00000000";
        ram_buffer(77749) := X"00000000";
        ram_buffer(77750) := X"00000000";
        ram_buffer(77751) := X"00000000";
        ram_buffer(77752) := X"00000000";
        ram_buffer(77753) := X"00000000";
        ram_buffer(77754) := X"00000000";
        ram_buffer(77755) := X"00000000";
        ram_buffer(77756) := X"00000000";
        ram_buffer(77757) := X"00000000";
        ram_buffer(77758) := X"00000000";
        ram_buffer(77759) := X"00000000";
        ram_buffer(77760) := X"00000000";
        ram_buffer(77761) := X"00000000";
        ram_buffer(77762) := X"00000000";
        ram_buffer(77763) := X"00000000";
        ram_buffer(77764) := X"00000000";
        ram_buffer(77765) := X"00000000";
        ram_buffer(77766) := X"00000000";
        ram_buffer(77767) := X"00000000";
        ram_buffer(77768) := X"00000000";
        ram_buffer(77769) := X"00000000";
        ram_buffer(77770) := X"00000000";
        ram_buffer(77771) := X"00000000";
        ram_buffer(77772) := X"00000000";
        ram_buffer(77773) := X"00000000";
        ram_buffer(77774) := X"00000000";
        ram_buffer(77775) := X"00000000";
        ram_buffer(77776) := X"00000000";
        ram_buffer(77777) := X"00000000";
        ram_buffer(77778) := X"00000000";
        ram_buffer(77779) := X"00000000";
        ram_buffer(77780) := X"00000000";
        ram_buffer(77781) := X"00000000";
        ram_buffer(77782) := X"00000000";
        ram_buffer(77783) := X"00000000";
        ram_buffer(77784) := X"00000000";
        ram_buffer(77785) := X"00000000";
        ram_buffer(77786) := X"00000000";
        ram_buffer(77787) := X"00000000";
        ram_buffer(77788) := X"00000000";
        ram_buffer(77789) := X"00000000";
        ram_buffer(77790) := X"00000000";
        ram_buffer(77791) := X"00000000";
        ram_buffer(77792) := X"00000000";
        ram_buffer(77793) := X"00000000";
        ram_buffer(77794) := X"00000000";
        ram_buffer(77795) := X"00000000";
        ram_buffer(77796) := X"00000000";
        ram_buffer(77797) := X"00000000";
        ram_buffer(77798) := X"00000000";
        ram_buffer(77799) := X"00000000";
        ram_buffer(77800) := X"00000000";
        ram_buffer(77801) := X"00000000";
        ram_buffer(77802) := X"00000000";
        ram_buffer(77803) := X"00000000";
        ram_buffer(77804) := X"00000000";
        ram_buffer(77805) := X"00000000";
        ram_buffer(77806) := X"00000000";
        ram_buffer(77807) := X"00000000";
        ram_buffer(77808) := X"00000000";
        ram_buffer(77809) := X"00000000";
        ram_buffer(77810) := X"00000000";
        ram_buffer(77811) := X"00000000";
        ram_buffer(77812) := X"00000000";
        ram_buffer(77813) := X"00000000";
        ram_buffer(77814) := X"00000000";
        ram_buffer(77815) := X"00000000";
        ram_buffer(77816) := X"00000000";
        ram_buffer(77817) := X"00000000";
        ram_buffer(77818) := X"00000000";
        ram_buffer(77819) := X"00000000";
        ram_buffer(77820) := X"00000000";
        ram_buffer(77821) := X"00000000";
        ram_buffer(77822) := X"00000000";
        ram_buffer(77823) := X"00000000";
        ram_buffer(77824) := X"00000000";
        ram_buffer(77825) := X"00000000";
        ram_buffer(77826) := X"00000000";
        ram_buffer(77827) := X"00000000";
        ram_buffer(77828) := X"00000000";
        ram_buffer(77829) := X"00000000";
        ram_buffer(77830) := X"00000000";
        ram_buffer(77831) := X"00000000";
        ram_buffer(77832) := X"00000000";
        ram_buffer(77833) := X"00000000";
        ram_buffer(77834) := X"00000000";
        ram_buffer(77835) := X"00000000";
        ram_buffer(77836) := X"00000000";
        ram_buffer(77837) := X"00000000";
        ram_buffer(77838) := X"00000000";
        ram_buffer(77839) := X"00000000";
        ram_buffer(77840) := X"00000000";
        ram_buffer(77841) := X"00000000";
        ram_buffer(77842) := X"00000000";
        ram_buffer(77843) := X"00000000";
        ram_buffer(77844) := X"00000000";
        ram_buffer(77845) := X"00000000";
        ram_buffer(77846) := X"00000000";
        ram_buffer(77847) := X"00000000";
        ram_buffer(77848) := X"00000000";
        ram_buffer(77849) := X"00000000";
        ram_buffer(77850) := X"00000000";
        ram_buffer(77851) := X"00000000";
        ram_buffer(77852) := X"00000000";
        ram_buffer(77853) := X"00000000";
        ram_buffer(77854) := X"00000000";
        ram_buffer(77855) := X"00000000";
        ram_buffer(77856) := X"00000000";
        ram_buffer(77857) := X"00000000";
        ram_buffer(77858) := X"00000000";
        ram_buffer(77859) := X"00000000";
        ram_buffer(77860) := X"00000000";
        ram_buffer(77861) := X"00000000";
        ram_buffer(77862) := X"00000000";
        ram_buffer(77863) := X"00000000";
        ram_buffer(77864) := X"00000000";
        ram_buffer(77865) := X"00000000";
        ram_buffer(77866) := X"00000000";
        ram_buffer(77867) := X"00000000";
        ram_buffer(77868) := X"00000000";
        ram_buffer(77869) := X"00000000";
        ram_buffer(77870) := X"00000000";
        ram_buffer(77871) := X"00000000";
        ram_buffer(77872) := X"00000000";
        ram_buffer(77873) := X"00000000";
        ram_buffer(77874) := X"00000000";
        ram_buffer(77875) := X"00000000";
        ram_buffer(77876) := X"00000000";
        ram_buffer(77877) := X"00000000";
        ram_buffer(77878) := X"00000000";
        ram_buffer(77879) := X"00000000";
        ram_buffer(77880) := X"00000000";
        ram_buffer(77881) := X"00000000";
        ram_buffer(77882) := X"00000000";
        ram_buffer(77883) := X"00000000";
        ram_buffer(77884) := X"00000000";
        ram_buffer(77885) := X"00000000";
        ram_buffer(77886) := X"00000000";
        ram_buffer(77887) := X"00000000";
        ram_buffer(77888) := X"00000000";
        ram_buffer(77889) := X"00000000";
        ram_buffer(77890) := X"00000000";
        ram_buffer(77891) := X"00000000";
        ram_buffer(77892) := X"00000000";
        ram_buffer(77893) := X"00000000";
        ram_buffer(77894) := X"00000000";
        ram_buffer(77895) := X"00000000";
        ram_buffer(77896) := X"00000000";
        ram_buffer(77897) := X"00000000";
        ram_buffer(77898) := X"00000000";
        ram_buffer(77899) := X"00000000";
        ram_buffer(77900) := X"00000000";
        ram_buffer(77901) := X"00000000";
        ram_buffer(77902) := X"00000000";
        ram_buffer(77903) := X"00000000";
        ram_buffer(77904) := X"00000000";
        ram_buffer(77905) := X"00000000";
        ram_buffer(77906) := X"00000000";
        ram_buffer(77907) := X"00000000";
        ram_buffer(77908) := X"00000000";
        ram_buffer(77909) := X"00000000";
        ram_buffer(77910) := X"00000000";
        ram_buffer(77911) := X"00000000";
        ram_buffer(77912) := X"00000000";
        ram_buffer(77913) := X"00000000";
        ram_buffer(77914) := X"00000000";
        ram_buffer(77915) := X"00000000";
        ram_buffer(77916) := X"00000000";
        ram_buffer(77917) := X"00000000";
        ram_buffer(77918) := X"00000000";
        ram_buffer(77919) := X"00000000";
        ram_buffer(77920) := X"00000000";
        ram_buffer(77921) := X"00000000";
        ram_buffer(77922) := X"00000000";
        ram_buffer(77923) := X"00000000";
        ram_buffer(77924) := X"00000000";
        ram_buffer(77925) := X"00000000";
        ram_buffer(77926) := X"00000000";
        ram_buffer(77927) := X"00000000";
        ram_buffer(77928) := X"00000000";
        ram_buffer(77929) := X"00000000";
        ram_buffer(77930) := X"00000000";
        ram_buffer(77931) := X"00000000";
        ram_buffer(77932) := X"00000000";
        ram_buffer(77933) := X"00000000";
        ram_buffer(77934) := X"00000000";
        ram_buffer(77935) := X"00000000";
        ram_buffer(77936) := X"00000000";
        ram_buffer(77937) := X"00000000";
        ram_buffer(77938) := X"00000000";
        ram_buffer(77939) := X"00000000";
        ram_buffer(77940) := X"00000000";
        ram_buffer(77941) := X"00000000";
        ram_buffer(77942) := X"00000000";
        ram_buffer(77943) := X"00000000";
        ram_buffer(77944) := X"00000000";
        ram_buffer(77945) := X"00000000";
        ram_buffer(77946) := X"00000000";
        ram_buffer(77947) := X"00000000";
        ram_buffer(77948) := X"00000000";
        ram_buffer(77949) := X"00000000";
        ram_buffer(77950) := X"00000000";
        ram_buffer(77951) := X"00000000";
        ram_buffer(77952) := X"00000000";
        ram_buffer(77953) := X"00000000";
        ram_buffer(77954) := X"00000000";
        ram_buffer(77955) := X"00000000";
        ram_buffer(77956) := X"00000000";
        ram_buffer(77957) := X"00000000";
        ram_buffer(77958) := X"00000000";
        ram_buffer(77959) := X"00000000";
        ram_buffer(77960) := X"00000000";
        ram_buffer(77961) := X"00000000";
        ram_buffer(77962) := X"00000000";
        ram_buffer(77963) := X"00000000";
        ram_buffer(77964) := X"00000000";
        ram_buffer(77965) := X"00000000";
        ram_buffer(77966) := X"00000000";
        ram_buffer(77967) := X"00000000";
        ram_buffer(77968) := X"00000000";
        ram_buffer(77969) := X"00000000";
        ram_buffer(77970) := X"00000000";
        ram_buffer(77971) := X"00000000";
        ram_buffer(77972) := X"00000000";
        ram_buffer(77973) := X"00000000";
        ram_buffer(77974) := X"00000000";
        ram_buffer(77975) := X"00000000";
        ram_buffer(77976) := X"00000000";
        ram_buffer(77977) := X"00000000";
        ram_buffer(77978) := X"00000000";
        ram_buffer(77979) := X"00000000";
        ram_buffer(77980) := X"00000000";
        ram_buffer(77981) := X"00000000";
        ram_buffer(77982) := X"00000000";
        ram_buffer(77983) := X"00000000";
        ram_buffer(77984) := X"00000000";
        ram_buffer(77985) := X"00000000";
        ram_buffer(77986) := X"00000000";
        ram_buffer(77987) := X"00000000";
        ram_buffer(77988) := X"00000000";
        ram_buffer(77989) := X"00000000";
        ram_buffer(77990) := X"00000000";
        ram_buffer(77991) := X"00000000";
        ram_buffer(77992) := X"00000000";
        ram_buffer(77993) := X"00000000";
        ram_buffer(77994) := X"00000000";
        ram_buffer(77995) := X"00000000";
        ram_buffer(77996) := X"00000000";
        ram_buffer(77997) := X"00000000";
        ram_buffer(77998) := X"00000000";
        ram_buffer(77999) := X"00000000";
        ram_buffer(78000) := X"00000000";
        ram_buffer(78001) := X"00000000";
        ram_buffer(78002) := X"00000000";
        ram_buffer(78003) := X"00000000";
        ram_buffer(78004) := X"00000000";
        ram_buffer(78005) := X"00000000";
        ram_buffer(78006) := X"00000000";
        ram_buffer(78007) := X"00000000";
        ram_buffer(78008) := X"00000000";
        ram_buffer(78009) := X"00000000";
        ram_buffer(78010) := X"00000000";
        ram_buffer(78011) := X"00000000";
        ram_buffer(78012) := X"00000000";
        ram_buffer(78013) := X"00000000";
        ram_buffer(78014) := X"00000000";
        ram_buffer(78015) := X"00000000";
        ram_buffer(78016) := X"00000000";
        ram_buffer(78017) := X"00000000";
        ram_buffer(78018) := X"00000000";
        ram_buffer(78019) := X"00000000";
        ram_buffer(78020) := X"00000000";
        ram_buffer(78021) := X"00000000";
        ram_buffer(78022) := X"00000000";
        ram_buffer(78023) := X"00000000";
        ram_buffer(78024) := X"00000000";
        ram_buffer(78025) := X"00000000";
        ram_buffer(78026) := X"00000000";
        ram_buffer(78027) := X"00000000";
        ram_buffer(78028) := X"00000000";
        ram_buffer(78029) := X"00000000";
        ram_buffer(78030) := X"00000000";
        ram_buffer(78031) := X"00000000";
        ram_buffer(78032) := X"00000000";
        ram_buffer(78033) := X"00000000";
        ram_buffer(78034) := X"00000000";
        ram_buffer(78035) := X"00000000";
        ram_buffer(78036) := X"00000000";
        ram_buffer(78037) := X"00000000";
        ram_buffer(78038) := X"00000000";
        ram_buffer(78039) := X"00000000";
        ram_buffer(78040) := X"00000000";
        ram_buffer(78041) := X"00000000";
        ram_buffer(78042) := X"00000000";
        ram_buffer(78043) := X"00000000";
        ram_buffer(78044) := X"00000000";
        ram_buffer(78045) := X"00000000";
        ram_buffer(78046) := X"00000000";
        ram_buffer(78047) := X"00000000";
        ram_buffer(78048) := X"00000000";
        ram_buffer(78049) := X"00000000";
        ram_buffer(78050) := X"00000000";
        ram_buffer(78051) := X"00000000";
        ram_buffer(78052) := X"00000000";
        ram_buffer(78053) := X"00000000";
        ram_buffer(78054) := X"00000000";
        ram_buffer(78055) := X"00000000";
        ram_buffer(78056) := X"00000000";
        ram_buffer(78057) := X"00000000";
        ram_buffer(78058) := X"00000000";
        ram_buffer(78059) := X"00000000";
        ram_buffer(78060) := X"00000000";
        ram_buffer(78061) := X"00000000";
        ram_buffer(78062) := X"00000000";
        ram_buffer(78063) := X"00000000";
        ram_buffer(78064) := X"00000000";
        ram_buffer(78065) := X"00000000";
        ram_buffer(78066) := X"00000000";
        ram_buffer(78067) := X"00000000";
        ram_buffer(78068) := X"00000000";
        ram_buffer(78069) := X"00000000";
        ram_buffer(78070) := X"00000000";
        ram_buffer(78071) := X"00000000";
        ram_buffer(78072) := X"00000000";
        ram_buffer(78073) := X"00000000";
        ram_buffer(78074) := X"00000000";
        ram_buffer(78075) := X"00000000";
        ram_buffer(78076) := X"00000000";
        ram_buffer(78077) := X"00000000";
        ram_buffer(78078) := X"00000000";
        ram_buffer(78079) := X"00000000";
        ram_buffer(78080) := X"00000000";
        ram_buffer(78081) := X"00000000";
        ram_buffer(78082) := X"00000000";
        ram_buffer(78083) := X"00000000";
        ram_buffer(78084) := X"00000000";
        ram_buffer(78085) := X"00000000";
        ram_buffer(78086) := X"00000000";
        ram_buffer(78087) := X"00000000";
        ram_buffer(78088) := X"00000000";
        ram_buffer(78089) := X"00000000";
        ram_buffer(78090) := X"00000000";
        ram_buffer(78091) := X"00000000";
        ram_buffer(78092) := X"00000000";
        ram_buffer(78093) := X"00000000";
        ram_buffer(78094) := X"00000000";
        ram_buffer(78095) := X"00000000";
        ram_buffer(78096) := X"00000000";
        ram_buffer(78097) := X"00000000";
        ram_buffer(78098) := X"00000000";
        ram_buffer(78099) := X"00000000";
        ram_buffer(78100) := X"00000000";
        ram_buffer(78101) := X"00000000";
        ram_buffer(78102) := X"00000000";
        ram_buffer(78103) := X"00000000";
        ram_buffer(78104) := X"00000000";
        ram_buffer(78105) := X"00000000";
        ram_buffer(78106) := X"00000000";
        ram_buffer(78107) := X"00000000";
        ram_buffer(78108) := X"00000000";
        ram_buffer(78109) := X"00000000";
        ram_buffer(78110) := X"00000000";
        ram_buffer(78111) := X"00000000";
        ram_buffer(78112) := X"00000000";
        ram_buffer(78113) := X"00000000";
        ram_buffer(78114) := X"00000000";
        ram_buffer(78115) := X"00000000";
        ram_buffer(78116) := X"00000000";
        ram_buffer(78117) := X"00000000";
        ram_buffer(78118) := X"00000000";
        ram_buffer(78119) := X"00000000";
        ram_buffer(78120) := X"00000000";
        ram_buffer(78121) := X"00000000";
        ram_buffer(78122) := X"00000000";
        ram_buffer(78123) := X"00000000";
        ram_buffer(78124) := X"00000000";
        ram_buffer(78125) := X"00000000";
        ram_buffer(78126) := X"00000000";
        ram_buffer(78127) := X"00000000";
        ram_buffer(78128) := X"00000000";
        ram_buffer(78129) := X"00000000";
        ram_buffer(78130) := X"00000000";
        ram_buffer(78131) := X"00000000";
        ram_buffer(78132) := X"00000000";
        ram_buffer(78133) := X"00000000";
        ram_buffer(78134) := X"00000000";
        ram_buffer(78135) := X"00000000";
        ram_buffer(78136) := X"00000000";
        ram_buffer(78137) := X"00000000";
        ram_buffer(78138) := X"00000000";
        ram_buffer(78139) := X"00000000";
        ram_buffer(78140) := X"00000000";
        ram_buffer(78141) := X"00000000";
        ram_buffer(78142) := X"00000000";
        ram_buffer(78143) := X"00000000";
        ram_buffer(78144) := X"00000000";
        ram_buffer(78145) := X"00000000";
        ram_buffer(78146) := X"00000000";
        ram_buffer(78147) := X"00000000";
        ram_buffer(78148) := X"00000000";
        ram_buffer(78149) := X"00000000";
        ram_buffer(78150) := X"00000000";
        ram_buffer(78151) := X"00000000";
        ram_buffer(78152) := X"00000000";
        ram_buffer(78153) := X"00000000";
        ram_buffer(78154) := X"00000000";
        ram_buffer(78155) := X"00000000";
        ram_buffer(78156) := X"00000000";
        ram_buffer(78157) := X"00000000";
        ram_buffer(78158) := X"00000000";
        ram_buffer(78159) := X"00000000";
        ram_buffer(78160) := X"00000000";
        ram_buffer(78161) := X"00000000";
        ram_buffer(78162) := X"00000000";
        ram_buffer(78163) := X"00000000";
        ram_buffer(78164) := X"00000000";
        ram_buffer(78165) := X"00000000";
        ram_buffer(78166) := X"00000000";
        ram_buffer(78167) := X"00000000";
        ram_buffer(78168) := X"00000000";
        ram_buffer(78169) := X"00000000";
        ram_buffer(78170) := X"00000000";
        ram_buffer(78171) := X"00000000";
        ram_buffer(78172) := X"00000000";
        ram_buffer(78173) := X"00000000";
        ram_buffer(78174) := X"00000000";
        ram_buffer(78175) := X"00000000";
        ram_buffer(78176) := X"00000000";
        ram_buffer(78177) := X"00000000";
        ram_buffer(78178) := X"00000000";
        ram_buffer(78179) := X"00000000";
        ram_buffer(78180) := X"00000000";
        ram_buffer(78181) := X"00000000";
        ram_buffer(78182) := X"00000000";
        ram_buffer(78183) := X"00000000";
        ram_buffer(78184) := X"00000000";
        ram_buffer(78185) := X"00000000";
        ram_buffer(78186) := X"00000000";
        ram_buffer(78187) := X"00000000";
        ram_buffer(78188) := X"00000000";
        ram_buffer(78189) := X"00000000";
        ram_buffer(78190) := X"00000000";
        ram_buffer(78191) := X"00000000";
        ram_buffer(78192) := X"00000000";
        ram_buffer(78193) := X"00000000";
        ram_buffer(78194) := X"00000000";
        ram_buffer(78195) := X"00000000";
        ram_buffer(78196) := X"00000000";
        ram_buffer(78197) := X"00000000";
        ram_buffer(78198) := X"00000000";
        ram_buffer(78199) := X"00000000";
        ram_buffer(78200) := X"00000000";
        ram_buffer(78201) := X"00000000";
        ram_buffer(78202) := X"00000000";
        ram_buffer(78203) := X"00000000";
        ram_buffer(78204) := X"00000000";
        ram_buffer(78205) := X"00000000";
        ram_buffer(78206) := X"00000000";
        ram_buffer(78207) := X"00000000";
        ram_buffer(78208) := X"00000000";
        ram_buffer(78209) := X"00000000";
        ram_buffer(78210) := X"00000000";
        ram_buffer(78211) := X"00000000";
        ram_buffer(78212) := X"00000000";
        ram_buffer(78213) := X"00000000";
        ram_buffer(78214) := X"00000000";
        ram_buffer(78215) := X"00000000";
        ram_buffer(78216) := X"00000000";
        ram_buffer(78217) := X"00000000";
        ram_buffer(78218) := X"00000000";
        ram_buffer(78219) := X"00000000";
        ram_buffer(78220) := X"00000000";
        ram_buffer(78221) := X"00000000";
        ram_buffer(78222) := X"00000000";
        ram_buffer(78223) := X"00000000";
        ram_buffer(78224) := X"00000000";
        ram_buffer(78225) := X"00000000";
        ram_buffer(78226) := X"00000000";
        ram_buffer(78227) := X"00000000";
        ram_buffer(78228) := X"00000000";
        ram_buffer(78229) := X"00000000";
        ram_buffer(78230) := X"00000000";
        ram_buffer(78231) := X"00000000";
        ram_buffer(78232) := X"00000000";
        ram_buffer(78233) := X"00000000";
        ram_buffer(78234) := X"00000000";
        ram_buffer(78235) := X"00000000";
        ram_buffer(78236) := X"00000000";
        ram_buffer(78237) := X"00000000";
        ram_buffer(78238) := X"00000000";
        ram_buffer(78239) := X"00000000";
        ram_buffer(78240) := X"00000000";
        ram_buffer(78241) := X"00000000";
        ram_buffer(78242) := X"00000000";
        ram_buffer(78243) := X"00000000";
        ram_buffer(78244) := X"00000000";
        ram_buffer(78245) := X"00000000";
        ram_buffer(78246) := X"00000000";
        ram_buffer(78247) := X"00000000";
        ram_buffer(78248) := X"00000000";
        ram_buffer(78249) := X"00000000";
        ram_buffer(78250) := X"00000000";
        ram_buffer(78251) := X"00000000";
        ram_buffer(78252) := X"00000000";
        ram_buffer(78253) := X"00000000";
        ram_buffer(78254) := X"00000000";
        ram_buffer(78255) := X"00000000";
        ram_buffer(78256) := X"00000000";
        ram_buffer(78257) := X"00000000";
        ram_buffer(78258) := X"00000000";
        ram_buffer(78259) := X"00000000";
        ram_buffer(78260) := X"00000000";
        ram_buffer(78261) := X"00000000";
        ram_buffer(78262) := X"00000000";
        ram_buffer(78263) := X"00000000";
        ram_buffer(78264) := X"00000000";
        ram_buffer(78265) := X"00000000";
        ram_buffer(78266) := X"00000000";
        ram_buffer(78267) := X"00000000";
        ram_buffer(78268) := X"00000000";
        ram_buffer(78269) := X"00000000";
        ram_buffer(78270) := X"00000000";
        ram_buffer(78271) := X"00000000";
        ram_buffer(78272) := X"00000000";
        ram_buffer(78273) := X"00000000";
        ram_buffer(78274) := X"00000000";
        ram_buffer(78275) := X"00000000";
        ram_buffer(78276) := X"00000000";
        ram_buffer(78277) := X"00000000";
        ram_buffer(78278) := X"00000000";
        ram_buffer(78279) := X"00000000";
        ram_buffer(78280) := X"00000000";
        ram_buffer(78281) := X"00000000";
        ram_buffer(78282) := X"00000000";
        ram_buffer(78283) := X"00000000";
        ram_buffer(78284) := X"00000000";
        ram_buffer(78285) := X"00000000";
        ram_buffer(78286) := X"00000000";
        ram_buffer(78287) := X"00000000";
        ram_buffer(78288) := X"00000000";
        ram_buffer(78289) := X"00000000";
        ram_buffer(78290) := X"00000000";
        ram_buffer(78291) := X"00000000";
        ram_buffer(78292) := X"00000000";
        ram_buffer(78293) := X"00000000";
        ram_buffer(78294) := X"00000000";
        ram_buffer(78295) := X"00000000";
        ram_buffer(78296) := X"00000000";
        ram_buffer(78297) := X"00000000";
        ram_buffer(78298) := X"00000000";
        ram_buffer(78299) := X"00000000";
        ram_buffer(78300) := X"00000000";
        ram_buffer(78301) := X"00000000";
        ram_buffer(78302) := X"00000000";
        ram_buffer(78303) := X"00000000";
        ram_buffer(78304) := X"00000000";
        ram_buffer(78305) := X"00000000";
        ram_buffer(78306) := X"00000000";
        ram_buffer(78307) := X"00000000";
        ram_buffer(78308) := X"00000000";
        ram_buffer(78309) := X"00000000";
        ram_buffer(78310) := X"00000000";
        ram_buffer(78311) := X"00000000";
        ram_buffer(78312) := X"FFFFFFFF";
        ram_buffer(78313) := X"00000000";
        ram_buffer(78314) := X"FFFFFFFF";
        ram_buffer(78315) := X"00000000";
        ram_buffer(78316) := X"00000000";
        ram_buffer(78317) := X"00000000";
        ram_buffer(78318) := X"00000000";
        ram_buffer(78319) := X"100CCAA4";
        ram_buffer(78320) := X"100CCB0C";
        ram_buffer(78321) := X"100CCB74";
        ram_buffer(78322) := X"00000000";
        ram_buffer(78323) := X"00000000";
        ram_buffer(78324) := X"00000000";
        ram_buffer(78325) := X"00000000";
        ram_buffer(78326) := X"00000000";
        ram_buffer(78327) := X"00000000";
        ram_buffer(78328) := X"00000000";
        ram_buffer(78329) := X"00000000";
        ram_buffer(78330) := X"00000000";
        ram_buffer(78331) := X"100CA070";
        ram_buffer(78332) := X"00000000";
        ram_buffer(78333) := X"00000000";
        ram_buffer(78334) := X"00000000";
        ram_buffer(78335) := X"00000000";
        ram_buffer(78336) := X"00000000";
        ram_buffer(78337) := X"00000000";
        ram_buffer(78338) := X"00000000";
        ram_buffer(78339) := X"00000000";
        ram_buffer(78340) := X"00000000";
        ram_buffer(78341) := X"00000000";
        ram_buffer(78342) := X"00000000";
        ram_buffer(78343) := X"00000000";
        ram_buffer(78344) := X"00000000";
        ram_buffer(78345) := X"00000000";
        ram_buffer(78346) := X"00000000";
        ram_buffer(78347) := X"00000000";
        ram_buffer(78348) := X"00000000";
        ram_buffer(78349) := X"00000000";
        ram_buffer(78350) := X"00000000";
        ram_buffer(78351) := X"00000000";
        ram_buffer(78352) := X"00000000";
        ram_buffer(78353) := X"00000000";
        ram_buffer(78354) := X"00000000";
        ram_buffer(78355) := X"00000000";
        ram_buffer(78356) := X"00000000";
        ram_buffer(78357) := X"00000000";
        ram_buffer(78358) := X"00000000";
        ram_buffer(78359) := X"00000000";
        ram_buffer(78360) := X"00000000";
        ram_buffer(78361) := X"00000001";
        ram_buffer(78362) := X"330EABCD";
        ram_buffer(78363) := X"1234E66D";
        ram_buffer(78364) := X"DEEC0005";
        ram_buffer(78365) := X"000B0000";
        ram_buffer(78366) := X"00000000";
        ram_buffer(78367) := X"00000000";
        ram_buffer(78368) := X"00000000";
        ram_buffer(78369) := X"00000000";
        ram_buffer(78370) := X"00000000";
        ram_buffer(78371) := X"00000000";
        ram_buffer(78372) := X"00000000";
        ram_buffer(78373) := X"00000000";
        ram_buffer(78374) := X"00000000";
        ram_buffer(78375) := X"00000000";
        ram_buffer(78376) := X"00000000";
        ram_buffer(78377) := X"00000000";
        ram_buffer(78378) := X"00000000";
        ram_buffer(78379) := X"00000000";
        ram_buffer(78380) := X"00000000";
        ram_buffer(78381) := X"00000000";
        ram_buffer(78382) := X"00000000";
        ram_buffer(78383) := X"00000000";
        ram_buffer(78384) := X"00000000";
        ram_buffer(78385) := X"00000000";
        ram_buffer(78386) := X"00000000";
        ram_buffer(78387) := X"00000000";
        ram_buffer(78388) := X"00000000";
        ram_buffer(78389) := X"00000000";
        ram_buffer(78390) := X"00000000";
        ram_buffer(78391) := X"00000000";
        ram_buffer(78392) := X"00000000";
        ram_buffer(78393) := X"00000000";
        ram_buffer(78394) := X"00000000";
        ram_buffer(78395) := X"00000000";
        ram_buffer(78396) := X"00000000";
        ram_buffer(78397) := X"00000000";
        ram_buffer(78398) := X"00000000";
        ram_buffer(78399) := X"00000000";
        ram_buffer(78400) := X"00000000";
        ram_buffer(78401) := X"00000000";
        ram_buffer(78402) := X"00000000";
        ram_buffer(78403) := X"00000000";
        ram_buffer(78404) := X"00000000";
        ram_buffer(78405) := X"00000000";
        ram_buffer(78406) := X"00000000";
        ram_buffer(78407) := X"00000000";
        ram_buffer(78408) := X"00000000";
        ram_buffer(78409) := X"00000000";
        ram_buffer(78410) := X"00000000";
        ram_buffer(78411) := X"00000000";
        ram_buffer(78412) := X"00000000";
        ram_buffer(78413) := X"00000000";
        ram_buffer(78414) := X"00000000";
        ram_buffer(78415) := X"00000000";
        ram_buffer(78416) := X"00000000";
        ram_buffer(78417) := X"00000000";
        ram_buffer(78418) := X"00000000";
        ram_buffer(78419) := X"00000000";
        ram_buffer(78420) := X"00000000";
        ram_buffer(78421) := X"00000000";
        ram_buffer(78422) := X"00000000";
        ram_buffer(78423) := X"00000000";
        ram_buffer(78424) := X"00000000";
        ram_buffer(78425) := X"00000000";
        ram_buffer(78426) := X"00000000";
        ram_buffer(78427) := X"00000000";
        ram_buffer(78428) := X"00000000";
        ram_buffer(78429) := X"00000000";
        ram_buffer(78430) := X"00000000";
        ram_buffer(78431) := X"00000000";
        ram_buffer(78432) := X"00000000";
        ram_buffer(78433) := X"00000000";
        ram_buffer(78434) := X"00000000";
        ram_buffer(78435) := X"00000000";
        ram_buffer(78436) := X"00000000";
        ram_buffer(78437) := X"00000000";
        ram_buffer(78438) := X"00000000";
        ram_buffer(78439) := X"00000000";
        ram_buffer(78440) := X"00000000";
        ram_buffer(78441) := X"00000000";
        ram_buffer(78442) := X"00000000";
        ram_buffer(78443) := X"00000000";
        ram_buffer(78444) := X"00000000";
        ram_buffer(78445) := X"00000000";
        ram_buffer(78446) := X"00000000";
        ram_buffer(78447) := X"00000000";
        ram_buffer(78448) := X"00000000";
        ram_buffer(78449) := X"00000000";
        ram_buffer(78450) := X"00000000";
        ram_buffer(78451) := X"00000000";
        ram_buffer(78452) := X"00000000";
        ram_buffer(78453) := X"00000000";
        ram_buffer(78454) := X"00000000";
        ram_buffer(78455) := X"00000000";
        ram_buffer(78456) := X"00000000";
        ram_buffer(78457) := X"00000000";
        ram_buffer(78458) := X"00000000";
        ram_buffer(78459) := X"00000000";
        ram_buffer(78460) := X"00000000";
        ram_buffer(78461) := X"00000000";
        ram_buffer(78462) := X"00000000";
        ram_buffer(78463) := X"00000000";
        ram_buffer(78464) := X"00000000";
        ram_buffer(78465) := X"00000000";
        ram_buffer(78466) := X"00000000";
        ram_buffer(78467) := X"00000000";
        ram_buffer(78468) := X"00000000";
        ram_buffer(78469) := X"00000000";
        ram_buffer(78470) := X"00000000";
        ram_buffer(78471) := X"00000000";
        ram_buffer(78472) := X"00000000";
        ram_buffer(78473) := X"00000000";
        ram_buffer(78474) := X"00000000";
        ram_buffer(78475) := X"00000000";
        ram_buffer(78476) := X"00000000";
        ram_buffer(78477) := X"00000000";
        ram_buffer(78478) := X"00000000";
        ram_buffer(78479) := X"00000000";
        ram_buffer(78480) := X"00000000";
        ram_buffer(78481) := X"00000000";
        ram_buffer(78482) := X"00000000";
        ram_buffer(78483) := X"00000000";
        ram_buffer(78484) := X"00000000";
        ram_buffer(78485) := X"00000000";
        ram_buffer(78486) := X"00000000";
        ram_buffer(78487) := X"00000000";
        ram_buffer(78488) := X"00000000";
        ram_buffer(78489) := X"00000000";
        ram_buffer(78490) := X"00000000";
        ram_buffer(78491) := X"00000000";
        ram_buffer(78492) := X"00000000";
        ram_buffer(78493) := X"00000000";
        ram_buffer(78494) := X"00000000";
        ram_buffer(78495) := X"00000000";
        ram_buffer(78496) := X"00000000";
        ram_buffer(78497) := X"00000000";
        ram_buffer(78498) := X"00000000";
        ram_buffer(78499) := X"00000000";
        ram_buffer(78500) := X"00000000";
        ram_buffer(78501) := X"00000000";
        ram_buffer(78502) := X"00000000";
        ram_buffer(78503) := X"00000000";
        ram_buffer(78504) := X"00000000";
        ram_buffer(78505) := X"00000000";
        ram_buffer(78506) := X"00000000";
        ram_buffer(78507) := X"00000000";
        ram_buffer(78508) := X"00000000";
        ram_buffer(78509) := X"00000000";
        ram_buffer(78510) := X"00000000";
        ram_buffer(78511) := X"00000000";
        ram_buffer(78512) := X"00000000";
        ram_buffer(78513) := X"00000000";
        ram_buffer(78514) := X"00000000";
        ram_buffer(78515) := X"00000000";
        ram_buffer(78516) := X"00000000";
        ram_buffer(78517) := X"00000000";
        ram_buffer(78518) := X"00000000";
        ram_buffer(78519) := X"00000000";
        ram_buffer(78520) := X"00000000";
        ram_buffer(78521) := X"00000000";
        ram_buffer(78522) := X"00000000";
        ram_buffer(78523) := X"00000000";
        ram_buffer(78524) := X"00000000";
        ram_buffer(78525) := X"00000000";
        ram_buffer(78526) := X"00000000";
        ram_buffer(78527) := X"00000000";
        ram_buffer(78528) := X"00000000";
        ram_buffer(78529) := X"00000000";
        ram_buffer(78530) := X"00000000";
        ram_buffer(78531) := X"00000000";
        ram_buffer(78532) := X"00000000";
        ram_buffer(78533) := X"00000000";
        ram_buffer(78534) := X"00000000";
        ram_buffer(78535) := X"00000000";
        ram_buffer(78536) := X"00000000";
        ram_buffer(78537) := X"00000000";
        ram_buffer(78538) := X"00000000";
        ram_buffer(78539) := X"00000000";
        ram_buffer(78540) := X"00000000";
        ram_buffer(78541) := X"00000000";
        ram_buffer(78542) := X"00000000";
        ram_buffer(78543) := X"00000000";
        ram_buffer(78544) := X"00000000";
        ram_buffer(78545) := X"00000000";
        ram_buffer(78546) := X"00000000";
        ram_buffer(78547) := X"00000000";
        ram_buffer(78548) := X"00000000";
        ram_buffer(78549) := X"00000000";
        ram_buffer(78550) := X"00000000";
        ram_buffer(78551) := X"00000000";
        ram_buffer(78552) := X"00000000";
        ram_buffer(78553) := X"00000000";
        ram_buffer(78554) := X"00000000";
        ram_buffer(78555) := X"00000000";
        ram_buffer(78556) := X"00000000";
        ram_buffer(78557) := X"00000000";
        ram_buffer(78558) := X"00000000";
        ram_buffer(78559) := X"00000000";
        ram_buffer(78560) := X"00000000";
        ram_buffer(78561) := X"00000000";
        ram_buffer(78562) := X"00000000";
        ram_buffer(78563) := X"00000000";
        ram_buffer(78564) := X"00000000";
        ram_buffer(78565) := X"00000000";
        ram_buffer(78566) := X"00000000";
        ram_buffer(78567) := X"00000000";
        ram_buffer(78568) := X"00000000";
        ram_buffer(78569) := X"00000000";
        ram_buffer(78570) := X"00000000";
        ram_buffer(78571) := X"00000000";
        ram_buffer(78572) := X"00000000";
        ram_buffer(78573) := X"00000000";
        ram_buffer(78574) := X"00000000";
        ram_buffer(78575) := X"00000000";
        ram_buffer(78576) := X"00000000";
        ram_buffer(78577) := X"00000000";
        ram_buffer(78578) := X"00000000";
        ram_buffer(78579) := X"00000000";
        ram_buffer(78580) := X"00000000";
        ram_buffer(78581) := X"00000000";
        ram_buffer(78582) := X"00000000";
        ram_buffer(78583) := X"00000000";
        ram_buffer(78584) := X"00000000";
        ram_buffer(78585) := X"00000000";
        ram_buffer(78586) := X"100CCBE0";
        ram_buffer(78587) := X"100CCBE0";
        ram_buffer(78588) := X"100CCBE8";
        ram_buffer(78589) := X"100CCBE8";
        ram_buffer(78590) := X"100CCBF0";
        ram_buffer(78591) := X"100CCBF0";
        ram_buffer(78592) := X"100CCBF8";
        ram_buffer(78593) := X"100CCBF8";
        ram_buffer(78594) := X"100CCC00";
        ram_buffer(78595) := X"100CCC00";
        ram_buffer(78596) := X"100CCC08";
        ram_buffer(78597) := X"100CCC08";
        ram_buffer(78598) := X"100CCC10";
        ram_buffer(78599) := X"100CCC10";
        ram_buffer(78600) := X"100CCC18";
        ram_buffer(78601) := X"100CCC18";
        ram_buffer(78602) := X"100CCC20";
        ram_buffer(78603) := X"100CCC20";
        ram_buffer(78604) := X"100CCC28";
        ram_buffer(78605) := X"100CCC28";
        ram_buffer(78606) := X"100CCC30";
        ram_buffer(78607) := X"100CCC30";
        ram_buffer(78608) := X"100CCC38";
        ram_buffer(78609) := X"100CCC38";
        ram_buffer(78610) := X"100CCC40";
        ram_buffer(78611) := X"100CCC40";
        ram_buffer(78612) := X"100CCC48";
        ram_buffer(78613) := X"100CCC48";
        ram_buffer(78614) := X"100CCC50";
        ram_buffer(78615) := X"100CCC50";
        ram_buffer(78616) := X"100CCC58";
        ram_buffer(78617) := X"100CCC58";
        ram_buffer(78618) := X"100CCC60";
        ram_buffer(78619) := X"100CCC60";
        ram_buffer(78620) := X"100CCC68";
        ram_buffer(78621) := X"100CCC68";
        ram_buffer(78622) := X"100CCC70";
        ram_buffer(78623) := X"100CCC70";
        ram_buffer(78624) := X"100CCC78";
        ram_buffer(78625) := X"100CCC78";
        ram_buffer(78626) := X"100CCC80";
        ram_buffer(78627) := X"100CCC80";
        ram_buffer(78628) := X"100CCC88";
        ram_buffer(78629) := X"100CCC88";
        ram_buffer(78630) := X"100CCC90";
        ram_buffer(78631) := X"100CCC90";
        ram_buffer(78632) := X"100CCC98";
        ram_buffer(78633) := X"100CCC98";
        ram_buffer(78634) := X"100CCCA0";
        ram_buffer(78635) := X"100CCCA0";
        ram_buffer(78636) := X"100CCCA8";
        ram_buffer(78637) := X"100CCCA8";
        ram_buffer(78638) := X"100CCCB0";
        ram_buffer(78639) := X"100CCCB0";
        ram_buffer(78640) := X"100CCCB8";
        ram_buffer(78641) := X"100CCCB8";
        ram_buffer(78642) := X"100CCCC0";
        ram_buffer(78643) := X"100CCCC0";
        ram_buffer(78644) := X"100CCCC8";
        ram_buffer(78645) := X"100CCCC8";
        ram_buffer(78646) := X"100CCCD0";
        ram_buffer(78647) := X"100CCCD0";
        ram_buffer(78648) := X"100CCCD8";
        ram_buffer(78649) := X"100CCCD8";
        ram_buffer(78650) := X"100CCCE0";
        ram_buffer(78651) := X"100CCCE0";
        ram_buffer(78652) := X"100CCCE8";
        ram_buffer(78653) := X"100CCCE8";
        ram_buffer(78654) := X"100CCCF0";
        ram_buffer(78655) := X"100CCCF0";
        ram_buffer(78656) := X"100CCCF8";
        ram_buffer(78657) := X"100CCCF8";
        ram_buffer(78658) := X"100CCD00";
        ram_buffer(78659) := X"100CCD00";
        ram_buffer(78660) := X"100CCD08";
        ram_buffer(78661) := X"100CCD08";
        ram_buffer(78662) := X"100CCD10";
        ram_buffer(78663) := X"100CCD10";
        ram_buffer(78664) := X"100CCD18";
        ram_buffer(78665) := X"100CCD18";
        ram_buffer(78666) := X"100CCD20";
        ram_buffer(78667) := X"100CCD20";
        ram_buffer(78668) := X"100CCD28";
        ram_buffer(78669) := X"100CCD28";
        ram_buffer(78670) := X"100CCD30";
        ram_buffer(78671) := X"100CCD30";
        ram_buffer(78672) := X"100CCD38";
        ram_buffer(78673) := X"100CCD38";
        ram_buffer(78674) := X"100CCD40";
        ram_buffer(78675) := X"100CCD40";
        ram_buffer(78676) := X"100CCD48";
        ram_buffer(78677) := X"100CCD48";
        ram_buffer(78678) := X"100CCD50";
        ram_buffer(78679) := X"100CCD50";
        ram_buffer(78680) := X"100CCD58";
        ram_buffer(78681) := X"100CCD58";
        ram_buffer(78682) := X"100CCD60";
        ram_buffer(78683) := X"100CCD60";
        ram_buffer(78684) := X"100CCD68";
        ram_buffer(78685) := X"100CCD68";
        ram_buffer(78686) := X"100CCD70";
        ram_buffer(78687) := X"100CCD70";
        ram_buffer(78688) := X"100CCD78";
        ram_buffer(78689) := X"100CCD78";
        ram_buffer(78690) := X"100CCD80";
        ram_buffer(78691) := X"100CCD80";
        ram_buffer(78692) := X"100CCD88";
        ram_buffer(78693) := X"100CCD88";
        ram_buffer(78694) := X"100CCD90";
        ram_buffer(78695) := X"100CCD90";
        ram_buffer(78696) := X"100CCD98";
        ram_buffer(78697) := X"100CCD98";
        ram_buffer(78698) := X"100CCDA0";
        ram_buffer(78699) := X"100CCDA0";
        ram_buffer(78700) := X"100CCDA8";
        ram_buffer(78701) := X"100CCDA8";
        ram_buffer(78702) := X"100CCDB0";
        ram_buffer(78703) := X"100CCDB0";
        ram_buffer(78704) := X"100CCDB8";
        ram_buffer(78705) := X"100CCDB8";
        ram_buffer(78706) := X"100CCDC0";
        ram_buffer(78707) := X"100CCDC0";
        ram_buffer(78708) := X"100CCDC8";
        ram_buffer(78709) := X"100CCDC8";
        ram_buffer(78710) := X"100CCDD0";
        ram_buffer(78711) := X"100CCDD0";
        ram_buffer(78712) := X"100CCDD8";
        ram_buffer(78713) := X"100CCDD8";
        ram_buffer(78714) := X"100CCDE0";
        ram_buffer(78715) := X"100CCDE0";
        ram_buffer(78716) := X"100CCDE8";
        ram_buffer(78717) := X"100CCDE8";
        ram_buffer(78718) := X"100CCDF0";
        ram_buffer(78719) := X"100CCDF0";
        ram_buffer(78720) := X"100CCDF8";
        ram_buffer(78721) := X"100CCDF8";
        ram_buffer(78722) := X"100CCE00";
        ram_buffer(78723) := X"100CCE00";
        ram_buffer(78724) := X"100CCE08";
        ram_buffer(78725) := X"100CCE08";
        ram_buffer(78726) := X"100CCE10";
        ram_buffer(78727) := X"100CCE10";
        ram_buffer(78728) := X"100CCE18";
        ram_buffer(78729) := X"100CCE18";
        ram_buffer(78730) := X"100CCE20";
        ram_buffer(78731) := X"100CCE20";
        ram_buffer(78732) := X"100CCE28";
        ram_buffer(78733) := X"100CCE28";
        ram_buffer(78734) := X"100CCE30";
        ram_buffer(78735) := X"100CCE30";
        ram_buffer(78736) := X"100CCE38";
        ram_buffer(78737) := X"100CCE38";
        ram_buffer(78738) := X"100CCE40";
        ram_buffer(78739) := X"100CCE40";
        ram_buffer(78740) := X"100CCE48";
        ram_buffer(78741) := X"100CCE48";
        ram_buffer(78742) := X"100CCE50";
        ram_buffer(78743) := X"100CCE50";
        ram_buffer(78744) := X"100CCE58";
        ram_buffer(78745) := X"100CCE58";
        ram_buffer(78746) := X"100CCE60";
        ram_buffer(78747) := X"100CCE60";
        ram_buffer(78748) := X"100CCE68";
        ram_buffer(78749) := X"100CCE68";
        ram_buffer(78750) := X"100CCE70";
        ram_buffer(78751) := X"100CCE70";
        ram_buffer(78752) := X"100CCE78";
        ram_buffer(78753) := X"100CCE78";
        ram_buffer(78754) := X"100CCE80";
        ram_buffer(78755) := X"100CCE80";
        ram_buffer(78756) := X"100CCE88";
        ram_buffer(78757) := X"100CCE88";
        ram_buffer(78758) := X"100CCE90";
        ram_buffer(78759) := X"100CCE90";
        ram_buffer(78760) := X"100CCE98";
        ram_buffer(78761) := X"100CCE98";
        ram_buffer(78762) := X"100CCEA0";
        ram_buffer(78763) := X"100CCEA0";
        ram_buffer(78764) := X"100CCEA8";
        ram_buffer(78765) := X"100CCEA8";
        ram_buffer(78766) := X"100CCEB0";
        ram_buffer(78767) := X"100CCEB0";
        ram_buffer(78768) := X"100CCEB8";
        ram_buffer(78769) := X"100CCEB8";
        ram_buffer(78770) := X"100CCEC0";
        ram_buffer(78771) := X"100CCEC0";
        ram_buffer(78772) := X"100CCEC8";
        ram_buffer(78773) := X"100CCEC8";
        ram_buffer(78774) := X"100CCED0";
        ram_buffer(78775) := X"100CCED0";
        ram_buffer(78776) := X"100CCED8";
        ram_buffer(78777) := X"100CCED8";
        ram_buffer(78778) := X"100CCEE0";
        ram_buffer(78779) := X"100CCEE0";
        ram_buffer(78780) := X"100CCEE8";
        ram_buffer(78781) := X"100CCEE8";
        ram_buffer(78782) := X"100CCEF0";
        ram_buffer(78783) := X"100CCEF0";
        ram_buffer(78784) := X"100CCEF8";
        ram_buffer(78785) := X"100CCEF8";
        ram_buffer(78786) := X"100CCF00";
        ram_buffer(78787) := X"100CCF00";
        ram_buffer(78788) := X"100CCF08";
        ram_buffer(78789) := X"100CCF08";
        ram_buffer(78790) := X"100CCF10";
        ram_buffer(78791) := X"100CCF10";
        ram_buffer(78792) := X"100CCF18";
        ram_buffer(78793) := X"100CCF18";
        ram_buffer(78794) := X"100CCF20";
        ram_buffer(78795) := X"100CCF20";
        ram_buffer(78796) := X"100CCF28";
        ram_buffer(78797) := X"100CCF28";
        ram_buffer(78798) := X"100CCF30";
        ram_buffer(78799) := X"100CCF30";
        ram_buffer(78800) := X"100CCF38";
        ram_buffer(78801) := X"100CCF38";
        ram_buffer(78802) := X"100CCF40";
        ram_buffer(78803) := X"100CCF40";
        ram_buffer(78804) := X"100CCF48";
        ram_buffer(78805) := X"100CCF48";
        ram_buffer(78806) := X"100CCF50";
        ram_buffer(78807) := X"100CCF50";
        ram_buffer(78808) := X"100CCF58";
        ram_buffer(78809) := X"100CCF58";
        ram_buffer(78810) := X"100CCF60";
        ram_buffer(78811) := X"100CCF60";
        ram_buffer(78812) := X"100CCF68";
        ram_buffer(78813) := X"100CCF68";
        ram_buffer(78814) := X"100CCF70";
        ram_buffer(78815) := X"100CCF70";
        ram_buffer(78816) := X"100CCF78";
        ram_buffer(78817) := X"100CCF78";
        ram_buffer(78818) := X"100CCF80";
        ram_buffer(78819) := X"100CCF80";
        ram_buffer(78820) := X"100CCF88";
        ram_buffer(78821) := X"100CCF88";
        ram_buffer(78822) := X"100CCF90";
        ram_buffer(78823) := X"100CCF90";
        ram_buffer(78824) := X"100CCF98";
        ram_buffer(78825) := X"100CCF98";
        ram_buffer(78826) := X"100CCFA0";
        ram_buffer(78827) := X"100CCFA0";
        ram_buffer(78828) := X"100CCFA8";
        ram_buffer(78829) := X"100CCFA8";
        ram_buffer(78830) := X"100CCFB0";
        ram_buffer(78831) := X"100CCFB0";
        ram_buffer(78832) := X"100CCFB8";
        ram_buffer(78833) := X"100CCFB8";
        ram_buffer(78834) := X"100CCFC0";
        ram_buffer(78835) := X"100CCFC0";
        ram_buffer(78836) := X"100CCFC8";
        ram_buffer(78837) := X"100CCFC8";
        ram_buffer(78838) := X"100CCFD0";
        ram_buffer(78839) := X"100CCFD0";
        ram_buffer(78840) := X"100CCFD8";
        ram_buffer(78841) := X"100CCFD8";
        ram_buffer(78842) := X"100CA91C";
        ram_buffer(78843) := X"100CA920";
        ram_buffer(78844) := X"100CA920";
        ram_buffer(78845) := X"100CA920";
        ram_buffer(78846) := X"100CA920";
        ram_buffer(78847) := X"100CA920";
        ram_buffer(78848) := X"100CA920";
        ram_buffer(78849) := X"100CA920";
        ram_buffer(78850) := X"100CA920";
        ram_buffer(78851) := X"100CA920";
        ram_buffer(78852) := X"7F7F7F7F";
        ram_buffer(78853) := X"7F7F7F7F";
        ram_buffer(78854) := X"7F7F7F7F";
        ram_buffer(78855) := X"7F7F0000";
        ram_buffer(78856) := X"41534349";
        ram_buffer(78857) := X"49000000";
        ram_buffer(78858) := X"00000000";
        ram_buffer(78859) := X"00000000";
        ram_buffer(78860) := X"00000000";
        ram_buffer(78861) := X"00000000";
        ram_buffer(78862) := X"00000000";
        ram_buffer(78863) := X"00000000";
        ram_buffer(78864) := X"41534349";
        ram_buffer(78865) := X"49000000";
        ram_buffer(78866) := X"00000000";
        ram_buffer(78867) := X"00000000";
        ram_buffer(78868) := X"00000000";
        ram_buffer(78869) := X"00000000";
        ram_buffer(78870) := X"00000000";
        ram_buffer(78871) := X"00000000";
        ram_buffer(78872) := X"00000000";
        ram_buffer(78873) := X"00000000";
        ram_buffer(78874) := X"412E8480";
        ram_buffer(78875) := X"00000000";
        ram_buffer(78876) := X"3FF00000";
        ram_buffer(78877) := X"00000000";
        ram_buffer(78878) := X"40200000";
        ram_buffer(78879) := X"00000000";
        ram_buffer(78880) := X"3FF00000";
        ram_buffer(78881) := X"00000000";
        ram_buffer(78882) := X"3FF63150";
        ram_buffer(78883) := X"B14861EF";
        ram_buffer(78884) := X"3FF4E7AE";
        ram_buffer(78885) := X"914D6FCA";
        ram_buffer(78886) := X"3FF2D062";
        ram_buffer(78887) := X"EF6C11AA";
        ram_buffer(78888) := X"3FE92469";
        ram_buffer(78889) := X"C0A7BF3B";
        ram_buffer(78890) := X"3FE1517A";
        ram_buffer(78891) := X"7BC720BB";
        ram_buffer(78892) := X"3FD1A855";
        ram_buffer(78893) := X"DE72AB5D";
        ram_buffer(78894) := X"46800100";
        ram_buffer(78895) := X"00000000";
        ram_buffer(78896) := X"3F3504F3";
        ram_buffer(78897) := X"3EC3EF15";
        ram_buffer(78898) := X"3F0A8BD4";
        ram_buffer(78899) := X"3FA73D75";
        ram_buffer(78900) := X"00000000";
        ram_buffer(78901) := X"00001388";
        ram_buffer(78902) := X"00000640";
        ram_buffer(78903) := X"00003E80";
        ram_buffer(78904) := X"100C9E6B";
        ram_buffer(78905) := X"100CD170";
        ram_buffer(78906) := X"100CC7B8";
        ram_buffer(78907) := X"100CC7B8";
        ram_buffer(78908) := X"00020000";
        ram_buffer(78909) := X"FFFFFFFF";
        ram_buffer(78910) := X"40200000";
        ram_buffer(78911) := X"00000000";
        ram_buffer(78912) := X"40300000";
        ram_buffer(78913) := X"00000000";
        ram_buffer(78914) := X"3FE00000";
        ram_buffer(78915) := X"00000000";
        ram_buffer(78916) := X"40200000";
        ram_buffer(78917) := X"00000000";
        ram_buffer(78918) := X"40300000";
        ram_buffer(78919) := X"00000000";
        ram_buffer(78920) := X"3FE00000";
        ram_buffer(78921) := X"00000000";
        ram_buffer(78922) := X"3FF80000";
        ram_buffer(78923) := X"00000000";
        ram_buffer(78924) := X"3FD287A7";
        ram_buffer(78925) := X"636F4361";
        ram_buffer(78926) := X"3FC68A28";
        ram_buffer(78927) := X"8B60C8B3";
        ram_buffer(78928) := X"3FD34413";
        ram_buffer(78929) := X"509F79FB";
        ram_buffer(78930) := X"3FF00000";
        ram_buffer(78931) := X"00000000";
        ram_buffer(78932) := X"40240000";
        ram_buffer(78933) := X"00000000";
        ram_buffer(78934) := X"401C0000";
        ram_buffer(78935) := X"00000000";
        ram_buffer(78936) := X"40140000";
        ram_buffer(78937) := X"00000000";
        ram_buffer(78938) := X"3FE00000";
        ram_buffer(78939) := X"00000000";
        ram_buffer(78940) := X"100CD218";
        ram_buffer(78941) := X"00000001";
        ram_buffer(78942) := X"100AF070";
        ram_buffer(78943) := X"00000000";
        ram_buffer(78944) := X"3FF00000";
        ram_buffer(78945) := X"00000000";
        ram_buffer(78946) := X"40240000";
        ram_buffer(78947) := X"00000000";
        ram_buffer(78948) := X"43500000";
        ram_buffer(78949) := X"00000000";
        ram_buffer(78950) := X"43500000";
        ram_buffer(78951) := X"00000000";
        ram_buffer(78952) := X"7FBFFFFF";
        ram_buffer(78953) := X"00000000";
        ram_buffer(78954) := X"40000000";
        ram_buffer(78955) := X"00000000";
        ram_buffer(78956) := X"3FF00000";
        ram_buffer(78957) := X"00000000";
        ram_buffer(78958) := X"BFF00000";
        ram_buffer(78959) := X"00000000";
        ram_buffer(78960) := X"3FE00000";
        ram_buffer(78961) := X"00000000";
        ram_buffer(78962) := X"41DFFFFF";
        ram_buffer(78963) := X"FFC00000";
        ram_buffer(78964) := X"3FDFFFFF";
        ram_buffer(78965) := X"94A03595";
        ram_buffer(78966) := X"3FE00000";
        ram_buffer(78967) := X"35AFE535";
        ram_buffer(78968) := X"3FCFFFFF";
        ram_buffer(78969) := X"94A03595";
        ram_buffer(78970) := X"100BECE4";
        return ram_buffer;
    end;
end;
