library ieee;
use ieee.std_logic_1164.all;

package boot_pack_zynq is

    constant cpu_width : integer := 32;
    constant ram_size : integer := 744;
    subtype word_type is std_logic_vector(cpu_width-1 downto 0);
    type ram_type is array(0 to ram_size-1) of word_type;
    function load_hex return ram_type;
end package;

package body boot_pack_zynq is

    function load_hex return ram_type is
        variable ram_buffer : ram_type := (others=>(others=>'0'));
    begin
        ram_buffer(0) := X"3C1C0001";
        ram_buffer(1) := X"279C8B90";
        ram_buffer(2) := X"3C050000";
        ram_buffer(3) := X"24A50BA0";
        ram_buffer(4) := X"3C040000";
        ram_buffer(5) := X"24840DC0";
        ram_buffer(6) := X"3C1D0000";
        ram_buffer(7) := X"27BD0DA8";
        ram_buffer(8) := X"ACA00000";
        ram_buffer(9) := X"00A4182A";
        ram_buffer(10) := X"1460FFFD";
        ram_buffer(11) := X"24A50004";
        ram_buffer(12) := X"0C00024F";
        ram_buffer(13) := X"00000000";
        ram_buffer(14) := X"0800000E";
        ram_buffer(15) := X"23BDFF98";
        ram_buffer(16) := X"AFA10010";
        ram_buffer(17) := X"AFA20014";
        ram_buffer(18) := X"AFA30018";
        ram_buffer(19) := X"AFA4001C";
        ram_buffer(20) := X"AFA50020";
        ram_buffer(21) := X"AFA60024";
        ram_buffer(22) := X"AFA70028";
        ram_buffer(23) := X"AFA8002C";
        ram_buffer(24) := X"AFA90030";
        ram_buffer(25) := X"AFAA0034";
        ram_buffer(26) := X"AFAB0038";
        ram_buffer(27) := X"AFAC003C";
        ram_buffer(28) := X"AFAD0040";
        ram_buffer(29) := X"AFAE0044";
        ram_buffer(30) := X"AFAF0048";
        ram_buffer(31) := X"AFB8004C";
        ram_buffer(32) := X"AFB90050";
        ram_buffer(33) := X"AFBF0054";
        ram_buffer(34) := X"401A7000";
        ram_buffer(35) := X"235AFFFC";
        ram_buffer(36) := X"AFBA0058";
        ram_buffer(37) := X"0000D810";
        ram_buffer(38) := X"AFBB005C";
        ram_buffer(39) := X"0000D812";
        ram_buffer(40) := X"AFBB0060";
        ram_buffer(41) := X"3C062000";
        ram_buffer(42) := X"8CC40020";
        ram_buffer(43) := X"8CC60010";
        ram_buffer(44) := X"00862024";
        ram_buffer(45) := X"0C0002B6";
        ram_buffer(46) := X"23A50000";
        ram_buffer(47) := X"8FA10010";
        ram_buffer(48) := X"8FA20014";
        ram_buffer(49) := X"8FA30018";
        ram_buffer(50) := X"8FA4001C";
        ram_buffer(51) := X"8FA50020";
        ram_buffer(52) := X"8FA60024";
        ram_buffer(53) := X"8FA70028";
        ram_buffer(54) := X"8FA8002C";
        ram_buffer(55) := X"8FA90030";
        ram_buffer(56) := X"8FAA0034";
        ram_buffer(57) := X"8FAB0038";
        ram_buffer(58) := X"8FAC003C";
        ram_buffer(59) := X"8FAD0040";
        ram_buffer(60) := X"8FAE0044";
        ram_buffer(61) := X"8FAF0048";
        ram_buffer(62) := X"8FB8004C";
        ram_buffer(63) := X"8FB90050";
        ram_buffer(64) := X"8FBF0054";
        ram_buffer(65) := X"8FBA0058";
        ram_buffer(66) := X"8FBB005C";
        ram_buffer(67) := X"03600011";
        ram_buffer(68) := X"8FBB0060";
        ram_buffer(69) := X"03600013";
        ram_buffer(70) := X"23BD0068";
        ram_buffer(71) := X"341B0001";
        ram_buffer(72) := X"03400008";
        ram_buffer(73) := X"409B6000";
        ram_buffer(74) := X"40026000";
        ram_buffer(75) := X"03E00008";
        ram_buffer(76) := X"40846000";
        ram_buffer(77) := X"3C050000";
        ram_buffer(78) := X"24A50160";
        ram_buffer(79) := X"8CA60000";
        ram_buffer(80) := X"AC06003C";
        ram_buffer(81) := X"8CA60004";
        ram_buffer(82) := X"AC060040";
        ram_buffer(83) := X"8CA60008";
        ram_buffer(84) := X"AC060044";
        ram_buffer(85) := X"8CA6000C";
        ram_buffer(86) := X"03E00008";
        ram_buffer(87) := X"AC060048";
        ram_buffer(88) := X"3C1A1000";
        ram_buffer(89) := X"375A003C";
        ram_buffer(90) := X"03400008";
        ram_buffer(91) := X"00000000";
        ram_buffer(92) := X"AC900000";
        ram_buffer(93) := X"AC910004";
        ram_buffer(94) := X"AC920008";
        ram_buffer(95) := X"AC93000C";
        ram_buffer(96) := X"AC940010";
        ram_buffer(97) := X"AC950014";
        ram_buffer(98) := X"AC960018";
        ram_buffer(99) := X"AC97001C";
        ram_buffer(100) := X"AC9E0020";
        ram_buffer(101) := X"AC9C0024";
        ram_buffer(102) := X"AC9D0028";
        ram_buffer(103) := X"AC9F002C";
        ram_buffer(104) := X"03E00008";
        ram_buffer(105) := X"34020000";
        ram_buffer(106) := X"8C900000";
        ram_buffer(107) := X"8C910004";
        ram_buffer(108) := X"8C920008";
        ram_buffer(109) := X"8C93000C";
        ram_buffer(110) := X"8C940010";
        ram_buffer(111) := X"8C950014";
        ram_buffer(112) := X"8C960018";
        ram_buffer(113) := X"8C97001C";
        ram_buffer(114) := X"8C9E0020";
        ram_buffer(115) := X"8C9C0024";
        ram_buffer(116) := X"8C9D0028";
        ram_buffer(117) := X"8C9F002C";
        ram_buffer(118) := X"03E00008";
        ram_buffer(119) := X"34A20000";
        ram_buffer(120) := X"00850019";
        ram_buffer(121) := X"00001012";
        ram_buffer(122) := X"00002010";
        ram_buffer(123) := X"03E00008";
        ram_buffer(124) := X"ACC40000";
        ram_buffer(125) := X"0000000C";
        ram_buffer(126) := X"03E00008";
        ram_buffer(127) := X"00000000";
        ram_buffer(128) := X"27BDFFE8";
        ram_buffer(129) := X"AFBE0014";
        ram_buffer(130) := X"03A0F021";
        ram_buffer(131) := X"3C042000";
        ram_buffer(132) := X"34840068";
        ram_buffer(133) := X"8C840000";
        ram_buffer(134) := X"00000000";
        ram_buffer(135) := X"AFC40004";
        ram_buffer(136) := X"AFC00000";
        ram_buffer(137) := X"3C042000";
        ram_buffer(138) := X"34840060";
        ram_buffer(139) := X"8C840000";
        ram_buffer(140) := X"00000000";
        ram_buffer(141) := X"AFC4000C";
        ram_buffer(142) := X"AFC00008";
        ram_buffer(143) := X"8FC4000C";
        ram_buffer(144) := X"00000000";
        ram_buffer(145) := X"00042000";
        ram_buffer(146) := X"AFC40008";
        ram_buffer(147) := X"AFC0000C";
        ram_buffer(148) := X"8FC4000C";
        ram_buffer(149) := X"00000000";
        ram_buffer(150) := X"00041000";
        ram_buffer(151) := X"00001821";
        ram_buffer(152) := X"8FC40000";
        ram_buffer(153) := X"00000000";
        ram_buffer(154) := X"00822025";
        ram_buffer(155) := X"AFC40000";
        ram_buffer(156) := X"8FC40004";
        ram_buffer(157) := X"00000000";
        ram_buffer(158) := X"00831025";
        ram_buffer(159) := X"AFC20004";
        ram_buffer(160) := X"8FC30004";
        ram_buffer(161) := X"8FC20000";
        ram_buffer(162) := X"03C0E821";
        ram_buffer(163) := X"8FBE0014";
        ram_buffer(164) := X"27BD0018";
        ram_buffer(165) := X"03E00008";
        ram_buffer(166) := X"00000000";
        ram_buffer(167) := X"27BDFFF0";
        ram_buffer(168) := X"AFBE000C";
        ram_buffer(169) := X"03A0F021";
        ram_buffer(170) := X"AFC40010";
        ram_buffer(171) := X"3C020000";
        ram_buffer(172) := X"24420BB0";
        ram_buffer(173) := X"A0400008";
        ram_buffer(174) := X"24020007";
        ram_buffer(175) := X"AFC20000";
        ram_buffer(176) := X"10000024";
        ram_buffer(177) := X"00000000";
        ram_buffer(178) := X"8FC20010";
        ram_buffer(179) := X"00000000";
        ram_buffer(180) := X"00021600";
        ram_buffer(181) := X"00021603";
        ram_buffer(182) := X"3042000F";
        ram_buffer(183) := X"A3C20004";
        ram_buffer(184) := X"83C20004";
        ram_buffer(185) := X"00000000";
        ram_buffer(186) := X"2842000A";
        ram_buffer(187) := X"10400004";
        ram_buffer(188) := X"00000000";
        ram_buffer(189) := X"24020030";
        ram_buffer(190) := X"10000002";
        ram_buffer(191) := X"00000000";
        ram_buffer(192) := X"24020037";
        ram_buffer(193) := X"93C30004";
        ram_buffer(194) := X"00000000";
        ram_buffer(195) := X"00431021";
        ram_buffer(196) := X"304200FF";
        ram_buffer(197) := X"00021E00";
        ram_buffer(198) := X"00031E03";
        ram_buffer(199) := X"3C020000";
        ram_buffer(200) := X"24440BB0";
        ram_buffer(201) := X"8FC20000";
        ram_buffer(202) := X"00000000";
        ram_buffer(203) := X"00821021";
        ram_buffer(204) := X"A0430000";
        ram_buffer(205) := X"8FC20010";
        ram_buffer(206) := X"00000000";
        ram_buffer(207) := X"00021102";
        ram_buffer(208) := X"AFC20010";
        ram_buffer(209) := X"8FC20000";
        ram_buffer(210) := X"00000000";
        ram_buffer(211) := X"2442FFFF";
        ram_buffer(212) := X"AFC20000";
        ram_buffer(213) := X"8FC20000";
        ram_buffer(214) := X"00000000";
        ram_buffer(215) := X"0441FFDA";
        ram_buffer(216) := X"00000000";
        ram_buffer(217) := X"3C020000";
        ram_buffer(218) := X"24420BB0";
        ram_buffer(219) := X"03C0E821";
        ram_buffer(220) := X"8FBE000C";
        ram_buffer(221) := X"27BD0010";
        ram_buffer(222) := X"03E00008";
        ram_buffer(223) := X"00000000";
        ram_buffer(224) := X"27BDFFD8";
        ram_buffer(225) := X"AFBF0024";
        ram_buffer(226) := X"AFBE0020";
        ram_buffer(227) := X"03A0F021";
        ram_buffer(228) := X"AFC00018";
        ram_buffer(229) := X"AFC00010";
        ram_buffer(230) := X"1000006E";
        ram_buffer(231) := X"00000000";
        ram_buffer(232) := X"0C0002C3";
        ram_buffer(233) := X"00000000";
        ram_buffer(234) := X"AFC2001C";
        ram_buffer(235) := X"8FC2001C";
        ram_buffer(236) := X"00000000";
        ram_buffer(237) := X"AFC20014";
        ram_buffer(238) := X"8FC30014";
        ram_buffer(239) := X"2402000A";
        ram_buffer(240) := X"10620069";
        ram_buffer(241) := X"00000000";
        ram_buffer(242) := X"8FC30014";
        ram_buffer(243) := X"2402000D";
        ram_buffer(244) := X"10620065";
        ram_buffer(245) := X"00000000";
        ram_buffer(246) := X"8FC20014";
        ram_buffer(247) := X"00000000";
        ram_buffer(248) := X"2C420030";
        ram_buffer(249) := X"1440000C";
        ram_buffer(250) := X"00000000";
        ram_buffer(251) := X"8FC20014";
        ram_buffer(252) := X"00000000";
        ram_buffer(253) := X"2C42003A";
        ram_buffer(254) := X"10400007";
        ram_buffer(255) := X"00000000";
        ram_buffer(256) := X"8FC20014";
        ram_buffer(257) := X"00000000";
        ram_buffer(258) := X"2442FFD0";
        ram_buffer(259) := X"AFC20014";
        ram_buffer(260) := X"10000040";
        ram_buffer(261) := X"00000000";
        ram_buffer(262) := X"8FC20014";
        ram_buffer(263) := X"00000000";
        ram_buffer(264) := X"2C420041";
        ram_buffer(265) := X"1440000C";
        ram_buffer(266) := X"00000000";
        ram_buffer(267) := X"8FC20014";
        ram_buffer(268) := X"00000000";
        ram_buffer(269) := X"2C42005B";
        ram_buffer(270) := X"10400007";
        ram_buffer(271) := X"00000000";
        ram_buffer(272) := X"8FC20014";
        ram_buffer(273) := X"00000000";
        ram_buffer(274) := X"2442FFC9";
        ram_buffer(275) := X"AFC20014";
        ram_buffer(276) := X"10000030";
        ram_buffer(277) := X"00000000";
        ram_buffer(278) := X"8FC20014";
        ram_buffer(279) := X"00000000";
        ram_buffer(280) := X"2C420061";
        ram_buffer(281) := X"1440000C";
        ram_buffer(282) := X"00000000";
        ram_buffer(283) := X"8FC20014";
        ram_buffer(284) := X"00000000";
        ram_buffer(285) := X"2C42007B";
        ram_buffer(286) := X"10400007";
        ram_buffer(287) := X"00000000";
        ram_buffer(288) := X"8FC20014";
        ram_buffer(289) := X"00000000";
        ram_buffer(290) := X"2442FFA9";
        ram_buffer(291) := X"AFC20014";
        ram_buffer(292) := X"10000020";
        ram_buffer(293) := X"00000000";
        ram_buffer(294) := X"8FC30014";
        ram_buffer(295) := X"24020008";
        ram_buffer(296) := X"1462001C";
        ram_buffer(297) := X"00000000";
        ram_buffer(298) := X"8FC20010";
        ram_buffer(299) := X"00000000";
        ram_buffer(300) := X"18400012";
        ram_buffer(301) := X"00000000";
        ram_buffer(302) := X"8FC20010";
        ram_buffer(303) := X"00000000";
        ram_buffer(304) := X"2442FFFF";
        ram_buffer(305) := X"AFC20010";
        ram_buffer(306) := X"8FC20014";
        ram_buffer(307) := X"00000000";
        ram_buffer(308) := X"00402021";
        ram_buffer(309) := X"0C00026E";
        ram_buffer(310) := X"00000000";
        ram_buffer(311) := X"24040020";
        ram_buffer(312) := X"0C00026E";
        ram_buffer(313) := X"00000000";
        ram_buffer(314) := X"8FC20014";
        ram_buffer(315) := X"00000000";
        ram_buffer(316) := X"00402021";
        ram_buffer(317) := X"0C00026E";
        ram_buffer(318) := X"00000000";
        ram_buffer(319) := X"8FC20018";
        ram_buffer(320) := X"00000000";
        ram_buffer(321) := X"00021102";
        ram_buffer(322) := X"AFC20018";
        ram_buffer(323) := X"10000011";
        ram_buffer(324) := X"00000000";
        ram_buffer(325) := X"8FC2001C";
        ram_buffer(326) := X"00000000";
        ram_buffer(327) := X"00402021";
        ram_buffer(328) := X"0C00026E";
        ram_buffer(329) := X"00000000";
        ram_buffer(330) := X"8FC20018";
        ram_buffer(331) := X"00000000";
        ram_buffer(332) := X"00021900";
        ram_buffer(333) := X"8FC20014";
        ram_buffer(334) := X"00000000";
        ram_buffer(335) := X"00621021";
        ram_buffer(336) := X"AFC20018";
        ram_buffer(337) := X"8FC20010";
        ram_buffer(338) := X"00000000";
        ram_buffer(339) := X"24420001";
        ram_buffer(340) := X"AFC20010";
        ram_buffer(341) := X"8FC20010";
        ram_buffer(342) := X"00000000";
        ram_buffer(343) := X"28420010";
        ram_buffer(344) := X"1440FF8F";
        ram_buffer(345) := X"00000000";
        ram_buffer(346) := X"2404000D";
        ram_buffer(347) := X"0C00026E";
        ram_buffer(348) := X"00000000";
        ram_buffer(349) := X"2404000A";
        ram_buffer(350) := X"0C00026E";
        ram_buffer(351) := X"00000000";
        ram_buffer(352) := X"8FC20018";
        ram_buffer(353) := X"03C0E821";
        ram_buffer(354) := X"8FBF0024";
        ram_buffer(355) := X"8FBE0020";
        ram_buffer(356) := X"27BD0028";
        ram_buffer(357) := X"03E00008";
        ram_buffer(358) := X"00000000";
        ram_buffer(359) := X"27BDFFE0";
        ram_buffer(360) := X"AFBF001C";
        ram_buffer(361) := X"AFBE0018";
        ram_buffer(362) := X"03A0F021";
        ram_buffer(363) := X"AFC40020";
        ram_buffer(364) := X"AFC00010";
        ram_buffer(365) := X"1000002A";
        ram_buffer(366) := X"00000000";
        ram_buffer(367) := X"8FC20010";
        ram_buffer(368) := X"8FC30020";
        ram_buffer(369) := X"00000000";
        ram_buffer(370) := X"00621021";
        ram_buffer(371) := X"8F838010";
        ram_buffer(372) := X"00000000";
        ram_buffer(373) := X"306300FF";
        ram_buffer(374) := X"A0430000";
        ram_buffer(375) := X"AFC00014";
        ram_buffer(376) := X"10000009";
        ram_buffer(377) := X"00000000";
        ram_buffer(378) := X"0C0002BF";
        ram_buffer(379) := X"00000000";
        ram_buffer(380) := X"1440000D";
        ram_buffer(381) := X"00000000";
        ram_buffer(382) := X"8FC20014";
        ram_buffer(383) := X"00000000";
        ram_buffer(384) := X"24420001";
        ram_buffer(385) := X"AFC20014";
        ram_buffer(386) := X"8FC30014";
        ram_buffer(387) := X"3C020001";
        ram_buffer(388) := X"344286A0";
        ram_buffer(389) := X"0062102A";
        ram_buffer(390) := X"1440FFF3";
        ram_buffer(391) := X"00000000";
        ram_buffer(392) := X"10000002";
        ram_buffer(393) := X"00000000";
        ram_buffer(394) := X"00000000";
        ram_buffer(395) := X"8FC30014";
        ram_buffer(396) := X"3C020001";
        ram_buffer(397) := X"344286A0";
        ram_buffer(398) := X"0062102A";
        ram_buffer(399) := X"1040000F";
        ram_buffer(400) := X"00000000";
        ram_buffer(401) := X"0C0002C3";
        ram_buffer(402) := X"00000000";
        ram_buffer(403) := X"AF828010";
        ram_buffer(404) := X"8FC20010";
        ram_buffer(405) := X"00000000";
        ram_buffer(406) := X"24420001";
        ram_buffer(407) := X"AFC20010";
        ram_buffer(408) := X"8FC30010";
        ram_buffer(409) := X"3C020020";
        ram_buffer(410) := X"0062102A";
        ram_buffer(411) := X"1440FFD3";
        ram_buffer(412) := X"00000000";
        ram_buffer(413) := X"10000002";
        ram_buffer(414) := X"00000000";
        ram_buffer(415) := X"00000000";
        ram_buffer(416) := X"00000000";
        ram_buffer(417) := X"03C0E821";
        ram_buffer(418) := X"8FBF001C";
        ram_buffer(419) := X"8FBE0018";
        ram_buffer(420) := X"27BD0020";
        ram_buffer(421) := X"03E00008";
        ram_buffer(422) := X"00000000";
        ram_buffer(423) := X"27BDFFE0";
        ram_buffer(424) := X"AFBF001C";
        ram_buffer(425) := X"AFBE0018";
        ram_buffer(426) := X"03A0F021";
        ram_buffer(427) := X"AFC40020";
        ram_buffer(428) := X"8FC20020";
        ram_buffer(429) := X"00000000";
        ram_buffer(430) := X"AFC20010";
        ram_buffer(431) := X"3C020000";
        ram_buffer(432) := X"24440B30";
        ram_buffer(433) := X"0C000277";
        ram_buffer(434) := X"00000000";
        ram_buffer(435) := X"8FC20010";
        ram_buffer(436) := X"00000000";
        ram_buffer(437) := X"00402021";
        ram_buffer(438) := X"0C0000A7";
        ram_buffer(439) := X"00000000";
        ram_buffer(440) := X"00402021";
        ram_buffer(441) := X"0C000277";
        ram_buffer(442) := X"00000000";
        ram_buffer(443) := X"3C020000";
        ram_buffer(444) := X"24440B44";
        ram_buffer(445) := X"0C000277";
        ram_buffer(446) := X"00000000";
        ram_buffer(447) := X"8FC20010";
        ram_buffer(448) := X"00000000";
        ram_buffer(449) := X"0040F809";
        ram_buffer(450) := X"00000000";
        ram_buffer(451) := X"00000000";
        ram_buffer(452) := X"03C0E821";
        ram_buffer(453) := X"8FBF001C";
        ram_buffer(454) := X"8FBE0018";
        ram_buffer(455) := X"27BD0020";
        ram_buffer(456) := X"03E00008";
        ram_buffer(457) := X"00000000";
        ram_buffer(458) := X"27BDFFD0";
        ram_buffer(459) := X"AFBF002C";
        ram_buffer(460) := X"AFBE0028";
        ram_buffer(461) := X"03A0F021";
        ram_buffer(462) := X"3C021050";
        ram_buffer(463) := X"AFC20018";
        ram_buffer(464) := X"AFC00010";
        ram_buffer(465) := X"1000000D";
        ram_buffer(466) := X"00000000";
        ram_buffer(467) := X"8FC20010";
        ram_buffer(468) := X"8FC30018";
        ram_buffer(469) := X"00000000";
        ram_buffer(470) := X"00621021";
        ram_buffer(471) := X"8FC30010";
        ram_buffer(472) := X"00000000";
        ram_buffer(473) := X"306300FF";
        ram_buffer(474) := X"A0430000";
        ram_buffer(475) := X"8FC20010";
        ram_buffer(476) := X"00000000";
        ram_buffer(477) := X"24420001";
        ram_buffer(478) := X"AFC20010";
        ram_buffer(479) := X"8FC20010";
        ram_buffer(480) := X"00000000";
        ram_buffer(481) := X"28420078";
        ram_buffer(482) := X"1440FFF0";
        ram_buffer(483) := X"00000000";
        ram_buffer(484) := X"3C020000";
        ram_buffer(485) := X"24440B48";
        ram_buffer(486) := X"0C000277";
        ram_buffer(487) := X"00000000";
        ram_buffer(488) := X"AFC00010";
        ram_buffer(489) := X"10000055";
        ram_buffer(490) := X"00000000";
        ram_buffer(491) := X"8FC20010";
        ram_buffer(492) := X"8FC30018";
        ram_buffer(493) := X"00000000";
        ram_buffer(494) := X"00621021";
        ram_buffer(495) := X"8C420000";
        ram_buffer(496) := X"00000000";
        ram_buffer(497) := X"AFC2001C";
        ram_buffer(498) := X"8FC20010";
        ram_buffer(499) := X"00000000";
        ram_buffer(500) := X"00021E00";
        ram_buffer(501) := X"8FC20010";
        ram_buffer(502) := X"00000000";
        ram_buffer(503) := X"24420001";
        ram_buffer(504) := X"00021400";
        ram_buffer(505) := X"00621821";
        ram_buffer(506) := X"8FC20010";
        ram_buffer(507) := X"00000000";
        ram_buffer(508) := X"24420002";
        ram_buffer(509) := X"00021200";
        ram_buffer(510) := X"00621821";
        ram_buffer(511) := X"8FC20010";
        ram_buffer(512) := X"00000000";
        ram_buffer(513) := X"24420003";
        ram_buffer(514) := X"00621021";
        ram_buffer(515) := X"AFC20020";
        ram_buffer(516) := X"8FC3001C";
        ram_buffer(517) := X"8FC20020";
        ram_buffer(518) := X"00000000";
        ram_buffer(519) := X"10620033";
        ram_buffer(520) := X"00000000";
        ram_buffer(521) := X"3C020000";
        ram_buffer(522) := X"24440B60";
        ram_buffer(523) := X"0C000277";
        ram_buffer(524) := X"00000000";
        ram_buffer(525) := X"3C020000";
        ram_buffer(526) := X"24440B84";
        ram_buffer(527) := X"0C000277";
        ram_buffer(528) := X"00000000";
        ram_buffer(529) := X"8FC2001C";
        ram_buffer(530) := X"00000000";
        ram_buffer(531) := X"00402021";
        ram_buffer(532) := X"0C0000A7";
        ram_buffer(533) := X"00000000";
        ram_buffer(534) := X"00402021";
        ram_buffer(535) := X"0C000277";
        ram_buffer(536) := X"00000000";
        ram_buffer(537) := X"AFC00014";
        ram_buffer(538) := X"10000005";
        ram_buffer(539) := X"00000000";
        ram_buffer(540) := X"8FC20014";
        ram_buffer(541) := X"00000000";
        ram_buffer(542) := X"24420001";
        ram_buffer(543) := X"AFC20014";
        ram_buffer(544) := X"8FC30014";
        ram_buffer(545) := X"3C02001E";
        ram_buffer(546) := X"34428480";
        ram_buffer(547) := X"0062102A";
        ram_buffer(548) := X"1440FFF7";
        ram_buffer(549) := X"00000000";
        ram_buffer(550) := X"3C020000";
        ram_buffer(551) := X"24440B8C";
        ram_buffer(552) := X"0C000277";
        ram_buffer(553) := X"00000000";
        ram_buffer(554) := X"8FC20020";
        ram_buffer(555) := X"00000000";
        ram_buffer(556) := X"00402021";
        ram_buffer(557) := X"0C0000A7";
        ram_buffer(558) := X"00000000";
        ram_buffer(559) := X"00402021";
        ram_buffer(560) := X"0C000277";
        ram_buffer(561) := X"00000000";
        ram_buffer(562) := X"240400FE";
        ram_buffer(563) := X"0C00026E";
        ram_buffer(564) := X"00000000";
        ram_buffer(565) := X"3C020000";
        ram_buffer(566) := X"24440B44";
        ram_buffer(567) := X"0C000277";
        ram_buffer(568) := X"00000000";
        ram_buffer(569) := X"1000FFFF";
        ram_buffer(570) := X"00000000";
        ram_buffer(571) := X"8FC20010";
        ram_buffer(572) := X"00000000";
        ram_buffer(573) := X"24420004";
        ram_buffer(574) := X"AFC20010";
        ram_buffer(575) := X"8FC20010";
        ram_buffer(576) := X"00000000";
        ram_buffer(577) := X"28420078";
        ram_buffer(578) := X"1440FFA8";
        ram_buffer(579) := X"00000000";
        ram_buffer(580) := X"3C020000";
        ram_buffer(581) := X"24440B98";
        ram_buffer(582) := X"0C000277";
        ram_buffer(583) := X"00000000";
        ram_buffer(584) := X"00000000";
        ram_buffer(585) := X"03C0E821";
        ram_buffer(586) := X"8FBF002C";
        ram_buffer(587) := X"8FBE0028";
        ram_buffer(588) := X"27BD0030";
        ram_buffer(589) := X"03E00008";
        ram_buffer(590) := X"00000000";
        ram_buffer(591) := X"27BDFFE0";
        ram_buffer(592) := X"AFBF001C";
        ram_buffer(593) := X"AFBE0018";
        ram_buffer(594) := X"03A0F021";
        ram_buffer(595) := X"3C021000";
        ram_buffer(596) := X"8C420000";
        ram_buffer(597) := X"00000000";
        ram_buffer(598) := X"AFC20010";
        ram_buffer(599) := X"8FC20010";
        ram_buffer(600) := X"00000000";
        ram_buffer(601) := X"00021603";
        ram_buffer(602) := X"AFC20014";
        ram_buffer(603) := X"8FC30014";
        ram_buffer(604) := X"2402003C";
        ram_buffer(605) := X"14620006";
        ram_buffer(606) := X"00000000";
        ram_buffer(607) := X"3C041000";
        ram_buffer(608) := X"0C0001A7";
        ram_buffer(609) := X"00000000";
        ram_buffer(610) := X"10000004";
        ram_buffer(611) := X"00000000";
        ram_buffer(612) := X"3C041008";
        ram_buffer(613) := X"0C0001A7";
        ram_buffer(614) := X"00000000";
        ram_buffer(615) := X"00001021";
        ram_buffer(616) := X"03C0E821";
        ram_buffer(617) := X"8FBF001C";
        ram_buffer(618) := X"8FBE0018";
        ram_buffer(619) := X"27BD0020";
        ram_buffer(620) := X"03E00008";
        ram_buffer(621) := X"00000000";
        ram_buffer(622) := X"3C032000";
        ram_buffer(623) := X"8C620020";
        ram_buffer(624) := X"00000000";
        ram_buffer(625) := X"30420002";
        ram_buffer(626) := X"1040FFFB";
        ram_buffer(627) := X"00000000";
        ram_buffer(628) := X"AC640000";
        ram_buffer(629) := X"03E00008";
        ram_buffer(630) := X"00001021";
        ram_buffer(631) := X"80820000";
        ram_buffer(632) := X"00000000";
        ram_buffer(633) := X"10400011";
        ram_buffer(634) := X"2406000A";
        ram_buffer(635) := X"2407000D";
        ram_buffer(636) := X"10460011";
        ram_buffer(637) := X"3C032000";
        ram_buffer(638) := X"24840001";
        ram_buffer(639) := X"8085FFFF";
        ram_buffer(640) := X"3C032000";
        ram_buffer(641) := X"8C620020";
        ram_buffer(642) := X"00000000";
        ram_buffer(643) := X"30420002";
        ram_buffer(644) := X"1040FFFB";
        ram_buffer(645) := X"00000000";
        ram_buffer(646) := X"AC650000";
        ram_buffer(647) := X"80820000";
        ram_buffer(648) := X"00000000";
        ram_buffer(649) := X"1440FFF2";
        ram_buffer(650) := X"00000000";
        ram_buffer(651) := X"03E00008";
        ram_buffer(652) := X"00001021";
        ram_buffer(653) := X"3C032000";
        ram_buffer(654) := X"8C620020";
        ram_buffer(655) := X"00000000";
        ram_buffer(656) := X"30420002";
        ram_buffer(657) := X"1040FFFB";
        ram_buffer(658) := X"00000000";
        ram_buffer(659) := X"AC670000";
        ram_buffer(660) := X"1000FFEA";
        ram_buffer(661) := X"24840001";
        ram_buffer(662) := X"2406001C";
        ram_buffer(663) := X"2407FFFC";
        ram_buffer(664) := X"00C41006";
        ram_buffer(665) := X"3042000F";
        ram_buffer(666) := X"2C43000A";
        ram_buffer(667) := X"1060000E";
        ram_buffer(668) := X"24450057";
        ram_buffer(669) := X"24450030";
        ram_buffer(670) := X"3C032000";
        ram_buffer(671) := X"8C620020";
        ram_buffer(672) := X"00000000";
        ram_buffer(673) := X"30420002";
        ram_buffer(674) := X"1040FFFB";
        ram_buffer(675) := X"00000000";
        ram_buffer(676) := X"24C6FFFC";
        ram_buffer(677) := X"AC650000";
        ram_buffer(678) := X"14C7FFF2";
        ram_buffer(679) := X"00C41006";
        ram_buffer(680) := X"03E00008";
        ram_buffer(681) := X"00000000";
        ram_buffer(682) := X"3C032000";
        ram_buffer(683) := X"8C620020";
        ram_buffer(684) := X"00000000";
        ram_buffer(685) := X"30420002";
        ram_buffer(686) := X"1040FFFB";
        ram_buffer(687) := X"00000000";
        ram_buffer(688) := X"24C6FFFC";
        ram_buffer(689) := X"AC650000";
        ram_buffer(690) := X"14C7FFE6";
        ram_buffer(691) := X"00C41006";
        ram_buffer(692) := X"1000FFF3";
        ram_buffer(693) := X"00000000";
        ram_buffer(694) := X"3C032000";
        ram_buffer(695) := X"8C620020";
        ram_buffer(696) := X"00000000";
        ram_buffer(697) := X"30420002";
        ram_buffer(698) := X"1040FFFC";
        ram_buffer(699) := X"24020049";
        ram_buffer(700) := X"AC620000";
        ram_buffer(701) := X"03E00008";
        ram_buffer(702) := X"00000000";
        ram_buffer(703) := X"3C022000";
        ram_buffer(704) := X"8C420020";
        ram_buffer(705) := X"03E00008";
        ram_buffer(706) := X"30420001";
        ram_buffer(707) := X"3C032000";
        ram_buffer(708) := X"8C620020";
        ram_buffer(709) := X"00000000";
        ram_buffer(710) := X"30420001";
        ram_buffer(711) := X"1040FFFB";
        ram_buffer(712) := X"00000000";
        ram_buffer(713) := X"8C620000";
        ram_buffer(714) := X"03E00008";
        ram_buffer(715) := X"00000000";
        ram_buffer(716) := X"4A756D70";
        ram_buffer(717) := X"696E6720";
        ram_buffer(718) := X"61742061";
        ram_buffer(719) := X"64647265";
        ram_buffer(720) := X"73732000";
        ram_buffer(721) := X"0A000000";
        ram_buffer(722) := X"43686563";
        ram_buffer(723) := X"6B696E67";
        ram_buffer(724) := X"20444452";
        ram_buffer(725) := X"202E2E2E";
        ram_buffer(726) := X"2E2E2E2E";
        ram_buffer(727) := X"20000000";
        ram_buffer(728) := X"4552524F";
        ram_buffer(729) := X"523A2043";
        ram_buffer(730) := X"616E6E6F";
        ram_buffer(731) := X"74206163";
        ram_buffer(732) := X"63657373";
        ram_buffer(733) := X"20444452";
        ram_buffer(734) := X"206D656D";
        ram_buffer(735) := X"6F727921";
        ram_buffer(736) := X"00000000";
        ram_buffer(737) := X"52656164";
        ram_buffer(738) := X"3A200000";
        ram_buffer(739) := X"45787065";
        ram_buffer(740) := X"63746564";
        ram_buffer(741) := X"3A200000";
        ram_buffer(742) := X"4F4B210A";
        ram_buffer(743) := X"00000000";
        return ram_buffer;
    end;
end;
