library ieee;
use ieee.std_logic_1164.all;

package main_pack_opcodes is

    constant cpu_width : integer := 32;
    constant ram_size : integer := 977;
    subtype word_type is std_logic_vector(cpu_width-1 downto 0);
    type ram_type is array(0 to ram_size-1) of word_type;
    function load_hex return ram_type;
end package;

package body main_pack_opcodes is

    function load_hex return ram_type is
		variable ram : ram_type := (others=>(others=>'0'));
    begin
        ram(0) := X"3C1C1001";
        ram(1) := X"279C8F4C";
        ram(2) := X"3C041000";
        ram(3) := X"24840F60";
        ram(4) := X"3C051000";
        ram(5) := X"24A50F60";
        ram(6) := X"00000000";
        ram(7) := X"00000000";
        ram(8) := X"10000009";
        ram(9) := X"00000000";
        ram(10) := X"00000000";
        ram(11) := X"3C1A1000";
        ram(12) := X"375A003C";
        ram(13) := X"03400008";
        ram(14) := X"00000000";
        ram(15) := X"401A7000";
        ram(16) := X"03400008";
        ram(17) := X"20840005";
        ram(18) := X"40806000";
        ram(19) := X"3C142000";
        ram(20) := X"3415000A";
        ram(21) := X"34160058";
        ram(22) := X"3417000D";
        ram(23) := X"34180F80";
        ram(24) := X"A2970000";
        ram(25) := X"A2950000";
        ram(26) := X"A2970000";
        ram(27) := X"A2950000";
        ram(28) := X"A2970000";
        ram(29) := X"A2950000";
        ram(30) := X"A2970000";
        ram(31) := X"A2950000";
        ram(32) := X"3C051000";
        ram(33) := X"24A5002C";
        ram(34) := X"20A6F000";
        ram(35) := X"18C00008";
        ram(36) := X"8CA60000";
        ram(37) := X"AC06003C";
        ram(38) := X"8CA60004";
        ram(39) := X"AC060040";
        ram(40) := X"8CA60008";
        ram(41) := X"AC060044";
        ram(42) := X"8CA6000C";
        ram(43) := X"AC060048";
        ram(44) := X"34020041";
        ram(45) := X"A2820000";
        ram(46) := X"34020072";
        ram(47) := X"A2820000";
        ram(48) := X"34020069";
        ram(49) := X"A2820000";
        ram(50) := X"34020074";
        ram(51) := X"A2820000";
        ram(52) := X"34020068";
        ram(53) := X"A2820000";
        ram(54) := X"A2970000";
        ram(55) := X"A2950000";
        ram(56) := X"34020061";
        ram(57) := X"A2820000";
        ram(58) := X"34030005";
        ram(59) := X"3404003C";
        ram(60) := X"00641020";
        ram(61) := X"A2820000";
        ram(62) := X"A2970000";
        ram(63) := X"A2950000";
        ram(64) := X"34020062";
        ram(65) := X"A2820000";
        ram(66) := X"3404003C";
        ram(67) := X"20820005";
        ram(68) := X"A2820000";
        ram(69) := X"A2970000";
        ram(70) := X"A2950000";
        ram(71) := X"34020063";
        ram(72) := X"A2820000";
        ram(73) := X"34040032";
        ram(74) := X"2485000F";
        ram(75) := X"A2850000";
        ram(76) := X"A2970000";
        ram(77) := X"A2950000";
        ram(78) := X"34020064";
        ram(79) := X"A2820000";
        ram(80) := X"34030005";
        ram(81) := X"3404003C";
        ram(82) := X"00641020";
        ram(83) := X"A2820000";
        ram(84) := X"A2970000";
        ram(85) := X"A2950000";
        ram(86) := X"34020065";
        ram(87) := X"A2820000";
        ram(88) := X"34021DDE";
        ram(89) := X"34030075";
        ram(90) := X"14600002";
        ram(91) := X"0043001A";
        ram(92) := X"0007000D";
        ram(93) := X"2401FFFF";
        ram(94) := X"14610004";
        ram(95) := X"3C018000";
        ram(96) := X"14410002";
        ram(97) := X"00000000";
        ram(98) := X"0006000D";
        ram(99) := X"00001012";
        ram(100) := X"00000000";
        ram(101) := X"00002012";
        ram(102) := X"A2840000";
        ram(103) := X"00002010";
        ram(104) := X"20840019";
        ram(105) := X"A2840000";
        ram(106) := X"2402FB07";
        ram(107) := X"34030013";
        ram(108) := X"14600002";
        ram(109) := X"0043001A";
        ram(110) := X"0007000D";
        ram(111) := X"2401FFFF";
        ram(112) := X"14610004";
        ram(113) := X"3C018000";
        ram(114) := X"14410002";
        ram(115) := X"00000000";
        ram(116) := X"0006000D";
        ram(117) := X"00001012";
        ram(118) := X"00000000";
        ram(119) := X"00002012";
        ram(120) := X"00042022";
        ram(121) := X"A2840000";
        ram(122) := X"3402061C";
        ram(123) := X"2403FFE9";
        ram(124) := X"14600002";
        ram(125) := X"0043001A";
        ram(126) := X"0007000D";
        ram(127) := X"2401FFFF";
        ram(128) := X"14610004";
        ram(129) := X"3C018000";
        ram(130) := X"14410002";
        ram(131) := X"00000000";
        ram(132) := X"0006000D";
        ram(133) := X"00001012";
        ram(134) := X"00000000";
        ram(135) := X"00002012";
        ram(136) := X"00042022";
        ram(137) := X"A2840000";
        ram(138) := X"2402FC7F";
        ram(139) := X"2403FFF3";
        ram(140) := X"14600002";
        ram(141) := X"0043001A";
        ram(142) := X"0007000D";
        ram(143) := X"2401FFFF";
        ram(144) := X"14610004";
        ram(145) := X"3C018000";
        ram(146) := X"14410002";
        ram(147) := X"00000000";
        ram(148) := X"0006000D";
        ram(149) := X"00001012";
        ram(150) := X"00002012";
        ram(151) := X"A2840000";
        ram(152) := X"2402FFFB";
        ram(153) := X"2403000C";
        ram(154) := X"14600002";
        ram(155) := X"0043001A";
        ram(156) := X"0007000D";
        ram(157) := X"2401FFFF";
        ram(158) := X"14610004";
        ram(159) := X"3C018000";
        ram(160) := X"14410002";
        ram(161) := X"00000000";
        ram(162) := X"0006000D";
        ram(163) := X"00001012";
        ram(164) := X"00002010";
        ram(165) := X"2484004B";
        ram(166) := X"A2840000";
        ram(167) := X"A2970000";
        ram(168) := X"A2950000";
        ram(169) := X"34020066";
        ram(170) := X"A2820000";
        ram(171) := X"3402034D";
        ram(172) := X"3403000D";
        ram(173) := X"14600002";
        ram(174) := X"0043001B";
        ram(175) := X"0007000D";
        ram(176) := X"00001012";
        ram(177) := X"00000000";
        ram(178) := X"00002012";
        ram(179) := X"A2840000";
        ram(180) := X"A2970000";
        ram(181) := X"A2950000";
        ram(182) := X"34020067";
        ram(183) := X"A2820000";
        ram(184) := X"34020005";
        ram(185) := X"3403000D";
        ram(186) := X"00430018";
        ram(187) := X"00000000";
        ram(188) := X"00002012";
        ram(189) := X"A2840000";
        ram(190) := X"2402FFFB";
        ram(191) := X"3403000D";
        ram(192) := X"00430018";
        ram(193) := X"00002810";
        ram(194) := X"00002012";
        ram(195) := X"00042022";
        ram(196) := X"00852021";
        ram(197) := X"20840002";
        ram(198) := X"A2840000";
        ram(199) := X"34020005";
        ram(200) := X"2403FFF3";
        ram(201) := X"00430018";
        ram(202) := X"00002810";
        ram(203) := X"00002012";
        ram(204) := X"00042022";
        ram(205) := X"00852021";
        ram(206) := X"20840003";
        ram(207) := X"A2840000";
        ram(208) := X"2402FFFB";
        ram(209) := X"2403FFF3";
        ram(210) := X"00430018";
        ram(211) := X"00002810";
        ram(212) := X"00002012";
        ram(213) := X"00852021";
        ram(214) := X"20840003";
        ram(215) := X"A2840000";
        ram(216) := X"3C04FE98";
        ram(217) := X"348462E5";
        ram(218) := X"3C050006";
        ram(219) := X"34A58DB8";
        ram(220) := X"00850018";
        ram(221) := X"00003010";
        ram(222) := X"24C7097A";
        ram(223) := X"A2870000";
        ram(224) := X"2402FFFF";
        ram(225) := X"24030000";
        ram(226) := X"00430018";
        ram(227) := X"00002010";
        ram(228) := X"24840046";
        ram(229) := X"A2840000";
        ram(230) := X"00620018";
        ram(231) := X"00002010";
        ram(232) := X"24840047";
        ram(233) := X"A2840000";
        ram(234) := X"A2970000";
        ram(235) := X"A2950000";
        ram(236) := X"34020068";
        ram(237) := X"A2820000";
        ram(238) := X"34020005";
        ram(239) := X"3403000D";
        ram(240) := X"00430019";
        ram(241) := X"00000000";
        ram(242) := X"00002012";
        ram(243) := X"A2840000";
        ram(244) := X"A2970000";
        ram(245) := X"A2950000";
        ram(246) := X"34020069";
        ram(247) := X"A2820000";
        ram(248) := X"3402000A";
        ram(249) := X"3403000C";
        ram(250) := X"0043202A";
        ram(251) := X"20850040";
        ram(252) := X"A2850000";
        ram(253) := X"0062202A";
        ram(254) := X"20850042";
        ram(255) := X"A2850000";
        ram(256) := X"2402FFF0";
        ram(257) := X"0043202A";
        ram(258) := X"20850042";
        ram(259) := X"A2850000";
        ram(260) := X"0062202A";
        ram(261) := X"20850044";
        ram(262) := X"A2850000";
        ram(263) := X"2403FFFF";
        ram(264) := X"0043202A";
        ram(265) := X"20850044";
        ram(266) := X"A2850000";
        ram(267) := X"0062202A";
        ram(268) := X"20850046";
        ram(269) := X"A2850000";
        ram(270) := X"A2970000";
        ram(271) := X"A2950000";
        ram(272) := X"3402006A";
        ram(273) := X"A2820000";
        ram(274) := X"3402000A";
        ram(275) := X"2844000C";
        ram(276) := X"20850040";
        ram(277) := X"A2850000";
        ram(278) := X"28440008";
        ram(279) := X"20850042";
        ram(280) := X"A2850000";
        ram(281) := X"A2970000";
        ram(282) := X"A2950000";
        ram(283) := X"3402006B";
        ram(284) := X"A2820000";
        ram(285) := X"3402000A";
        ram(286) := X"2C44000C";
        ram(287) := X"20850040";
        ram(288) := X"A2850000";
        ram(289) := X"2C440008";
        ram(290) := X"20850042";
        ram(291) := X"A2850000";
        ram(292) := X"A2970000";
        ram(293) := X"A2950000";
        ram(294) := X"3402006C";
        ram(295) := X"A2820000";
        ram(296) := X"3402000A";
        ram(297) := X"3403000C";
        ram(298) := X"0043202A";
        ram(299) := X"20850040";
        ram(300) := X"A2850000";
        ram(301) := X"0062202A";
        ram(302) := X"20850042";
        ram(303) := X"A2850000";
        ram(304) := X"A2970000";
        ram(305) := X"A2950000";
        ram(306) := X"3402006D";
        ram(307) := X"A2820000";
        ram(308) := X"34030046";
        ram(309) := X"34040005";
        ram(310) := X"00641022";
        ram(311) := X"A2820000";
        ram(312) := X"A2970000";
        ram(313) := X"A2950000";
        ram(314) := X"3402006E";
        ram(315) := X"A2820000";
        ram(316) := X"34030046";
        ram(317) := X"34040005";
        ram(318) := X"00641022";
        ram(319) := X"A2820000";
        ram(320) := X"A2970000";
        ram(321) := X"A2950000";
        ram(322) := X"34020042";
        ram(323) := X"A2820000";
        ram(324) := X"34020072";
        ram(325) := X"A2820000";
        ram(326) := X"34020061";
        ram(327) := X"A2820000";
        ram(328) := X"3402006E";
        ram(329) := X"A2820000";
        ram(330) := X"34020063";
        ram(331) := X"A2820000";
        ram(332) := X"34020068";
        ram(333) := X"A2820000";
        ram(334) := X"A2970000";
        ram(335) := X"A2950000";
        ram(336) := X"34020061";
        ram(337) := X"A2820000";
        ram(338) := X"340A0041";
        ram(339) := X"340B0042";
        ram(340) := X"10000002";
        ram(341) := X"A28A0000";
        ram(342) := X"A2960000";
        ram(343) := X"A28B0000";
        ram(344) := X"A2970000";
        ram(345) := X"A2950000";
        ram(346) := X"34020062";
        ram(347) := X"A2820000";
        ram(348) := X"340A0041";
        ram(349) := X"340B0042";
        ram(350) := X"340C0043";
        ram(351) := X"340D0044";
        ram(352) := X"340E0045";
        ram(353) := X"340F0058";
        ram(354) := X"04110005";
        ram(355) := X"A28A0000";
        ram(356) := X"A28D0000";
        ram(357) := X"10000006";
        ram(358) := X"A28E0000";
        ram(359) := X"A28F0000";
        ram(360) := X"A28B0000";
        ram(361) := X"03E00008";
        ram(362) := X"A28C0000";
        ram(363) := X"A2960000";
        ram(364) := X"A2970000";
        ram(365) := X"A2950000";
        ram(366) := X"34020063";
        ram(367) := X"A2820000";
        ram(368) := X"340A0041";
        ram(369) := X"340B0042";
        ram(370) := X"340C0043";
        ram(371) := X"340D0044";
        ram(372) := X"34020064";
        ram(373) := X"3403007B";
        ram(374) := X"3404007B";
        ram(375) := X"10430005";
        ram(376) := X"A28A0000";
        ram(377) := X"A28B0000";
        ram(378) := X"10640002";
        ram(379) := X"A28C0000";
        ram(380) := X"A2960000";
        ram(381) := X"A28D0000";
        ram(382) := X"A2970000";
        ram(383) := X"A2950000";
        ram(384) := X"34020064";
        ram(385) := X"A2820000";
        ram(386) := X"340A0041";
        ram(387) := X"340B0042";
        ram(388) := X"340C0043";
        ram(389) := X"340D0044";
        ram(390) := X"340F0058";
        ram(391) := X"34020064";
        ram(392) := X"3C03FFFF";
        ram(393) := X"34631234";
        ram(394) := X"3404007B";
        ram(395) := X"04610005";
        ram(396) := X"A28A0000";
        ram(397) := X"A28B0000";
        ram(398) := X"04410002";
        ram(399) := X"A28C0000";
        ram(400) := X"A2960000";
        ram(401) := X"04010002";
        ram(402) := X"00000000";
        ram(403) := X"A28F0000";
        ram(404) := X"A28D0000";
        ram(405) := X"A2970000";
        ram(406) := X"A2950000";
        ram(407) := X"34020065";
        ram(408) := X"A2820000";
        ram(409) := X"340A0041";
        ram(410) := X"340B0042";
        ram(411) := X"340C0043";
        ram(412) := X"340D0044";
        ram(413) := X"340E0045";
        ram(414) := X"340F0058";
        ram(415) := X"3C03FFFF";
        ram(416) := X"34631234";
        ram(417) := X"04710008";
        ram(418) := X"00000000";
        ram(419) := X"A28A0000";
        ram(420) := X"04110005";
        ram(421) := X"00000000";
        ram(422) := X"A28D0000";
        ram(423) := X"10000006";
        ram(424) := X"A28E0000";
        ram(425) := X"A28F0000";
        ram(426) := X"A28B0000";
        ram(427) := X"03E00008";
        ram(428) := X"A28C0000";
        ram(429) := X"A2960000";
        ram(430) := X"A2970000";
        ram(431) := X"A2950000";
        ram(432) := X"34020066";
        ram(433) := X"A2820000";
        ram(434) := X"340A0041";
        ram(435) := X"340B0042";
        ram(436) := X"340C0043";
        ram(437) := X"340D0044";
        ram(438) := X"34020064";
        ram(439) := X"3C03FFFF";
        ram(440) := X"34631234";
        ram(441) := X"1C600005";
        ram(442) := X"A28A0000";
        ram(443) := X"A28B0000";
        ram(444) := X"1C400002";
        ram(445) := X"A28C0000";
        ram(446) := X"A2960000";
        ram(447) := X"A28D0000";
        ram(448) := X"A2970000";
        ram(449) := X"A2950000";
        ram(450) := X"34020067";
        ram(451) := X"A2820000";
        ram(452) := X"340A0041";
        ram(453) := X"340B0042";
        ram(454) := X"340C0043";
        ram(455) := X"340D0044";
        ram(456) := X"34020064";
        ram(457) := X"3C03FFFF";
        ram(458) := X"34631234";
        ram(459) := X"18400005";
        ram(460) := X"A28A0000";
        ram(461) := X"A28B0000";
        ram(462) := X"18600002";
        ram(463) := X"A28C0000";
        ram(464) := X"A2960000";
        ram(465) := X"18000002";
        ram(466) := X"00000000";
        ram(467) := X"A2960000";
        ram(468) := X"A28D0000";
        ram(469) := X"A2970000";
        ram(470) := X"A2950000";
        ram(471) := X"34020068";
        ram(472) := X"A2820000";
        ram(473) := X"340A0041";
        ram(474) := X"340B0042";
        ram(475) := X"340C0043";
        ram(476) := X"340D0044";
        ram(477) := X"340E0045";
        ram(478) := X"34020064";
        ram(479) := X"3C03FFFF";
        ram(480) := X"34631234";
        ram(481) := X"34040000";
        ram(482) := X"04400005";
        ram(483) := X"A28A0000";
        ram(484) := X"A28B0000";
        ram(485) := X"04600002";
        ram(486) := X"A28C0000";
        ram(487) := X"A2960000";
        ram(488) := X"04800002";
        ram(489) := X"00000000";
        ram(490) := X"A28D0000";
        ram(491) := X"A28E0000";
        ram(492) := X"A2970000";
        ram(493) := X"A2950000";
        ram(494) := X"34020069";
        ram(495) := X"A2820000";
        ram(496) := X"340A0041";
        ram(497) := X"340B0042";
        ram(498) := X"340C0043";
        ram(499) := X"340D0044";
        ram(500) := X"340E0045";
        ram(501) := X"340F0058";
        ram(502) := X"3C03FFFF";
        ram(503) := X"34631234";
        ram(504) := X"04100008";
        ram(505) := X"00000000";
        ram(506) := X"A28A0000";
        ram(507) := X"04700005";
        ram(508) := X"00000000";
        ram(509) := X"A28D0000";
        ram(510) := X"10000006";
        ram(511) := X"A28E0000";
        ram(512) := X"A28F0000";
        ram(513) := X"A28B0000";
        ram(514) := X"03E00008";
        ram(515) := X"A28C0000";
        ram(516) := X"A2960000";
        ram(517) := X"A2970000";
        ram(518) := X"A2950000";
        ram(519) := X"3402006A";
        ram(520) := X"A2820000";
        ram(521) := X"340A0041";
        ram(522) := X"340B0042";
        ram(523) := X"340C0043";
        ram(524) := X"340D0044";
        ram(525) := X"34020064";
        ram(526) := X"3403007B";
        ram(527) := X"3404007B";
        ram(528) := X"14640005";
        ram(529) := X"A28A0000";
        ram(530) := X"A28B0000";
        ram(531) := X"14430002";
        ram(532) := X"A28C0000";
        ram(533) := X"A2960000";
        ram(534) := X"A28D0000";
        ram(535) := X"A2970000";
        ram(536) := X"A2950000";
        ram(537) := X"3402006B";
        ram(538) := X"A2820000";
        ram(539) := X"340A0041";
        ram(540) := X"340B0042";
        ram(541) := X"340F0058";
        ram(542) := X"08000221";
        ram(543) := X"A28A0000";
        ram(544) := X"A28F0000";
        ram(545) := X"A28B0000";
        ram(546) := X"A2970000";
        ram(547) := X"A2950000";
        ram(548) := X"3402006C";
        ram(549) := X"A2820000";
        ram(550) := X"340A0041";
        ram(551) := X"340B0042";
        ram(552) := X"340C0043";
        ram(553) := X"340D0044";
        ram(554) := X"340E0045";
        ram(555) := X"340F0058";
        ram(556) := X"0C000232";
        ram(557) := X"A28A0000";
        ram(558) := X"A28D0000";
        ram(559) := X"10000006";
        ram(560) := X"A28E0000";
        ram(561) := X"A28F0000";
        ram(562) := X"A28B0000";
        ram(563) := X"03E00008";
        ram(564) := X"A28C0000";
        ram(565) := X"A2960000";
        ram(566) := X"A2970000";
        ram(567) := X"A2950000";
        ram(568) := X"3402006D";
        ram(569) := X"A2820000";
        ram(570) := X"340A0041";
        ram(571) := X"340B0042";
        ram(572) := X"340C0043";
        ram(573) := X"340D0044";
        ram(574) := X"340E0045";
        ram(575) := X"340F0058";
        ram(576) := X"3C031000";
        ram(577) := X"24630920";
        ram(578) := X"0060F809";
        ram(579) := X"A28A0000";
        ram(580) := X"A28D0000";
        ram(581) := X"10000006";
        ram(582) := X"A28E0000";
        ram(583) := X"A28F0000";
        ram(584) := X"A28B0000";
        ram(585) := X"03E00008";
        ram(586) := X"A28C0000";
        ram(587) := X"A2960000";
        ram(588) := X"A2970000";
        ram(589) := X"A2950000";
        ram(590) := X"3402006E";
        ram(591) := X"A2820000";
        ram(592) := X"340A0041";
        ram(593) := X"340B0042";
        ram(594) := X"340F0058";
        ram(595) := X"3C031000";
        ram(596) := X"24630960";
        ram(597) := X"00600008";
        ram(598) := X"A28A0000";
        ram(599) := X"A28F0000";
        ram(600) := X"A28B0000";
        ram(601) := X"A2970000";
        ram(602) := X"A2950000";
        ram(603) := X"3402006F";
        ram(604) := X"A2820000";
        ram(605) := X"34020041";
        ram(606) := X"00000000";
        ram(607) := X"A2820000";
        ram(608) := X"A2970000";
        ram(609) := X"A2950000";
        ram(610) := X"34020070";
        ram(611) := X"A2820000";
        ram(612) := X"3402007A";
        ram(613) := X"3404003B";
        ram(614) := X"0000000D";
        ram(615) := X"20840001";
        ram(616) := X"A2840000";
        ram(617) := X"A2970000";
        ram(618) := X"A2950000";
        ram(619) := X"34020071";
        ram(620) := X"A2820000";
        ram(621) := X"3404003D";
        ram(622) := X"0000000C";
        ram(623) := X"2084FFFF";
        ram(624) := X"A2840000";
        ram(625) := X"A2970000";
        ram(626) := X"A2950000";
        ram(627) := X"3402004C";
        ram(628) := X"A2820000";
        ram(629) := X"3402006F";
        ram(630) := X"A2820000";
        ram(631) := X"34020061";
        ram(632) := X"A2820000";
        ram(633) := X"34020064";
        ram(634) := X"A2820000";
        ram(635) := X"A2970000";
        ram(636) := X"A2950000";
        ram(637) := X"34020061";
        ram(638) := X"A2820000";
        ram(639) := X"00181025";
        ram(640) := X"3C034142";
        ram(641) := X"346343FC";
        ram(642) := X"AC430010";
        ram(643) := X"80440010";
        ram(644) := X"A2840000";
        ram(645) := X"80440011";
        ram(646) := X"A2840000";
        ram(647) := X"80440012";
        ram(648) := X"A2840000";
        ram(649) := X"80420013";
        ram(650) := X"00021A03";
        ram(651) := X"20630045";
        ram(652) := X"A2830000";
        ram(653) := X"20420049";
        ram(654) := X"A2820000";
        ram(655) := X"A2970000";
        ram(656) := X"A2950000";
        ram(657) := X"34020062";
        ram(658) := X"A2820000";
        ram(659) := X"00181025";
        ram(660) := X"3C034142";
        ram(661) := X"34634344";
        ram(662) := X"AC430010";
        ram(663) := X"80440010";
        ram(664) := X"A2840000";
        ram(665) := X"80440011";
        ram(666) := X"A2840000";
        ram(667) := X"80440012";
        ram(668) := X"A2840000";
        ram(669) := X"80420013";
        ram(670) := X"A2820000";
        ram(671) := X"A2970000";
        ram(672) := X"A2950000";
        ram(673) := X"34020063";
        ram(674) := X"A2820000";
        ram(675) := X"00181025";
        ram(676) := X"3C030041";
        ram(677) := X"34630042";
        ram(678) := X"AC430010";
        ram(679) := X"84440010";
        ram(680) := X"A2840000";
        ram(681) := X"84420012";
        ram(682) := X"A2820000";
        ram(683) := X"A2970000";
        ram(684) := X"A2950000";
        ram(685) := X"34020064";
        ram(686) := X"A2820000";
        ram(687) := X"00181025";
        ram(688) := X"3C030041";
        ram(689) := X"34630042";
        ram(690) := X"AC430010";
        ram(691) := X"84440010";
        ram(692) := X"A2840000";
        ram(693) := X"84420012";
        ram(694) := X"A2820000";
        ram(695) := X"A2970000";
        ram(696) := X"A2950000";
        ram(697) := X"34020065";
        ram(698) := X"A2820000";
        ram(699) := X"00181025";
        ram(700) := X"24030041";
        ram(701) := X"AC430010";
        ram(702) := X"34030000";
        ram(703) := X"8C420010";
        ram(704) := X"A2820000";
        ram(705) := X"A2970000";
        ram(706) := X"A2950000";
        ram(707) := X"34020066";
        ram(708) := X"A2820000";
        ram(709) := X"00181025";
        ram(710) := X"24030041";
        ram(711) := X"AC430010";
        ram(712) := X"34030000";
        ram(713) := X"88420010";
        ram(714) := X"98420010";
        ram(715) := X"A2820000";
        ram(716) := X"A2970000";
        ram(717) := X"A2950000";
        ram(718) := X"34020067";
        ram(719) := X"A2820000";
        ram(720) := X"34020041";
        ram(721) := X"A2820000";
        ram(722) := X"A2970000";
        ram(723) := X"A2950000";
        ram(724) := X"34020068";
        ram(725) := X"A2820000";
        ram(726) := X"00182025";
        ram(727) := X"34024142";
        ram(728) := X"A4820010";
        ram(729) := X"80830010";
        ram(730) := X"A2830000";
        ram(731) := X"80820011";
        ram(732) := X"A2820000";
        ram(733) := X"A2970000";
        ram(734) := X"A2950000";
        ram(735) := X"34020069";
        ram(736) := X"A2820000";
        ram(737) := X"00181025";
        ram(738) := X"3C034142";
        ram(739) := X"34634344";
        ram(740) := X"AC430010";
        ram(741) := X"80440010";
        ram(742) := X"A2840000";
        ram(743) := X"80440011";
        ram(744) := X"A2840000";
        ram(745) := X"80440012";
        ram(746) := X"A2840000";
        ram(747) := X"80420013";
        ram(748) := X"A2820000";
        ram(749) := X"A2970000";
        ram(750) := X"A2950000";
        ram(751) := X"3402006A";
        ram(752) := X"A2820000";
        ram(753) := X"00181025";
        ram(754) := X"3C034142";
        ram(755) := X"34634344";
        ram(756) := X"A8430010";
        ram(757) := X"B8430010";
        ram(758) := X"80440010";
        ram(759) := X"A2840000";
        ram(760) := X"80440011";
        ram(761) := X"A2840000";
        ram(762) := X"80440012";
        ram(763) := X"A2840000";
        ram(764) := X"80420013";
        ram(765) := X"A2820000";
        ram(766) := X"A2970000";
        ram(767) := X"A2950000";
        ram(768) := X"3402004C";
        ram(769) := X"A2820000";
        ram(770) := X"3402006F";
        ram(771) := X"A2820000";
        ram(772) := X"34020067";
        ram(773) := X"A2820000";
        ram(774) := X"34020069";
        ram(775) := X"A2820000";
        ram(776) := X"34020063";
        ram(777) := X"A2820000";
        ram(778) := X"A2970000";
        ram(779) := X"A2950000";
        ram(780) := X"34020061";
        ram(781) := X"A2820000";
        ram(782) := X"34020741";
        ram(783) := X"340360F3";
        ram(784) := X"00432024";
        ram(785) := X"A2840000";
        ram(786) := X"A2970000";
        ram(787) := X"A2950000";
        ram(788) := X"34020062";
        ram(789) := X"A2820000";
        ram(790) := X"34020741";
        ram(791) := X"304460F3";
        ram(792) := X"A2840000";
        ram(793) := X"A2970000";
        ram(794) := X"A2950000";
        ram(795) := X"34020063";
        ram(796) := X"A2820000";
        ram(797) := X"3C020041";
        ram(798) := X"00021C02";
        ram(799) := X"A2830000";
        ram(800) := X"A2970000";
        ram(801) := X"A2950000";
        ram(802) := X"34020064";
        ram(803) := X"A2820000";
        ram(804) := X"3C02F0FF";
        ram(805) := X"3442F08E";
        ram(806) := X"3C030F0F";
        ram(807) := X"34630F30";
        ram(808) := X"00432027";
        ram(809) := X"A2840000";
        ram(810) := X"A2970000";
        ram(811) := X"A2950000";
        ram(812) := X"34020065";
        ram(813) := X"A2820000";
        ram(814) := X"34020040";
        ram(815) := X"34030001";
        ram(816) := X"00432025";
        ram(817) := X"A2840000";
        ram(818) := X"A2970000";
        ram(819) := X"A2950000";
        ram(820) := X"34020066";
        ram(821) := X"A2820000";
        ram(822) := X"34020040";
        ram(823) := X"34440001";
        ram(824) := X"A2840000";
        ram(825) := X"A2970000";
        ram(826) := X"A2950000";
        ram(827) := X"34020067";
        ram(828) := X"A2820000";
        ram(829) := X"3402F043";
        ram(830) := X"3403F002";
        ram(831) := X"00432026";
        ram(832) := X"A2840000";
        ram(833) := X"A2970000";
        ram(834) := X"A2950000";
        ram(835) := X"34020068";
        ram(836) := X"A2820000";
        ram(837) := X"3402F043";
        ram(838) := X"3844F002";
        ram(839) := X"A2840000";
        ram(840) := X"A2970000";
        ram(841) := X"A2950000";
        ram(842) := X"3402004D";
        ram(843) := X"A2820000";
        ram(844) := X"3402006F";
        ram(845) := X"A2820000";
        ram(846) := X"34020076";
        ram(847) := X"A2820000";
        ram(848) := X"34020065";
        ram(849) := X"A2820000";
        ram(850) := X"A2970000";
        ram(851) := X"A2950000";
        ram(852) := X"34020061";
        ram(853) := X"A2820000";
        ram(854) := X"34020041";
        ram(855) := X"00400011";
        ram(856) := X"00001810";
        ram(857) := X"A2830000";
        ram(858) := X"A2970000";
        ram(859) := X"A2950000";
        ram(860) := X"34020062";
        ram(861) := X"A2820000";
        ram(862) := X"34020041";
        ram(863) := X"00400013";
        ram(864) := X"00001812";
        ram(865) := X"A2830000";
        ram(866) := X"A2970000";
        ram(867) := X"A2950000";
        ram(868) := X"34020063";
        ram(869) := X"A2820000";
        ram(870) := X"34020041";
        ram(871) := X"00400011";
        ram(872) := X"00001810";
        ram(873) := X"A2830000";
        ram(874) := X"A2970000";
        ram(875) := X"A2950000";
        ram(876) := X"34020064";
        ram(877) := X"A2820000";
        ram(878) := X"34020041";
        ram(879) := X"00400013";
        ram(880) := X"00001812";
        ram(881) := X"A2830000";
        ram(882) := X"A2970000";
        ram(883) := X"A2950000";
        ram(884) := X"34020053";
        ram(885) := X"A2820000";
        ram(886) := X"34020068";
        ram(887) := X"A2820000";
        ram(888) := X"34020069";
        ram(889) := X"A2820000";
        ram(890) := X"34020066";
        ram(891) := X"A2820000";
        ram(892) := X"34020074";
        ram(893) := X"A2820000";
        ram(894) := X"A2970000";
        ram(895) := X"A2950000";
        ram(896) := X"34020061";
        ram(897) := X"A2820000";
        ram(898) := X"3C024041";
        ram(899) := X"34424243";
        ram(900) := X"00021A00";
        ram(901) := X"00031E02";
        ram(902) := X"A2830000";
        ram(903) := X"A2970000";
        ram(904) := X"A2950000";
        ram(905) := X"34020062";
        ram(906) := X"A2820000";
        ram(907) := X"3C024041";
        ram(908) := X"34424243";
        ram(909) := X"34030008";
        ram(910) := X"00621804";
        ram(911) := X"00031E02";
        ram(912) := X"A2830000";
        ram(913) := X"A2970000";
        ram(914) := X"A2950000";
        ram(915) := X"34020063";
        ram(916) := X"A2820000";
        ram(917) := X"3C024041";
        ram(918) := X"34424243";
        ram(919) := X"00021C03";
        ram(920) := X"A2830000";
        ram(921) := X"3C028400";
        ram(922) := X"00021E43";
        ram(923) := X"2063FF80";
        ram(924) := X"A2830000";
        ram(925) := X"A2970000";
        ram(926) := X"A2950000";
        ram(927) := X"34020064";
        ram(928) := X"A2820000";
        ram(929) := X"3C024041";
        ram(930) := X"34424243";
        ram(931) := X"34030010";
        ram(932) := X"00621807";
        ram(933) := X"A2830000";
        ram(934) := X"34030019";
        ram(935) := X"3C028400";
        ram(936) := X"00621807";
        ram(937) := X"2063FF80";
        ram(938) := X"A2830000";
        ram(939) := X"A2970000";
        ram(940) := X"A2950000";
        ram(941) := X"34020065";
        ram(942) := X"A2820000";
        ram(943) := X"3C024041";
        ram(944) := X"34424243";
        ram(945) := X"00021C02";
        ram(946) := X"A2830000";
        ram(947) := X"3C028400";
        ram(948) := X"00021E42";
        ram(949) := X"A2830000";
        ram(950) := X"A2970000";
        ram(951) := X"A2950000";
        ram(952) := X"34020066";
        ram(953) := X"A2820000";
        ram(954) := X"3C024041";
        ram(955) := X"34424243";
        ram(956) := X"34030010";
        ram(957) := X"00622006";
        ram(958) := X"A2840000";
        ram(959) := X"34030019";
        ram(960) := X"3C028400";
        ram(961) := X"00621806";
        ram(962) := X"A2830000";
        ram(963) := X"A2970000";
        ram(964) := X"A2950000";
        ram(965) := X"34020044";
        ram(966) := X"A2820000";
        ram(967) := X"3402006F";
        ram(968) := X"A2820000";
        ram(969) := X"3402006E";
        ram(970) := X"A2820000";
        ram(971) := X"34020065";
        ram(972) := X"A2820000";
        ram(973) := X"A2970000";
        ram(974) := X"A2950000";
        ram(975) := X"080003CF";
        ram(976) := X"00000000";
        return ram;
    end;
end;
